module hidden_5 (I0, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I16, I17, I18, I19, I20, I21, I22, I23, I24, I26, I27, I28, I29, I30, I31, I32, I34, I36, I38, I39, I40, I42, I43, I44, I45, I46, I48, I49, I50, I51, I52, I54, I55, I56, I57, I58, I60, I61, I62, I64, I65, I66, I68, I70, I71, I72, I74, I75, I76, I78, I79, I80, I81, I82, I84, I85, I86, I88, I90, I91, I92, I94, I95, I96, I98, I100, I102, I103, I104, I106, I108, I109, I110, I111, I112, I113, I114, I115, I116, I117, I118, I120, I121, I122, I123, I124, I126, I128, I130, I132, I134, I135, I136, I137, I138, I140, I142, I144, I145, I146, I147, I148, I150, I151, I152, I153, I154, I156, I157, I158, I160, I161, I162, I163, I164, I165, I166, I168, I169, I170, I171, I172, I174, I175, I176, I178, I179, I180, I181, I182, I184, I185, I186, I188, I190, I191, I192, I193, I194, I195, I196, I197, I198, O0, O1, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15, O16, O17, O18, O19, O20, O21, O22, O23, O24, O25, O26, O27, O28, O29, O30, O31, O32, O33, O34, O35, O36, O37, O38, O39, O40, O41, O42, O43, O44, O45, O46, O47, O48, O49, O50, O51, O52, O53, O54, O55, O56, O57, O58, O59, O60, O61, O62, O63, O64, O65, O66, O67, O68, O69, O70, O71, O72, O73, O74, O75, O76, O77, O78, O79, O80, O81, O82, O83, O84, O85, O86, O87, O88, O89, O90, O91, O92, O93, O94, O95, O96, O97, O98, O99, O100, O101, O102, O103, O104, O105, O106, O107, O108, O109, O110, O111, O112, O113, O114, O115, O116, O117, O118, O119, O120, O121, O122, O123, O124, O125, O126, O127, O128, O129, O130, O131, O132, O133, O134, O135, O136, O137, O138, O139, O140, O141, O142, O143, O144, O145, O146, O147, O148, O149, O150, O151, O152, O153, O154, O155, O156, O157, O158, O159, O160, O161, O162, O163, O164, O165, O166, O167, O168, O169, O170, O171, O172, O173, O174, O175, O176, O177, O178, O179, O180, O181, O182, O183, O184, O185, O186, O187, O188, O189, O190, O191, O192, O193, O194, O195, O196, O197, O198, O199, O200, O201, O202, O203, O204, O205, O206, O207, O208, O209, O210, O211, O212, O213, O214, O215, O216, O217, O218, O219, O220, O221, O222, O223, O224, O225, O226, O227, O228, O229, O230, O231, O232, O233, O234, O235, O236, O237, O238, O239, O240, O241, O242, O243, O244, O245, O246, O247, O248, O249, O250, O251, O252, O253, O254, O255, O256, O257, O258, O259, O260, O261, O262, O263, O264, O265, O266, O267, O268, O269, O270, O271, O272, O273, O274, O275, O276, O277, O278, O279, O280, O281, O282, O283, O284, O285, O286, O287, O288, O289, O290, O291, O292, O293, O294, O295, O296, O297, O298, O299, O300, O301, O302, O303, O304, O305, O306, O307, O308, O309, O310, O311, O312, O313, O314, O315, O316, O317, O318, O319, O320, O321, O322, O323, O324, O325, O326, O327, O328, O329, O330, O331, O332, O333, O334, O335, O336, O337, O338, O339, O340, O341, O342, O343, O344, O345, O346, O347, O348, O349, O350, O351, O352, O353, O354, O355, O356, O357, O358, O359, O360, O361, O362, O363, O364, O365, O366, O367, O368, O369, O370, O371, O372, O373, O374, O375, O376, O377, O378, O379, O380, O381, O382, O383, O384, O385, O386, O387, O388, O389, O390, O391, O392, O393, O394, O395, O396, O397, O398, O399, O400, O401, O402, O403, O404, O405, O406, O407, O408, O409, O410, O411, O412, O413, O414, O415, O416, O417, O418, O419, O420, O421, O422, O423, O424, O425, O426, O427, O428, O429, O430, O431, O432, O433, O434, O435, O436, O437, O438, O439, O440, O441, O442, O443, O444, O445, O446, O447, O448, O449, O450, O451, O452, O453, O454, O455, O456, O457, O458, O459, O460, O461, O462, O463, O464, O465, O466, O467, O468, O469, O470, O471, O472, O473, O474, O475, O476, O477, O478, O479, O480, O481, O482, O483, O484, O485, O486, O487, O488, O489, O490, O491, O492, O493, O494, O495, O496, O497, O498, O499, O500, O501, O502, O503, O504, O505, O506, O507, O508, O509, O510, O511, O512, O513, O514, O515, O516, O517, O518, O519, O520, O521, O522, O523, O524, O525, O526, O527, O528, O529, O530, O531, O532, O533, O534, O535, O536, O537, O538, O539, O540, O541, O542, O543, O544, O545, O546, O547, O548, O549, O550, O551, O552, O553, O554, O555, O556, O557, O558, O559, O560, O561, O562, O563, O564, O565, O566, O567, O568, O569, O570, O571, O572, O573, O574, O575, O576, O577, O578, O579, O580, O581, O582, O583, O584, O585, O586, O587, O588, O589, O590, O591, O592, O593, O594, O595, O596, O597, O598, O599, O600, O601, O602, O603, O604, O605, O606, O607, O608, O609, O610, O611, O612, O613, O614, O615, O616, O617, O618, O619, O620, O621, O622, O623, O624, O625, O626, O627, O628, O629, O630, O631, O632, O633, O634, O635, O636, O637, O638, O639, O640, O641, O642, O643, O644, O645, O646, O647, O648, O649, O650, O651, O652, O653, O654, O655, O656, O657, O658, O659, O660, O661, O662, O663, O664, O665, O666, O667, O668, O669, O670, O671, O672, O673, O674, O675, O676, O677, O678, O679, O680, O681, O682, O683, O684, O685, O686, O687, O688, O689, O690, O691, O692, O693, O694, O695, O696, O697, O698, O699, O700, O701, O702, O703, O704, O705, O706, O707, O708, O709, O710, O711, O712, O713, O714, O715, O716, O717, O718, O719, O720, O721, O722, O723, O724, O725, O726, O727, O728, O729, O730, O731, O732, O733, O734, O735, O736, O737, O738, O739, O740, O741, O742, O743, O744, O745, O746, O747, O748, O749, O750, O751, O752, O753, O754, O755, O756, O757, O758, O759, O760, O761, O762, O763, O764, O765, O766, O767, O768, O769, O770, O771, O772, O773, O774, O775, O776, O777, O778, O779, O780, O781, O782, O783, O784, O785, O786, O787, O788, O789, O790, O791, O792, O793, O794, O795, O796, O797, O798, O799, O800, O801, O802, O803, O804, O805, O806, O807, O808, O809, O810, O811, O812, O813, O814, O815, O816, O817, O818, O819, O820, O821, O822, O823, O824, O825, O826, O827, O828, O829, O830, O831, O832, O833, O834, O835, O836, O837, O838, O839, O840, O841, O842, O843, O844, O845, O846, O847, O848, O849, O850, O851, O852, O853, O854, O855, O856, O857, O858, O859, O860, O861, O862, O863, O864, O865, O866, O867, O868, O869, O870, O871, O872, O873, O874, O875, O876, O877, O878, O879, O880, O881, O882, O883, O884, O885, O886, O887, O888, O889, O890, O891, O892, O893, O894, O895, O896, O897, O898, O899, O900, O901, O902, O903, O904, O905, O906, O907, O908, O909, O910, O911, O912, O913, O914, O915, O916, O917, O918, O919, O920, O921, O922, O923, O924, O925, O926, O927, O928, O929, O930, O931, O932, O933, O934, O935, O936, O937, O938, O939, O940, O941, O942, O943, O944, O945, O946, O947, O948, O949, O950, O951, O952, O953, O954, O955, O956, O957, O958, O959, O960, O961, O962, O963, O964, O965, O966, O967, O968, O969, O970, O971, O972, O973, O974, O975, O976, O977, O978, O979, O980, O981, O982, O983, O984, O985, O986, O987, O988, O989, O990, O991, O992, O993, O994, O995, O996, O997, O998, O999, O1000, O1001, O1002, O1003, O1004, O1005, O1006, O1007, O1008, O1009, O1010, O1011, O1012, O1013, O1014, O1015, O1016, O1017, O1018, O1019, O1020, O1021, O1022, O1023, O1024, O1025, O1026, O1027, O1028, O1029, O1030, O1031, O1032, O1033, O1034, O1035, O1036, O1037, O1038, O1039, O1040, O1041, O1042, O1043, O1044, O1045, O1046, O1047, O1048, O1049, O1050, O1051, O1052, O1053, O1054, O1055, O1056, O1057, O1058, O1059, O1060, O1061, O1062, O1063, O1064, O1065, O1066, O1067, O1068, O1069, O1070, O1071, O1072, O1073, O1074, O1075, O1076, O1077, O1078, O1079, O1080, O1081, O1082, O1083, O1084, O1085, O1086, O1087, O1088, O1089, O1090, O1091, O1092, O1093, O1094, O1095, O1096, O1097, O1098, O1099, O1100, O1101, O1102, O1103, O1104, O1105, O1106, O1107, O1108, O1109, O1110, O1111, O1112, O1113, O1114, O1115, O1116, O1117, O1118, O1119, O1120, O1121, O1122, O1123, O1124, O1125, O1126, O1127, O1128, O1129, O1130, O1131, O1132, O1133, O1134, O1135, O1136, O1137, O1138, O1139, O1140, O1141, O1142, O1143, O1144, O1145, O1146, O1147, O1148, O1149, O1150, O1151, O1152, O1153, O1154, O1155, O1156, O1157, O1158, O1159, O1160, O1161, O1162, O1163, O1164, O1165, O1166, O1167, O1168, O1169, O1170, O1171, O1172, O1173, O1174, O1175, O1176, O1177, O1178, O1179, O1180, O1181, O1182, O1183, O1184, O1185, O1186, O1187, O1188, O1189, O1190, O1191, O1192, O1193, O1194, O1195, O1196, O1197, O1198, O1199, O1200, O1201, O1202, O1203, O1204, O1205, O1206, O1207, O1208, O1209, O1210, O1211, O1212, O1213, O1214, O1215, O1216, O1217, O1218, O1219, O1220, O1221, O1222, O1223, O1224, O1225, O1226, O1227, O1228, O1229, O1230, O1231, O1232, O1233, O1234, O1235, O1236, O1237, O1238, O1239, O1240, O1241, O1242, O1243, O1244, O1245, O1246, O1247, O1248, O1249, O1250, O1251, O1252, O1253, O1254, O1255, O1256, O1257, O1258, O1259, O1260, O1261, O1262, O1263, O1264, O1265, O1266, O1267, O1268, O1269, O1270, O1271, O1272, O1273, O1274, O1275, O1276, O1277, O1278, O1279, O1280, O1281, O1282, O1283, O1284, O1285, O1286, O1287, O1288, O1289, O1290, O1291, O1292, O1293, O1294, O1295, O1296, O1297, O1298, O1299, O1300, O1301, O1302, O1303, O1304, O1305, O1306, O1307, O1308, O1309, O1310, O1311, O1312, O1313, O1314, O1315, O1316, O1317, O1318, O1319, O1320, O1321, O1322, O1323, O1324, O1325, O1326, O1327, O1328, O1329, O1330, O1331, O1332, O1333, O1334, O1335, O1336, O1337, O1338, O1339, O1340, O1341, O1342, O1343, O1344, O1345, O1346, O1347, O1348, O1349, O1350, O1351, O1352, O1353, O1354, O1355, O1356, O1357, O1358, O1359, O1360, O1361, O1362, O1363, O1364, O1365, O1366, O1367, O1368, O1369, O1370, O1371, O1372, O1373, O1374, O1375, O1376, O1377, O1378, O1379, O1380, O1381, O1382, O1383, O1384, O1385, O1386, O1387, O1388, O1389, O1390, O1391, O1392, O1393, O1394, O1395, O1396, O1397, O1398, O1399, O1400, O1401, O1402, O1403, O1404, O1405, O1406, O1407, O1408, O1409, O1410, O1411, O1412, O1413, O1414, O1415, O1416, O1417, O1418, O1419, O1420, O1421, O1422, O1423, O1424, O1425, O1426, O1427, O1428, O1429, O1430, O1431, O1432, O1433, O1434, O1435, O1436, O1437, O1438, O1439, O1440, O1441, O1442, O1443, O1444, O1445, O1446, O1447, O1448, O1449, O1450, O1451, O1452, O1453, O1454, O1455, O1456, O1457, O1458, O1459, O1460, O1461, O1462, O1463, O1464, O1465, O1466, O1467, O1468, O1469, O1470, O1471, O1472, O1473, O1474, O1475, O1476, O1477, O1478, O1479, O1480, O1481, O1482, O1483, O1484, O1485, O1486, O1487, O1488, O1489, O1490, O1491, O1492, O1493, O1494, O1495, O1496, O1497, O1498, O1499, O1500, O1501, O1502, O1503, O1504, O1505, O1506, O1507, O1508, O1509, O1510, O1511, O1512, O1513, O1514, O1515, O1516, O1517, O1518, O1519, O1520, O1521, O1522, O1523, O1524, O1525, O1526, O1527, O1528, O1529, O1530, O1531, O1532, O1533, O1534, O1535, O1536, O1537, O1538, O1539, O1540, O1541, O1542, O1543, O1544, O1545, O1546, O1547, O1548, O1549, O1550, O1551, O1552, O1553, O1554, O1555, O1556, O1557, O1558, O1559, O1560, O1561, O1562, O1563, O1564, O1565, O1566, O1567, O1568, O1569, O1570, O1571, O1572, O1573, O1574, O1575, O1576, O1577, O1578, O1579, O1580, O1581, O1582, O1583, O1584, O1585, O1586, O1587, O1588, O1589, O1590, O1591, O1592, O1593, O1594, O1595, O1596, O1597, O1598, O1599, O1600, O1601, O1602, O1603, O1604, O1605, O1606, O1607, O1608, O1609, O1610, O1611, O1612, O1613, O1614, O1615, O1616, O1617, O1618, O1619, O1620, O1621, O1622, O1623, O1624, O1625, O1626, O1627, O1628, O1629, O1630, O1631, O1632, O1633);
  input I0, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I16, I17, I18, I19, I20, I21, I22, I23, I24, I26, I27, I28, I29, I30, I31, I32, I34, I36, I38, I39, I40, I42, I43, I44, I45, I46, I48, I49, I50, I51, I52, I54, I55, I56, I57, I58, I60, I61, I62, I64, I65, I66, I68, I70, I71, I72, I74, I75, I76, I78, I79, I80, I81, I82, I84, I85, I86, I88, I90, I91, I92, I94, I95, I96, I98, I100, I102, I103, I104, I106, I108, I109, I110, I111, I112, I113, I114, I115, I116, I117, I118, I120, I121, I122, I123, I124, I126, I128, I130, I132, I134, I135, I136, I137, I138, I140, I142, I144, I145, I146, I147, I148, I150, I151, I152, I153, I154, I156, I157, I158, I160, I161, I162, I163, I164, I165, I166, I168, I169, I170, I171, I172, I174, I175, I176, I178, I179, I180, I181, I182, I184, I185, I186, I188, I190, I191, I192, I193, I194, I195, I196, I197, I198;
  output O0, O1, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15, O16, O17, O18, O19, O20, O21, O22, O23, O24, O25, O26, O27, O28, O29, O30, O31, O32, O33, O34, O35, O36, O37, O38, O39, O40, O41, O42, O43, O44, O45, O46, O47, O48, O49, O50, O51, O52, O53, O54, O55, O56, O57, O58, O59, O60, O61, O62, O63, O64, O65, O66, O67, O68, O69, O70, O71, O72, O73, O74, O75, O76, O77, O78, O79, O80, O81, O82, O83, O84, O85, O86, O87, O88, O89, O90, O91, O92, O93, O94, O95, O96, O97, O98, O99, O100, O101, O102, O103, O104, O105, O106, O107, O108, O109, O110, O111, O112, O113, O114, O115, O116, O117, O118, O119, O120, O121, O122, O123, O124, O125, O126, O127, O128, O129, O130, O131, O132, O133, O134, O135, O136, O137, O138, O139, O140, O141, O142, O143, O144, O145, O146, O147, O148, O149, O150, O151, O152, O153, O154, O155, O156, O157, O158, O159, O160, O161, O162, O163, O164, O165, O166, O167, O168, O169, O170, O171, O172, O173, O174, O175, O176, O177, O178, O179, O180, O181, O182, O183, O184, O185, O186, O187, O188, O189, O190, O191, O192, O193, O194, O195, O196, O197, O198, O199, O200, O201, O202, O203, O204, O205, O206, O207, O208, O209, O210, O211, O212, O213, O214, O215, O216, O217, O218, O219, O220, O221, O222, O223, O224, O225, O226, O227, O228, O229, O230, O231, O232, O233, O234, O235, O236, O237, O238, O239, O240, O241, O242, O243, O244, O245, O246, O247, O248, O249, O250, O251, O252, O253, O254, O255, O256, O257, O258, O259, O260, O261, O262, O263, O264, O265, O266, O267, O268, O269, O270, O271, O272, O273, O274, O275, O276, O277, O278, O279, O280, O281, O282, O283, O284, O285, O286, O287, O288, O289, O290, O291, O292, O293, O294, O295, O296, O297, O298, O299, O300, O301, O302, O303, O304, O305, O306, O307, O308, O309, O310, O311, O312, O313, O314, O315, O316, O317, O318, O319, O320, O321, O322, O323, O324, O325, O326, O327, O328, O329, O330, O331, O332, O333, O334, O335, O336, O337, O338, O339, O340, O341, O342, O343, O344, O345, O346, O347, O348, O349, O350, O351, O352, O353, O354, O355, O356, O357, O358, O359, O360, O361, O362, O363, O364, O365, O366, O367, O368, O369, O370, O371, O372, O373, O374, O375, O376, O377, O378, O379, O380, O381, O382, O383, O384, O385, O386, O387, O388, O389, O390, O391, O392, O393, O394, O395, O396, O397, O398, O399, O400, O401, O402, O403, O404, O405, O406, O407, O408, O409, O410, O411, O412, O413, O414, O415, O416, O417, O418, O419, O420, O421, O422, O423, O424, O425, O426, O427, O428, O429, O430, O431, O432, O433, O434, O435, O436, O437, O438, O439, O440, O441, O442, O443, O444, O445, O446, O447, O448, O449, O450, O451, O452, O453, O454, O455, O456, O457, O458, O459, O460, O461, O462, O463, O464, O465, O466, O467, O468, O469, O470, O471, O472, O473, O474, O475, O476, O477, O478, O479, O480, O481, O482, O483, O484, O485, O486, O487, O488, O489, O490, O491, O492, O493, O494, O495, O496, O497, O498, O499, O500, O501, O502, O503, O504, O505, O506, O507, O508, O509, O510, O511, O512, O513, O514, O515, O516, O517, O518, O519, O520, O521, O522, O523, O524, O525, O526, O527, O528, O529, O530, O531, O532, O533, O534, O535, O536, O537, O538, O539, O540, O541, O542, O543, O544, O545, O546, O547, O548, O549, O550, O551, O552, O553, O554, O555, O556, O557, O558, O559, O560, O561, O562, O563, O564, O565, O566, O567, O568, O569, O570, O571, O572, O573, O574, O575, O576, O577, O578, O579, O580, O581, O582, O583, O584, O585, O586, O587, O588, O589, O590, O591, O592, O593, O594, O595, O596, O597, O598, O599, O600, O601, O602, O603, O604, O605, O606, O607, O608, O609, O610, O611, O612, O613, O614, O615, O616, O617, O618, O619, O620, O621, O622, O623, O624, O625, O626, O627, O628, O629, O630, O631, O632, O633, O634, O635, O636, O637, O638, O639, O640, O641, O642, O643, O644, O645, O646, O647, O648, O649, O650, O651, O652, O653, O654, O655, O656, O657, O658, O659, O660, O661, O662, O663, O664, O665, O666, O667, O668, O669, O670, O671, O672, O673, O674, O675, O676, O677, O678, O679, O680, O681, O682, O683, O684, O685, O686, O687, O688, O689, O690, O691, O692, O693, O694, O695, O696, O697, O698, O699, O700, O701, O702, O703, O704, O705, O706, O707, O708, O709, O710, O711, O712, O713, O714, O715, O716, O717, O718, O719, O720, O721, O722, O723, O724, O725, O726, O727, O728, O729, O730, O731, O732, O733, O734, O735, O736, O737, O738, O739, O740, O741, O742, O743, O744, O745, O746, O747, O748, O749, O750, O751, O752, O753, O754, O755, O756, O757, O758, O759, O760, O761, O762, O763, O764, O765, O766, O767, O768, O769, O770, O771, O772, O773, O774, O775, O776, O777, O778, O779, O780, O781, O782, O783, O784, O785, O786, O787, O788, O789, O790, O791, O792, O793, O794, O795, O796, O797, O798, O799, O800, O801, O802, O803, O804, O805, O806, O807, O808, O809, O810, O811, O812, O813, O814, O815, O816, O817, O818, O819, O820, O821, O822, O823, O824, O825, O826, O827, O828, O829, O830, O831, O832, O833, O834, O835, O836, O837, O838, O839, O840, O841, O842, O843, O844, O845, O846, O847, O848, O849, O850, O851, O852, O853, O854, O855, O856, O857, O858, O859, O860, O861, O862, O863, O864, O865, O866, O867, O868, O869, O870, O871, O872, O873, O874, O875, O876, O877, O878, O879, O880, O881, O882, O883, O884, O885, O886, O887, O888, O889, O890, O891, O892, O893, O894, O895, O896, O897, O898, O899, O900, O901, O902, O903, O904, O905, O906, O907, O908, O909, O910, O911, O912, O913, O914, O915, O916, O917, O918, O919, O920, O921, O922, O923, O924, O925, O926, O927, O928, O929, O930, O931, O932, O933, O934, O935, O936, O937, O938, O939, O940, O941, O942, O943, O944, O945, O946, O947, O948, O949, O950, O951, O952, O953, O954, O955, O956, O957, O958, O959, O960, O961, O962, O963, O964, O965, O966, O967, O968, O969, O970, O971, O972, O973, O974, O975, O976, O977, O978, O979, O980, O981, O982, O983, O984, O985, O986, O987, O988, O989, O990, O991, O992, O993, O994, O995, O996, O997, O998, O999, O1000, O1001, O1002, O1003, O1004, O1005, O1006, O1007, O1008, O1009, O1010, O1011, O1012, O1013, O1014, O1015, O1016, O1017, O1018, O1019, O1020, O1021, O1022, O1023, O1024, O1025, O1026, O1027, O1028, O1029, O1030, O1031, O1032, O1033, O1034, O1035, O1036, O1037, O1038, O1039, O1040, O1041, O1042, O1043, O1044, O1045, O1046, O1047, O1048, O1049, O1050, O1051, O1052, O1053, O1054, O1055, O1056, O1057, O1058, O1059, O1060, O1061, O1062, O1063, O1064, O1065, O1066, O1067, O1068, O1069, O1070, O1071, O1072, O1073, O1074, O1075, O1076, O1077, O1078, O1079, O1080, O1081, O1082, O1083, O1084, O1085, O1086, O1087, O1088, O1089, O1090, O1091, O1092, O1093, O1094, O1095, O1096, O1097, O1098, O1099, O1100, O1101, O1102, O1103, O1104, O1105, O1106, O1107, O1108, O1109, O1110, O1111, O1112, O1113, O1114, O1115, O1116, O1117, O1118, O1119, O1120, O1121, O1122, O1123, O1124, O1125, O1126, O1127, O1128, O1129, O1130, O1131, O1132, O1133, O1134, O1135, O1136, O1137, O1138, O1139, O1140, O1141, O1142, O1143, O1144, O1145, O1146, O1147, O1148, O1149, O1150, O1151, O1152, O1153, O1154, O1155, O1156, O1157, O1158, O1159, O1160, O1161, O1162, O1163, O1164, O1165, O1166, O1167, O1168, O1169, O1170, O1171, O1172, O1173, O1174, O1175, O1176, O1177, O1178, O1179, O1180, O1181, O1182, O1183, O1184, O1185, O1186, O1187, O1188, O1189, O1190, O1191, O1192, O1193, O1194, O1195, O1196, O1197, O1198, O1199, O1200, O1201, O1202, O1203, O1204, O1205, O1206, O1207, O1208, O1209, O1210, O1211, O1212, O1213, O1214, O1215, O1216, O1217, O1218, O1219, O1220, O1221, O1222, O1223, O1224, O1225, O1226, O1227, O1228, O1229, O1230, O1231, O1232, O1233, O1234, O1235, O1236, O1237, O1238, O1239, O1240, O1241, O1242, O1243, O1244, O1245, O1246, O1247, O1248, O1249, O1250, O1251, O1252, O1253, O1254, O1255, O1256, O1257, O1258, O1259, O1260, O1261, O1262, O1263, O1264, O1265, O1266, O1267, O1268, O1269, O1270, O1271, O1272, O1273, O1274, O1275, O1276, O1277, O1278, O1279, O1280, O1281, O1282, O1283, O1284, O1285, O1286, O1287, O1288, O1289, O1290, O1291, O1292, O1293, O1294, O1295, O1296, O1297, O1298, O1299, O1300, O1301, O1302, O1303, O1304, O1305, O1306, O1307, O1308, O1309, O1310, O1311, O1312, O1313, O1314, O1315, O1316, O1317, O1318, O1319, O1320, O1321, O1322, O1323, O1324, O1325, O1326, O1327, O1328, O1329, O1330, O1331, O1332, O1333, O1334, O1335, O1336, O1337, O1338, O1339, O1340, O1341, O1342, O1343, O1344, O1345, O1346, O1347, O1348, O1349, O1350, O1351, O1352, O1353, O1354, O1355, O1356, O1357, O1358, O1359, O1360, O1361, O1362, O1363, O1364, O1365, O1366, O1367, O1368, O1369, O1370, O1371, O1372, O1373, O1374, O1375, O1376, O1377, O1378, O1379, O1380, O1381, O1382, O1383, O1384, O1385, O1386, O1387, O1388, O1389, O1390, O1391, O1392, O1393, O1394, O1395, O1396, O1397, O1398, O1399, O1400, O1401, O1402, O1403, O1404, O1405, O1406, O1407, O1408, O1409, O1410, O1411, O1412, O1413, O1414, O1415, O1416, O1417, O1418, O1419, O1420, O1421, O1422, O1423, O1424, O1425, O1426, O1427, O1428, O1429, O1430, O1431, O1432, O1433, O1434, O1435, O1436, O1437, O1438, O1439, O1440, O1441, O1442, O1443, O1444, O1445, O1446, O1447, O1448, O1449, O1450, O1451, O1452, O1453, O1454, O1455, O1456, O1457, O1458, O1459, O1460, O1461, O1462, O1463, O1464, O1465, O1466, O1467, O1468, O1469, O1470, O1471, O1472, O1473, O1474, O1475, O1476, O1477, O1478, O1479, O1480, O1481, O1482, O1483, O1484, O1485, O1486, O1487, O1488, O1489, O1490, O1491, O1492, O1493, O1494, O1495, O1496, O1497, O1498, O1499, O1500, O1501, O1502, O1503, O1504, O1505, O1506, O1507, O1508, O1509, O1510, O1511, O1512, O1513, O1514, O1515, O1516, O1517, O1518, O1519, O1520, O1521, O1522, O1523, O1524, O1525, O1526, O1527, O1528, O1529, O1530, O1531, O1532, O1533, O1534, O1535, O1536, O1537, O1538, O1539, O1540, O1541, O1542, O1543, O1544, O1545, O1546, O1547, O1548, O1549, O1550, O1551, O1552, O1553, O1554, O1555, O1556, O1557, O1558, O1559, O1560, O1561, O1562, O1563, O1564, O1565, O1566, O1567, O1568, O1569, O1570, O1571, O1572, O1573, O1574, O1575, O1576, O1577, O1578, O1579, O1580, O1581, O1582, O1583, O1584, O1585, O1586, O1587, O1588, O1589, O1590, O1591, O1592, O1593, O1594, O1595, O1596, O1597, O1598, O1599, O1600, O1601, O1602, O1603, O1604, O1605, O1606, O1607, O1608, O1609, O1610, O1611, O1612, O1613, O1614, O1615, O1616, O1617, O1618, O1619, O1620, O1621, O1622, O1623, O1624, O1625, O1626, O1627, O1628, O1629, O1630, O1631, O1632, O1633;
  wire W1214, W1230, W2842, W1224, W2846, W1221, W2851, W2855, W1215, W1213, W2863, W1207, W1200, W2871, W1193, W2884, W1264, W1255, W1253, W1252, W1251, W1249, W1246, W2823, W1244, W2829, W1238, W1237, W1236, W2834, W1122, W1144, W1143, W1142, W2921, W1137, W1134, W1130, W2937, W1125, W2939, W1147, W2943, W2945, W1114, W1112, W2956, W1107, W2885, W2893, W1181, W1180, W1178, W1175, W1174, W1171, W1169, W1268, W1167, W1166, W1165, W1163, W1160, W1159, W1153, W1151, W1149, W1364, W1378, W2702, W1375, W1374, W2705, W1372, W1371, W1370, W1369, W2709, W2714, W1359, W1357, W1356, W1354, W1353, W2721, W1351, W2666, W2646, W2651, W1416, W2654, W1411, W1410, W1349, W2674, W2680, W2684, W1387, W2689, W1307, W1306, W2773, W2779, W1296, W1294, W2781, W1290, W2786, W2767, W2791, W1283, W2802, W1275, W1273, W1272, W1271, W2745, W1346, W1344, W2737, W1333, W1332, W1330, W2741, W2957, W1326, W1321, W2753, W2761, W2765, W2766, W3196, W906, W3190, W901, W899, W896, W893, W892, W911, W887, W3213, W882, W880, W876, W3132, W3140, W946, W3144, W942, W940, W939, W928, W925, W922, W831, W829, W827, W825, W824, W822, W819, W818, W3272, W811, W809, W808, W3279, W805, W855, W3221, W3225, W870, W868, W864, W863, W862, W861, W856, W958, W852, W845, W843, W842, W841, W840, W839, W1069, W1068, W1066, W1062, W1057, W3008, W3034, W1042, W3043, W1038, W1035, W1034, W2958, W1104, W2959, W1102, W1101, W2961, W1097, W1096, W2973, W1032, W1089, W2978, W2985, W2988, W2993, W1078, W1072, W3007, W972, W992, W986, W3104, W982, W3107, W980, W3108, W971, W970, W967, W3123, W963, W962, W960, W959, W1014, W3050, W3052, W3053, W1024, W1022, W3060, W1016, W1013, W3077, W3080, W1003, W998, W994, W1848, W2212, W1838, W2223, W2210, W1824, W2238, W2239, W2241, W2242, W2246, W2185, W1886, W1884, W1883, W1881, W1880, W1877, W1875, W1810, W2195, W1865, W1864, W2196, W2202, W1856, W1855, W1854, W2206, W2320, W1759, W2304, W1757, W2309, W1752, W1751, W2317, W2318, W1745, W1742, W1741, W1740, W2323, W2325, W1736, W1734, W1733, W1786, W2257, W1799, W1798, W2268, W1792, W1790, W2271, W1788, W1783, W1781, W1780, W1778, W1767, W1980, W2066, W2069, W1995, W1993, W2072, W2074, W1989, W2077, W2081, W1983, W2087, W2091, W1975, W2092, W2093, W1970, W2100, W2101, W1966, W2018, W2034, W2035, W2036, W2031, W2027, W2044, W2025, W2023, W2048, W2104, W2017, W2050, W2015, W2014, W2051, W2054, W2056, W2006, W1907, W2138, W1922, W2146, W2148, W2150, W2157, W1909, W1925, W2159, W1904, W2165, W1894, W2171, W1890, W1946, W2109, W2110, W1956, W1955, W2117, W2119, W2121, W1730, W2123, W1943, W2129, W1934, W1931, W2134, W1541, W2517, W1533, W1531, W2529, W1528, W2534, W1525, W1524, W1523, W1519, W1514, W1513, W2555, W1507, W1506, W1504, W2559, W2560, W1501, W2496, W1576, W2491, W1568, W2494, W2495, W1562, W1500, W1560, W1559, W2497, W2500, W1551, W2507, W2510, W1437, W2623, W1448, W1447, W1445, W1444, W1442, W1440, W1439, W2633, W1435, W1433, W1430, W1428, W2639, W1426, W2642, W1482, W2561, W1498, W1495, W1491, W1490, W1488, W1487, W2577, W1483, W1577, W2583, W1479, W1474, W2598, W2601, W1464, W2611, W2612, W1691, W1684, W2378, W2384, W1677, W1676, W1671, W2392, W1698, W1668, W1664, W2398, W1659, W1658, W2400, W2402, W1655, W1727, W2333, W2336, W1722, W2337, W2339, W1718, W2340, W1714, W1653, W2344, W2345, W2348, W1706, W1702, W1701, W2465, W1616, W1614, W2440, W2449, W2450, W2451, W1600, W2460, W2462, W2466, W1584, W2482, W1578, W1650, W2408, W1645, W1644, W2412, W2421, W1630, W2424, W2426, W1623, W1620, W2436, W184, W486, W185, W187, W483, W482, W481, W188, W189, W194, W196, W197, W3634, W176, W505, W504, W503, W173, W501, W174, W178, W3603, W179, W180, W490, W182, W183, W3663, W205, W206, W3893, W209, W453, W210, W451, W212, W448, W213, W3666, W201, W472, W198, W468, W467, W466, W465, W202, W463, W3650, W456, W142, W3537, W3538, W144, W147, W568, W554, W153, W578, W127, W586, W579, W133, W134, W135, W138, W571, W140, W3583, W523, W521, W520, W517, W530, W171, W514, W511, W510, W172, W507, W541, W154, W156, W544, W158, W159, W160, W218, W539, W537, W534, W532, W531, W260, W346, W339, W268, W271, W329, W272, W274, W275, W356, W366, W365, W3741, W355, W254, W256, W257, W258, W350, W307, W306, W304, W303, W302, W300, W298, W295, W294, W324, W323, W279, W280, W281, W283, W3799, W315, W3802, W310, W230, W3704, W3705, W411, W410, W409, W408, W406, W405, W403, W401, W231, W430, W436, W219, W220, W221, W431, W400, W428, W425, W422, W421, W241, W237, W238, W377, W376, W375, W374, W372, W379, W244, W3735, W245, W246, W248, W388, W399, W398, W397, W396, W233, W390, W3560, W386, W384, W382, W380, W700, W57, W60, W61, W702, W709, W698, W696, W694, W692, W3392, W688, W687, W3360, W724, W45, W721, W3365, W3372, W55, W712, W3375, W710, W56, W85, W668, W666, W665, W84, W80, W658, W655, W654, W87, W3397, W680, W3357, W73, W75, W76, W3416, W670, W775, W782, W781, W10, W779, W13, W15, W774, W773, W772, W768, W3292, W3, W4, W3289, W796, W5, W3290, W3291, W21, W792, W791, W788, W785, W35, W748, W747, W32, W3339, W738, W750, W733, W37, W731, W39, W40, W3356, W757, W3310, W3313, W24, W761, W760, W3322, W25, W693, W756, W754, W3332, W28, W119, W107, W3458, W3489, W103, W635, W629, W3494, W600, W599, W96, W639, W3981, W619, W110, W621, W109, W589, W625, W3978, W3485, W627, W590, W3435, W652, W89, W3442, W90, W653, W3438, W122, W651, W92, W95, W124, W593, W2411, W2065, W2409, W2245, W2064, W2214, W2240, W2259, W2079, W2394, W2396, W2258, W2075, W2251, W2403, W2070, W2194, W3854, W2443, W2232, W2217, W2230, W2438, W2439, W2441, W2442, W2205, W2445, W2446, W2226, W2224, W2043, W2198, W2059, W2200, W2234, W2433, W2434, W2132, W2286, W2331, W2287, W2330, W3886, W2126, W2128, W2280, W2302, W2162, W2161, W2154, W2314, W2160, W2167, W2289, W2327, W2168, W2141, W2143, W2352, W2166, W2290, W2147, W2322, W2094, W2382, W2380, W2269, W2105, W2376, W2375, W2106, W2089, W2260, W2186, W2653, W2390, W2261, W2385, W2354, W2120, W2122, W2369, W2367, W2366, W2272, W2082, W2360, W2357, W3037, W3035, W3031, W3027, W3451, W3022, W3015, W3472, W2992, W2990, W2986, W3088, W3085, W3081, W3072, W3421, W3066, W3432, W3058, W3054, W3047, W3443, W3039, W2909, W2922, W2919, W2918, W3525, W3528, W2915, W2926, W2907, W2906, W2902, W2900, W2967, W3487, W3492, W3414, W3500, W2946, W2938, W2934, W2931, W2930, W3323, W3230, W3226, W3334, W3341, W3344, W3193, W3353, W3264, W3188, W3299, W3245, W3117, W3382, W3139, W3389, W3400, W3187, W3179, W3367, W3162, W2599, W2627, W2624, W2620, W2615, W2606, W2597, W2594, W2588, W2581, W3750, W2575, W2700, W2686, W2662, W2637, W2636, W2505, W2523, W2519, W2518, W2516, W2509, W3793, W2525, W2502, W2489, W2487, W2483, W2471, W2469, W2567, W3755, W2551, W2544, W2542, W3774, W2537, W2535, W2531, W3579, W3580, W3582, W2828, W2827, W2825, W3584, W2822, W2820, W2819, W2818, W2808, W3599, W2804, W2876, W2897, W2891, W2889, W2887, W3562, W2868, W2867, W2864, W3568, W2853, W2724, W2736, W2733, W2728, W2722, W2720, W3668, W2719, W2708, W3609, W2468, W2772, W3633, W2754, W2752, W474, W1335, W459, W462, W464, W469, W1320, W470, W471, W1316, W1315, W1338, W476, W1311, W477, W478, W479, W1303, W1301, W1300, W1297, W485, W487, W447, W1383, W1382, W1381, W440, W1376, W1373, W1367, W1366, W444, W445, W446, W488, W1360, W450, W1355, W452, W455, W1345, W1343, W1341, W1340, W1339, W457, W1209, W525, W1226, W526, W527, W1223, W528, W535, W536, W1217, W1216, W543, W545, W524, W1208, W1205, W1204, W1203, W546, W1198, W1196, W549, W551, W552, W553, W1261, W489, W1281, W1280, W494, W1278, W1277, W1276, W1274, W496, W1265, W497, W498, W1384, W1260, W1258, W502, W1256, W508, W509, W512, W513, W1239, W1235, W516, W1233, W1232, W1508, W325, W327, W1526, W328, W1520, W1518, W331, W336, W1515, W1511, W1529, W341, W1502, W1494, W344, W347, W349, W1489, W351, W352, W354, W358, W1552, W297, W1579, W1573, W1571, W1570, W301, W1567, W309, W1553, W360, W312, W1544, W1543, W1542, W1539, W1538, W317, W1535, W320, W321, W322, W1406, W412, W1422, W1419, W415, W416, W1418, W1417, W1414, W418, W419, W1408, W1424, W1403, W426, W1401, W427, W1397, W1396, W1395, W1394, W1392, W1391, W1390, W1388, W1455, W361, W1473, W362, W1470, W368, W1468, W1461, W1460, W1459, W373, W1458, W1457, W1194, W1454, W381, W387, W389, W391, W1446, W392, W1441, W1429, W404, W407, W931, W705, W706, W949, W708, W941, W938, W936, W715, W934, W933, W716, W932, W953, W717, W930, W929, W722, W723, W727, W921, W920, W728, W916, W730, W912, W908, W683, W995, W993, W991, W673, W675, W987, W985, W677, W679, W981, W682, W978, W977, W734, W974, W685, W686, W689, W690, W965, W964, W695, W961, W697, W699, W703, W954, W784, W765, W850, W766, W847, W846, W776, W835, W834, W778, W828, W826, W854, W823, W787, W815, W794, W795, W797, W799, W810, W807, W806, W804, W800, W907, W739, W902, W900, W897, W894, W891, W741, W890, W742, W889, W885, W749, W751, W883, W879, W755, W872, W871, W758, W866, W860, W764, W1111, W573, W574, W1135, W577, W1132, W1128, W581, W1126, W582, W1120, W587, W1113, W1110, W1109, W588, W1103, W592, W1095, W1093, W595, W1091, W1090, W1087, W555, W1190, W557, W1186, W559, W1179, W561, W562, W605, W1168, W1164, W564, W1158, W565, W1156, W1154, W1150, W1148, W1146, W1145, W1141, W656, W633, W1043, W636, W640, W1030, W644, W1028, W1027, W1026, W645, W647, W648, W1020, W632, W1015, W657, W1010, W1009, W661, W663, W667, W1005, W1001, W999, W997, W996, W615, W1086, W606, W1084, W607, W1081, W1080, W1079, W610, W1077, W1076, W613, W614, W2032, W1074, W1073, W624, W1064, W1060, W1059, W1056, W1055, W1054, W631, W1050, W1048, W1773, W1801, W1796, W139, W1794, W146, W148, W150, W1777, W151, W1802, W1771, W1769, W155, W162, W163, W164, W1762, W1758, W1821, W1846, W1845, W111, W1837, W1831, W1830, W116, W117, W120, W121, W1822, W1756, W125, W1818, W1815, W128, W1809, W1806, W131, W1803, W204, W199, W1708, W1707, W1703, W203, W1696, W1694, W1693, W1690, W1710, W215, W217, W223, W224, W225, W1680, W227, W1731, W1754, W167, W1748, W1747, W1744, W1739, W170, W1737, W1732, W1729, W1728, W177, W1725, W186, W190, W192, W195, W42, W1988, W1987, W19, W22, W1985, W27, W30, W1974, W1969, W1990, W1963, W47, W1954, W1953, W1952, W1949, W51, W1940, W2011, W1, W2, W6, W2028, W8, W2020, W2019, W9, W2012, W11, W1938, W2009, W2007, W14, W2000, W1998, W1991, W1874, W97, W1872, W1871, W98, W1870, W1869, W101, W1889, W102, W104, W1858, W105, W1857, W1852, W106, W1851, W1937, W1932, W1930, W54, W58, W1921, W67, W68, W1916, W293, W1910, W1905, W72, W1902, W78, W82, W1893, W1891, W1636, W1631, W252, W262, W1667, W284, W235, W1670, W263, W1587, W1625, W288, W1593, W232, W1589, W286, W1605, W269, W1591, W1592, W1646, W242, W1638, W1610, W287, W236, W1666, W1586, W1615, W292, W1651, W276, W229, W266, W265, W1678, W1674, W277, W1612, W1652, W259, W290, W1654, W1599, W240, W1618, W1603, W255, W1595, W1624, W289, W1601, W264, W70, W671, W3417, W662, W669, W69, W64, W664, W59, W3404, W326, W684, W62, W53, W270, W52, W3407, W63, W674, W65, W66, W330, W626, W3466, W628, W630, W94, W337, W93, W91, W616, W609, W3481, W611, W99, W340, W338, W617, W618, W622, W623, W267, W334, W83, W79, W50, W77, W646, W335, W3436, W74, W86, W649, W650, W333, W3781, W71, W659, W332, W3452, W634, W88, W637, W660, W638, W641, W642, W643, W3324, W311, W16, W759, W3320, W17, W763, W3314, W746, W20, W743, W745, W18, W752, W753, W299, W786, W789, W793, W3822, W7, W291, W296, W3286, W2033, W424, W767, W308, W770, W771, W12, W3302, W305, W777, W783, W46, W49, W48, W714, W316, W0, W44, W282, W43, W41, W719, W319, W691, W4044, W273, W3387, W704, W720, W318, W3380, W3379, W707, W31, W34, W735, W736, W737, W33, W732, W313, W29, W740, W26, W3343, W23, W285, W38, W3363, W3361, W725, W3359, W726, W314, W729, W36, W3352, W3622, W3621, W169, W168, W484, W480, W3614, W492, W475, W239, W402, W473, W395, W493, W394, W3631, W393, W175, W3587, W247, W506, W3590, W161, W157, W515, W249, W518, W495, W3607, W166, W378, W243, W499, W500, W434, W437, W211, W208, W438, W439, W216, W207, W441, W442, W417, W228, W226, W423, W429, W3685, W432, W222, W433, W461, W193, W458, W3708, W191, W460, W3654, W3870, W181, W414, W443, W3702, W449, W3661, W454, W200, W413, W3521, W114, W113, W112, W584, W585, W572, W123, W3748, W359, W357, W118, W569, W3509, W575, W576, W353, W261, W115, W580, W348, W601, W345, W602, W603, W604, W3490, W598, W608, W343, W342, W3999, W591, W594, W108, W3498, W596, W597, W3952, W538, W540, W251, W542, W149, W370, W145, W369, W547, W143, W548, W519, W522, W152, W529, W533, W371, W3731, W363, W130, W129, W563, W126, W566, W567, W556, W141, W137, W550, W100, W136, W132, W367, W558, W364, W1598, W1585, W2477, W2474, W2473, W2472, W1590, W1594, W1596, W2480, W2455, W2453, W2452, W2448, W1604, W1606, W1609, W1534, W1536, W2520, W1537, W1540, W1545, W1546, W2508, W1548, W1613, W2501, W1555, W2498, W1563, W1564, W1569, W1575, W1581, W1582, W2481, W1669, W1672, W2388, W1665, W2373, W2372, W2370, W1685, W2368, W1686, W1687, W1688, W1692, W1619, W1622, W2432, W2429, W1628, W1629, W1532, W2420, W1634, W1635, W2404, W2401, W2608, W1449, W1450, W2625, W1451, W1452, W1453, W2628, W1462, W2605, W1465, W2603, W1466, W1467, W2600, W1469, W1471, W2593, W1420, W1405, W1407, W1409, W1412, W2659, W2658, W2657, W2656, W2655, W2650, W1421, W1427, W2632, W1443, W1499, W1503, W1505, W2556, W1512, W2548, W2547, W2545, W1516, W2562, W1517, W2538, W1522, W2533, W1527, W2527, W1530, W1472, W2589, W1475, W1476, W1478, W1480, W1481, W2580, W2579, W1695, W1484, W2573, W1497, W2563, W1912, W2152, W2149, W1917, W1919, W1920, W2145, W2144, W2142, W1923, W2139, W1911, W1926, W1927, W1933, W1935, W1942, W1944, W1948, W2116, W1957, W1958, W2175, W2192, W2189, W1876, W2183, W2182, W2179, W2178, W1885, W1887, W2112, W1892, W2170, W1895, W1896, W1897, W1899, W1903, W1906, W2156, W2155, W2055, W2078, W1996, W2067, W2001, W2002, W2003, W2060, W2010, W2080, W2013, W2016, W2022, W2026, W2041, W2029, W2037, W2095, W1960, W1961, W2107, W1965, W2103, W2102, W1967, W2097, W2096, W1973, W1976, W1978, W1979, W2086, W2084, W1982, W1984, W2293, W2311, W2310, W1755, W2306, W2305, W1761, W2301, W2295, W2294, W2292, W2291, W1766, W1770, W1772, W1774, W1775, W1776, W2278, W1779, W1723, W1697, W2351, W2350, W2347, W1712, W1715, W2341, W1716, W1719, W1784, W2335, W2334, W1726, W2324, W1738, W1746, W2316, W2315, W1820, W1823, W2231, W1825, W1829, W1832, W1834, W2222, W1835, W1839, W1842, W1847, W2207, W2203, W1862, W2255, W1787, W2266, W1795, W2263, W2262, W1800, W2254, W2253, W2252, W1805, W2248, W1812, W1814, W1819, W3089, W3084, W1002, W1004, W1006, W1007, W989, W3074, W1012, W1017, W1018, W1019, W1023, W1025, W973, W957, W3129, W3128, W3124, W3120, W966, W968, W969, W3114, W976, W979, W3105, W984, W3099, W988, W3019, W3017, W1061, W1063, W3013, W3011, W1067, W1070, W1071, W3020, W1075, W2997, W2996, W1083, W1085, W3056, W3055, W1029, W3049, W1031, W1036, W1037, W1040, W1041, W3042, W3038, W1045, W1046, W1047, W1049, W1051, W1053, W867, W849, W3243, W3242, W3239, W853, W857, W858, W859, W865, W869, W875, W877, W881, W3214, W884, W821, W802, W803, W3278, W812, W813, W814, W816, W3263, W832, W833, W3254, W836, W837, W838, W844, W3249, W3168, W924, W3165, W926, W927, W3161, W935, W3169, W943, W944, W948, W950, W951, W3137, W952, W955, W3207, W886, W3200, W3198, W895, W903, W2984, W905, W3184, W909, W910, W913, W914, W915, W917, W923, W3170, W1308, W1289, W1292, W1293, W1298, W1299, W2774, W1304, W1305, W1288, W2764, W2763, W1314, W2756, W2755, W1318, W1322, W1269, W1248, W2821, W1250, W2813, W1262, W1263, W1267, W1323, W1270, W1279, W1282, W1285, W1286, W2787, W2691, W1363, W1377, W1379, W1380, W2697, W1362, W1385, W1389, W2678, W2677, W1398, W2673, W1402, W1324, W2747, W1325, W2744, W1329, W1331, W1334, W1337, W2730, W1347, W1348, W1350, W1352, W2717, W1361, W2713, W2927, W1116, W1117, W1118, W1119, W1121, W1124, W1127, W2935, W2933, W1131, W1133, W1115, W1136, W2924, W1138, W2920, W2913, W2911, W1157, W2964, W2979, W2974, W1092, W1094, W1161, W2963, W1098, W1099, W1100, W1105, W1108, W2952, W2950, W2947, W2857, W1212, W1218, W1219, W2850, W1222, W1225, W1210, W1227, W1228, W1234, W2832, W2830, W1240, W2826, W1195, W1162, W1170, W1172, W1176, W1177, W1183, W1185, W1192, W2881, W801, W2873, W1201, W1202, W2861, W2860;

  NOR2X1 G0 (.A1(W349), .A2(W163), .ZN(W1214));
  NOR2X1 G1 (.A1(I157), .A2(W1012), .ZN(W1230));
  NOR2X1 G2 (.A1(W638), .A2(W982), .ZN(O82));
  NOR2X1 G3 (.A1(W1070), .A2(W1650), .ZN(O658));
  NOR2X1 G4 (.A1(W637), .A2(W2084), .ZN(W2842));
  NOR2X1 G5 (.A1(W746), .A2(W2245), .ZN(O663));
  NOR2X1 G6 (.A1(W700), .A2(W338), .ZN(W1224));
  NOR2X1 G7 (.A1(W521), .A2(W1171), .ZN(W2846));
  NOR2X1 G8 (.A1(W850), .A2(W129), .ZN(W1221));
  NOR2X1 G9 (.A1(W1320), .A2(W1459), .ZN(W2851));
  NOR2X1 G10 (.A1(W1160), .A2(W46), .ZN(O668));
  NOR2X1 G11 (.A1(W5), .A2(W443), .ZN(W2855));
  NOR2X1 G12 (.A1(W145), .A2(W696), .ZN(W1215));
  NOR2X1 G13 (.A1(W129), .A2(W1028), .ZN(O83));
  NOR2X1 G14 (.A1(W249), .A2(W519), .ZN(W1213));
  NOR2X1 G15 (.A1(W748), .A2(W454), .ZN(O669));
  NOR2X1 G16 (.A1(W786), .A2(W1715), .ZN(O670));
  NOR2X1 G17 (.A1(W2853), .A2(W270), .ZN(W2863));
  NOR2X1 G18 (.A1(W753), .A2(W339), .ZN(W1207));
  NOR2X1 G19 (.A1(W911), .A2(W273), .ZN(O674));
  NOR2X1 G20 (.A1(W168), .A2(W999), .ZN(W1200));
  NOR2X1 G21 (.A1(W2752), .A2(W2261), .ZN(W2871));
  NOR2X1 G22 (.A1(W2037), .A2(W2579), .ZN(O684));
  NOR2X1 G23 (.A1(W322), .A2(W140), .ZN(W1193));
  NOR2X1 G24 (.A1(I115), .A2(W426), .ZN(W2884));
  NOR2X1 G25 (.A1(W92), .A2(W449), .ZN(O88));
  NOR2X1 G26 (.A1(W2625), .A2(W178), .ZN(O643));
  NOR2X1 G27 (.A1(W256), .A2(W747), .ZN(W1264));
  NOR2X1 G28 (.A1(W56), .A2(W1472), .ZN(O645));
  NOR2X1 G29 (.A1(W1204), .A2(W636), .ZN(O646));
  NOR2X1 G30 (.A1(W1454), .A2(W1142), .ZN(O647));
  NOR2X1 G31 (.A1(W478), .A2(I174), .ZN(O91));
  NOR2X1 G32 (.A1(W641), .A2(W771), .ZN(O90));
  NOR2X1 G33 (.A1(W121), .A2(W366), .ZN(W1255));
  NOR2X1 G34 (.A1(W13), .A2(W175), .ZN(W1253));
  NOR2X1 G35 (.A1(W1096), .A2(W1194), .ZN(W1252));
  NOR2X1 G36 (.A1(W908), .A2(W249), .ZN(W1251));
  NOR2X1 G37 (.A1(W1215), .A2(W95), .ZN(W1249));
  NOR2X1 G38 (.A1(W806), .A2(W805), .ZN(O76));
  NOR2X1 G39 (.A1(W949), .A2(W1009), .ZN(W1246));
  NOR2X1 G40 (.A1(I191), .A2(W632), .ZN(W2823));
  NOR2X1 G41 (.A1(W683), .A2(W70), .ZN(W1244));
  NOR2X1 G42 (.A1(W389), .A2(W173), .ZN(O84));
  NOR2X1 G43 (.A1(W2471), .A2(I51), .ZN(W2829));
  NOR2X1 G44 (.A1(W836), .A2(W1071), .ZN(W1238));
  NOR2X1 G45 (.A1(W257), .A2(W282), .ZN(W1237));
  NOR2X1 G46 (.A1(W846), .A2(W260), .ZN(W1236));
  NOR2X1 G47 (.A1(W1790), .A2(W959), .ZN(W2834));
  NOR2X1 G48 (.A1(W1005), .A2(W390), .ZN(O654));
  NOR2X1 G49 (.A1(W1099), .A2(W2351), .ZN(O655));
  NOR2X1 G50 (.A1(W819), .A2(W1119), .ZN(W1122));
  NOR2X1 G51 (.A1(W1061), .A2(I180), .ZN(W1144));
  NOR2X1 G52 (.A1(W1120), .A2(W952), .ZN(W1143));
  NOR2X1 G53 (.A1(W280), .A2(W994), .ZN(W1142));
  NOR2X1 G54 (.A1(W935), .A2(W1214), .ZN(W2921));
  NOR2X1 G55 (.A1(W418), .A2(W461), .ZN(W1137));
  NOR2X1 G56 (.A1(W2529), .A2(W198), .ZN(O707));
  NOR2X1 G57 (.A1(W6), .A2(W159), .ZN(W1134));
  NOR2X1 G58 (.A1(W137), .A2(W311), .ZN(W1130));
  NOR2X1 G59 (.A1(W417), .A2(W602), .ZN(O65));
  NOR2X1 G60 (.A1(W2646), .A2(W705), .ZN(W2937));
  NOR2X1 G61 (.A1(W1109), .A2(W147), .ZN(W1125));
  NOR2X1 G62 (.A1(W2189), .A2(W294), .ZN(W2939));
  NOR2X1 G63 (.A1(W809), .A2(W66), .ZN(W1147));
  NOR2X1 G64 (.A1(W1026), .A2(W223), .ZN(O711));
  NOR2X1 G65 (.A1(W1426), .A2(W227), .ZN(O712));
  NOR2X1 G66 (.A1(W2655), .A2(W2378), .ZN(W2943));
  NOR2X1 G67 (.A1(W1635), .A2(W1427), .ZN(O714));
  NOR2X1 G68 (.A1(W1180), .A2(I138), .ZN(W2945));
  NOR2X1 G69 (.A1(W631), .A2(W733), .ZN(W1114));
  NOR2X1 G70 (.A1(W1599), .A2(W852), .ZN(O716));
  NOR2X1 G71 (.A1(W72), .A2(W905), .ZN(W1112));
  NOR2X1 G72 (.A1(W673), .A2(W577), .ZN(O720));
  NOR2X1 G73 (.A1(W2314), .A2(W1437), .ZN(W2956));
  NOR2X1 G74 (.A1(W33), .A2(W456), .ZN(W1107));
  NOR2X1 G75 (.A1(W1395), .A2(W1014), .ZN(O695));
  NOR2X1 G76 (.A1(W784), .A2(W1343), .ZN(W2885));
  NOR2X1 G77 (.A1(W1210), .A2(W633), .ZN(O689));
  NOR2X1 G78 (.A1(W2767), .A2(W2421), .ZN(W2893));
  NOR2X1 G79 (.A1(W106), .A2(W1160), .ZN(O71));
  NOR2X1 G80 (.A1(W953), .A2(I38), .ZN(W1181));
  NOR2X1 G81 (.A1(W151), .A2(W342), .ZN(W1180));
  NOR2X1 G82 (.A1(W615), .A2(I17), .ZN(W1178));
  NOR2X1 G83 (.A1(W1005), .A2(W2744), .ZN(O692));
  NOR2X1 G84 (.A1(W127), .A2(W883), .ZN(W1175));
  NOR2X1 G85 (.A1(I178), .A2(W793), .ZN(W1174));
  NOR2X1 G86 (.A1(W444), .A2(W540), .ZN(W1171));
  NOR2X1 G87 (.A1(I98), .A2(W608), .ZN(W1169));
  NOR2X1 G88 (.A1(W275), .A2(W121), .ZN(W1268));
  NOR2X1 G89 (.A1(W19), .A2(W893), .ZN(W1167));
  NOR2X1 G90 (.A1(W349), .A2(W689), .ZN(W1166));
  NOR2X1 G91 (.A1(I31), .A2(W72), .ZN(W1165));
  NOR2X1 G92 (.A1(W831), .A2(I152), .ZN(W1163));
  NOR2X1 G93 (.A1(W2025), .A2(W1029), .ZN(O697));
  NOR2X1 G94 (.A1(W536), .A2(W970), .ZN(W1160));
  NOR2X1 G95 (.A1(W730), .A2(W920), .ZN(W1159));
  NOR2X1 G96 (.A1(W1912), .A2(W1983), .ZN(O700));
  NOR2X1 G97 (.A1(W366), .A2(I86), .ZN(W1153));
  NOR2X1 G98 (.A1(W862), .A2(W371), .ZN(W1151));
  NOR2X1 G99 (.A1(W841), .A2(W786), .ZN(W1149));
  NOR2X1 G100 (.A1(W748), .A2(W186), .ZN(W1364));
  NOR2X1 G101 (.A1(W141), .A2(W186), .ZN(W1378));
  NOR2X1 G102 (.A1(W119), .A2(I44), .ZN(W2702));
  NOR2X1 G103 (.A1(I164), .A2(W451), .ZN(O580));
  NOR2X1 G104 (.A1(W1332), .A2(W348), .ZN(W1375));
  NOR2X1 G105 (.A1(W1235), .A2(W1154), .ZN(W1374));
  NOR2X1 G106 (.A1(W2178), .A2(W372), .ZN(W2705));
  NOR2X1 G107 (.A1(W827), .A2(W608), .ZN(W1372));
  NOR2X1 G108 (.A1(W586), .A2(W661), .ZN(W1371));
  NOR2X1 G109 (.A1(W409), .A2(W1289), .ZN(W1370));
  NOR2X1 G110 (.A1(W304), .A2(W78), .ZN(W1369));
  NOR2X1 G111 (.A1(W871), .A2(W951), .ZN(O582));
  NOR2X1 G112 (.A1(W2183), .A2(W104), .ZN(W2709));
  NOR2X1 G113 (.A1(W135), .A2(I166), .ZN(O574));
  NOR2X1 G114 (.A1(W2347), .A2(W296), .ZN(O583));
  NOR2X1 G115 (.A1(W2117), .A2(I86), .ZN(O585));
  NOR2X1 G116 (.A1(W21), .A2(I188), .ZN(W2714));
  NOR2X1 G117 (.A1(W2600), .A2(W1331), .ZN(O586));
  NOR2X1 G118 (.A1(W261), .A2(W166), .ZN(W1359));
  NOR2X1 G119 (.A1(W1192), .A2(W125), .ZN(W1357));
  NOR2X1 G120 (.A1(W136), .A2(W1177), .ZN(W1356));
  NOR2X1 G121 (.A1(W502), .A2(W1224), .ZN(W1354));
  NOR2X1 G122 (.A1(W1275), .A2(W846), .ZN(W1353));
  NOR2X1 G123 (.A1(W1886), .A2(W1570), .ZN(W2721));
  NOR2X1 G124 (.A1(I184), .A2(W1019), .ZN(W1351));
  NOR2X1 G125 (.A1(W1955), .A2(W2372), .ZN(W2666));
  NOR2X1 G126 (.A1(W709), .A2(W1948), .ZN(W2646));
  NOR2X1 G127 (.A1(W1240), .A2(W977), .ZN(O547));
  NOR2X1 G128 (.A1(W2436), .A2(W591), .ZN(W2651));
  NOR2X1 G129 (.A1(W1298), .A2(I196), .ZN(W1416));
  NOR2X1 G130 (.A1(W504), .A2(W38), .ZN(O117));
  NOR2X1 G131 (.A1(W580), .A2(W2350), .ZN(W2654));
  NOR2X1 G132 (.A1(W421), .A2(W642), .ZN(O116));
  NOR2X1 G133 (.A1(W694), .A2(W908), .ZN(W1411));
  NOR2X1 G134 (.A1(W615), .A2(W1167), .ZN(W1410));
  NOR2X1 G135 (.A1(W124), .A2(W727), .ZN(O552));
  NOR2X1 G136 (.A1(I150), .A2(W2434), .ZN(O554));
  NOR2X1 G137 (.A1(W375), .A2(W957), .ZN(O115));
  NOR2X1 G138 (.A1(W25), .A2(W1275), .ZN(W1349));
  NOR2X1 G139 (.A1(W1895), .A2(W1185), .ZN(O556));
  NOR2X1 G140 (.A1(W2523), .A2(W1540), .ZN(O558));
  NOR2X1 G141 (.A1(W857), .A2(W692), .ZN(W2674));
  NOR2X1 G142 (.A1(W210), .A2(W791), .ZN(W2680));
  NOR2X1 G143 (.A1(W429), .A2(W1064), .ZN(O112));
  NOR2X1 G144 (.A1(W1348), .A2(W2054), .ZN(W2684));
  NOR2X1 G145 (.A1(W266), .A2(W716), .ZN(W1387));
  NOR2X1 G146 (.A1(W196), .A2(W462), .ZN(O111));
  NOR2X1 G147 (.A1(W294), .A2(W2404), .ZN(W2689));
  NOR2X1 G148 (.A1(W2424), .A2(W330), .ZN(O570));
  NOR2X1 G149 (.A1(W640), .A2(W1506), .ZN(O573));
  NOR2X1 G150 (.A1(I164), .A2(W2074), .ZN(O626));
  NOR2X1 G151 (.A1(W160), .A2(W235), .ZN(W1307));
  NOR2X1 G152 (.A1(W929), .A2(W338), .ZN(W1306));
  NOR2X1 G153 (.A1(W19), .A2(W216), .ZN(O614));
  NOR2X1 G154 (.A1(W2445), .A2(W914), .ZN(W2773));
  NOR2X1 G155 (.A1(W2678), .A2(W2581), .ZN(W2779));
  NOR2X1 G156 (.A1(I81), .A2(W310), .ZN(W1296));
  NOR2X1 G157 (.A1(W15), .A2(I2), .ZN(W1294));
  NOR2X1 G158 (.A1(W1902), .A2(W2589), .ZN(W2781));
  NOR2X1 G159 (.A1(W2755), .A2(W1273), .ZN(O623));
  NOR2X1 G160 (.A1(W2507), .A2(W1757), .ZN(O624));
  NOR2X1 G161 (.A1(W359), .A2(W116), .ZN(W1290));
  NOR2X1 G162 (.A1(W1917), .A2(W2087), .ZN(W2786));
  NOR2X1 G163 (.A1(W2646), .A2(W2202), .ZN(W2767));
  NOR2X1 G164 (.A1(W908), .A2(W2680), .ZN(W2791));
  NOR2X1 G165 (.A1(W1054), .A2(W763), .ZN(W1283));
  NOR2X1 G166 (.A1(W1667), .A2(W1426), .ZN(O634));
  NOR2X1 G167 (.A1(W589), .A2(W601), .ZN(O637));
  NOR2X1 G168 (.A1(W2451), .A2(W329), .ZN(O638));
  NOR2X1 G169 (.A1(W458), .A2(W1646), .ZN(W2802));
  NOR2X1 G170 (.A1(W673), .A2(W403), .ZN(W1275));
  NOR2X1 G171 (.A1(W350), .A2(W140), .ZN(W1273));
  NOR2X1 G172 (.A1(W832), .A2(I170), .ZN(W1272));
  NOR2X1 G173 (.A1(W531), .A2(W446), .ZN(W1271));
  NOR2X1 G174 (.A1(W885), .A2(W2501), .ZN(O640));
  NOR2X1 G175 (.A1(W1441), .A2(W473), .ZN(W2745));
  NOR2X1 G176 (.A1(W2271), .A2(W1984), .ZN(O589));
  NOR2X1 G177 (.A1(W333), .A2(W237), .ZN(W1346));
  NOR2X1 G178 (.A1(W417), .A2(W717), .ZN(W1344));
  NOR2X1 G179 (.A1(W1921), .A2(W1548), .ZN(O592));
  NOR2X1 G180 (.A1(W2102), .A2(W1845), .ZN(O597));
  NOR2X1 G181 (.A1(I148), .A2(W1183), .ZN(O106));
  NOR2X1 G182 (.A1(W485), .A2(W698), .ZN(W2737));
  NOR2X1 G183 (.A1(W1113), .A2(W483), .ZN(W1333));
  NOR2X1 G184 (.A1(W928), .A2(W228), .ZN(W1332));
  NOR2X1 G185 (.A1(W1091), .A2(W624), .ZN(W1330));
  NOR2X1 G186 (.A1(W2100), .A2(W2192), .ZN(W2741));
  NOR2X1 G187 (.A1(W1007), .A2(W1084), .ZN(O602));
  NOR2X1 G188 (.A1(I130), .A2(W434), .ZN(W2957));
  NOR2X1 G189 (.A1(W381), .A2(W1224), .ZN(W1326));
  NOR2X1 G190 (.A1(W1109), .A2(W197), .ZN(O603));
  NOR2X1 G191 (.A1(I182), .A2(I192), .ZN(W1321));
  NOR2X1 G192 (.A1(W1715), .A2(W231), .ZN(W2753));
  NOR2X1 G193 (.A1(W367), .A2(W2489), .ZN(O609));
  NOR2X1 G194 (.A1(W1382), .A2(W2186), .ZN(O610));
  NOR2X1 G195 (.A1(W2055), .A2(W2059), .ZN(O611));
  NOR2X1 G196 (.A1(W267), .A2(W1253), .ZN(O101));
  NOR2X1 G197 (.A1(W222), .A2(W402), .ZN(W2761));
  NOR2X1 G198 (.A1(W1832), .A2(W107), .ZN(W2765));
  NOR2X1 G199 (.A1(W2473), .A2(W1874), .ZN(W2766));
  NOR2X1 G200 (.A1(W1078), .A2(W2195), .ZN(W3196));
  NOR2X1 G201 (.A1(W3072), .A2(W1163), .ZN(O862));
  NOR2X1 G202 (.A1(W172), .A2(W1131), .ZN(O865));
  NOR2X1 G203 (.A1(W437), .A2(I44), .ZN(O866));
  NOR2X1 G204 (.A1(I166), .A2(I154), .ZN(W906));
  NOR2X1 G205 (.A1(W2252), .A2(W3074), .ZN(W3190));
  NOR2X1 G206 (.A1(W782), .A2(W358), .ZN(W901));
  NOR2X1 G207 (.A1(W960), .A2(W2573), .ZN(O869));
  NOR2X1 G208 (.A1(W123), .A2(W476), .ZN(W899));
  NOR2X1 G209 (.A1(W117), .A2(W469), .ZN(W896));
  NOR2X1 G210 (.A1(W863), .A2(W2367), .ZN(O871));
  NOR2X1 G211 (.A1(W536), .A2(W288), .ZN(W893));
  NOR2X1 G212 (.A1(W775), .A2(I112), .ZN(W892));
  NOR2X1 G213 (.A1(W557), .A2(W624), .ZN(W911));
  NOR2X1 G214 (.A1(W2611), .A2(W1304), .ZN(O874));
  NOR2X1 G215 (.A1(W1330), .A2(W109), .ZN(O875));
  NOR2X1 G216 (.A1(W1967), .A2(W2495), .ZN(O876));
  NOR2X1 G217 (.A1(I71), .A2(W724), .ZN(W887));
  NOR2X1 G218 (.A1(W1179), .A2(W976), .ZN(O885));
  NOR2X1 G219 (.A1(W113), .A2(W1518), .ZN(W3213));
  NOR2X1 G220 (.A1(W378), .A2(W770), .ZN(W882));
  NOR2X1 G221 (.A1(W333), .A2(W864), .ZN(W880));
  NOR2X1 G222 (.A1(I176), .A2(W267), .ZN(O38));
  NOR2X1 G223 (.A1(W2016), .A2(W739), .ZN(O888));
  NOR2X1 G224 (.A1(W564), .A2(W585), .ZN(W876));
  NOR2X1 G225 (.A1(W1801), .A2(W938), .ZN(O837));
  NOR2X1 G226 (.A1(W145), .A2(W2823), .ZN(W3132));
  NOR2X1 G227 (.A1(W367), .A2(W1164), .ZN(O826));
  NOR2X1 G228 (.A1(W215), .A2(W949), .ZN(O827));
  NOR2X1 G229 (.A1(W1569), .A2(W2198), .ZN(W3140));
  NOR2X1 G230 (.A1(W2673), .A2(W334), .ZN(O831));
  NOR2X1 G231 (.A1(I56), .A2(W386), .ZN(O46));
  NOR2X1 G232 (.A1(W427), .A2(W114), .ZN(W946));
  NOR2X1 G233 (.A1(W302), .A2(W484), .ZN(W3144));
  NOR2X1 G234 (.A1(W939), .A2(W2161), .ZN(O835));
  NOR2X1 G235 (.A1(W355), .A2(W868), .ZN(W942));
  NOR2X1 G236 (.A1(W369), .A2(W79), .ZN(W940));
  NOR2X1 G237 (.A1(W511), .A2(W193), .ZN(W939));
  NOR2X1 G238 (.A1(W823), .A2(W2251), .ZN(O889));
  NOR2X1 G239 (.A1(W2317), .A2(W893), .ZN(O843));
  NOR2X1 G240 (.A1(W2196), .A2(W1668), .ZN(O845));
  NOR2X1 G241 (.A1(W1402), .A2(W532), .ZN(O849));
  NOR2X1 G242 (.A1(W897), .A2(W778), .ZN(W928));
  NOR2X1 G243 (.A1(W707), .A2(W416), .ZN(W925));
  NOR2X1 G244 (.A1(W720), .A2(I104), .ZN(W922));
  NOR2X1 G245 (.A1(W54), .A2(W1067), .ZN(O855));
  NOR2X1 G246 (.A1(I62), .A2(W496), .ZN(O43));
  NOR2X1 G247 (.A1(W773), .A2(W120), .ZN(O42));
  NOR2X1 G248 (.A1(W687), .A2(W122), .ZN(O859));
  NOR2X1 G249 (.A1(W2747), .A2(W365), .ZN(O861));
  NOR2X1 G250 (.A1(I5), .A2(W144), .ZN(O31));
  NOR2X1 G251 (.A1(W1780), .A2(W6), .ZN(O915));
  NOR2X1 G252 (.A1(W2029), .A2(W722), .ZN(O917));
  NOR2X1 G253 (.A1(W2159), .A2(W899), .ZN(O920));
  NOR2X1 G254 (.A1(W235), .A2(W0), .ZN(W831));
  NOR2X1 G255 (.A1(I158), .A2(I172), .ZN(W829));
  NOR2X1 G256 (.A1(W473), .A2(W477), .ZN(W827));
  NOR2X1 G257 (.A1(W204), .A2(I145), .ZN(W825));
  NOR2X1 G258 (.A1(W600), .A2(W239), .ZN(W824));
  NOR2X1 G259 (.A1(W532), .A2(W249), .ZN(W822));
  NOR2X1 G260 (.A1(W1133), .A2(W64), .ZN(O925));
  NOR2X1 G261 (.A1(W588), .A2(W328), .ZN(W819));
  NOR2X1 G262 (.A1(W596), .A2(W552), .ZN(W818));
  NOR2X1 G263 (.A1(W1411), .A2(W1568), .ZN(O913));
  NOR2X1 G264 (.A1(W2138), .A2(W2119), .ZN(O927));
  NOR2X1 G265 (.A1(W2451), .A2(W2330), .ZN(O928));
  NOR2X1 G266 (.A1(W811), .A2(W2483), .ZN(W3272));
  NOR2X1 G267 (.A1(W1616), .A2(W2376), .ZN(O932));
  NOR2X1 G268 (.A1(W273), .A2(W685), .ZN(W811));
  NOR2X1 G269 (.A1(W2747), .A2(W65), .ZN(O934));
  NOR2X1 G270 (.A1(W473), .A2(W511), .ZN(W809));
  NOR2X1 G271 (.A1(W543), .A2(W12), .ZN(W808));
  NOR2X1 G272 (.A1(W1578), .A2(W1728), .ZN(W3279));
  NOR2X1 G273 (.A1(W639), .A2(W264), .ZN(W805));
  NOR2X1 G274 (.A1(W2067), .A2(W1418), .ZN(O937));
  NOR2X1 G275 (.A1(W52), .A2(W59), .ZN(W855));
  NOR2X1 G276 (.A1(W1919), .A2(I174), .ZN(W3221));
  NOR2X1 G277 (.A1(W2561), .A2(W266), .ZN(W3225));
  NOR2X1 G278 (.A1(W742), .A2(I74), .ZN(W870));
  NOR2X1 G279 (.A1(W436), .A2(W635), .ZN(W868));
  NOR2X1 G280 (.A1(I32), .A2(W569), .ZN(W864));
  NOR2X1 G281 (.A1(W800), .A2(W609), .ZN(W863));
  NOR2X1 G282 (.A1(W17), .A2(W747), .ZN(W862));
  NOR2X1 G283 (.A1(W471), .A2(W470), .ZN(W861));
  NOR2X1 G284 (.A1(I79), .A2(W1385), .ZN(O900));
  NOR2X1 G285 (.A1(W1872), .A2(W1494), .ZN(O902));
  NOR2X1 G286 (.A1(W980), .A2(W2112), .ZN(O903));
  NOR2X1 G287 (.A1(I197), .A2(W114), .ZN(W856));
  NOR2X1 G288 (.A1(W509), .A2(W630), .ZN(W958));
  NOR2X1 G289 (.A1(W2700), .A2(W3077), .ZN(O904));
  NOR2X1 G290 (.A1(W805), .A2(W99), .ZN(W852));
  NOR2X1 G291 (.A1(W542), .A2(W1112), .ZN(O906));
  NOR2X1 G292 (.A1(W2248), .A2(W2722), .ZN(O907));
  NOR2X1 G293 (.A1(W3108), .A2(W936), .ZN(O911));
  NOR2X1 G294 (.A1(W27), .A2(W47), .ZN(W845));
  NOR2X1 G295 (.A1(W301), .A2(W590), .ZN(W843));
  NOR2X1 G296 (.A1(W761), .A2(W210), .ZN(W842));
  NOR2X1 G297 (.A1(I84), .A2(W717), .ZN(W841));
  NOR2X1 G298 (.A1(I169), .A2(W213), .ZN(W840));
  NOR2X1 G299 (.A1(W538), .A2(W313), .ZN(W839));
  NOR2X1 G300 (.A1(W2765), .A2(W2963), .ZN(O762));
  NOR2X1 G301 (.A1(W179), .A2(W399), .ZN(W1069));
  NOR2X1 G302 (.A1(W844), .A2(I78), .ZN(W1068));
  NOR2X1 G303 (.A1(W1668), .A2(W1405), .ZN(O751));
  NOR2X1 G304 (.A1(W759), .A2(W770), .ZN(W1066));
  NOR2X1 G305 (.A1(W29), .A2(W720), .ZN(O60));
  NOR2X1 G306 (.A1(W2182), .A2(W2633), .ZN(O754));
  NOR2X1 G307 (.A1(W942), .A2(W526), .ZN(W1062));
  NOR2X1 G308 (.A1(W2662), .A2(W1670), .ZN(O755));
  NOR2X1 G309 (.A1(W351), .A2(W21), .ZN(O758));
  NOR2X1 G310 (.A1(W115), .A2(W870), .ZN(W1057));
  NOR2X1 G311 (.A1(W549), .A2(W1778), .ZN(O760));
  NOR2X1 G312 (.A1(W293), .A2(W495), .ZN(O58));
  NOR2X1 G313 (.A1(W1581), .A2(W825), .ZN(W3008));
  NOR2X1 G314 (.A1(W1592), .A2(W1103), .ZN(O765));
  NOR2X1 G315 (.A1(W2598), .A2(W883), .ZN(W3034));
  NOR2X1 G316 (.A1(W490), .A2(W544), .ZN(O57));
  NOR2X1 G317 (.A1(W586), .A2(W752), .ZN(W1042));
  NOR2X1 G318 (.A1(W1824), .A2(W1830), .ZN(W3043));
  NOR2X1 G319 (.A1(W2915), .A2(W1726), .ZN(O770));
  NOR2X1 G320 (.A1(W164), .A2(W2873), .ZN(O771));
  NOR2X1 G321 (.A1(W174), .A2(W595), .ZN(W1038));
  NOR2X1 G322 (.A1(W56), .A2(W314), .ZN(W1035));
  NOR2X1 G323 (.A1(I147), .A2(I9), .ZN(W1034));
  NOR2X1 G324 (.A1(I46), .A2(I165), .ZN(O55));
  NOR2X1 G325 (.A1(W652), .A2(W797), .ZN(O730));
  NOR2X1 G326 (.A1(W1195), .A2(W2141), .ZN(W2958));
  NOR2X1 G327 (.A1(W218), .A2(W118), .ZN(W1104));
  NOR2X1 G328 (.A1(W496), .A2(W130), .ZN(W2959));
  NOR2X1 G329 (.A1(W307), .A2(W127), .ZN(W1102));
  NOR2X1 G330 (.A1(W691), .A2(W8), .ZN(W1101));
  NOR2X1 G331 (.A1(W451), .A2(W2205), .ZN(W2961));
  NOR2X1 G332 (.A1(I7), .A2(W66), .ZN(W1097));
  NOR2X1 G333 (.A1(W242), .A2(W339), .ZN(W1096));
  NOR2X1 G334 (.A1(W1248), .A2(W2720), .ZN(O723));
  NOR2X1 G335 (.A1(W2651), .A2(W2947), .ZN(O724));
  NOR2X1 G336 (.A1(W2730), .A2(W618), .ZN(O726));
  NOR2X1 G337 (.A1(W1373), .A2(W68), .ZN(W2973));
  NOR2X1 G338 (.A1(I92), .A2(W613), .ZN(W1032));
  NOR2X1 G339 (.A1(W907), .A2(W614), .ZN(W1089));
  NOR2X1 G340 (.A1(I150), .A2(W1268), .ZN(O731));
  NOR2X1 G341 (.A1(W386), .A2(I8), .ZN(W2978));
  NOR2X1 G342 (.A1(W2034), .A2(W616), .ZN(W2985));
  NOR2X1 G343 (.A1(W2013), .A2(W1156), .ZN(W2988));
  NOR2X1 G344 (.A1(W738), .A2(W2440), .ZN(W2993));
  NOR2X1 G345 (.A1(I42), .A2(W511), .ZN(W1078));
  NOR2X1 G346 (.A1(W1814), .A2(W1218), .ZN(O742));
  NOR2X1 G347 (.A1(W2491), .A2(W159), .ZN(O749));
  NOR2X1 G348 (.A1(I42), .A2(I172), .ZN(W1072));
  NOR2X1 G349 (.A1(I84), .A2(W2144), .ZN(W3007));
  NOR2X1 G350 (.A1(W398), .A2(W670), .ZN(W972));
  NOR2X1 G351 (.A1(W326), .A2(W577), .ZN(W992));
  NOR2X1 G352 (.A1(W55), .A2(W1954), .ZN(O798));
  NOR2X1 G353 (.A1(W1414), .A2(W2500), .ZN(O803));
  NOR2X1 G354 (.A1(W2495), .A2(W2056), .ZN(O804));
  NOR2X1 G355 (.A1(W375), .A2(I14), .ZN(W986));
  NOR2X1 G356 (.A1(W1732), .A2(W1917), .ZN(W3104));
  NOR2X1 G357 (.A1(W310), .A2(W534), .ZN(O49));
  NOR2X1 G358 (.A1(I111), .A2(W754), .ZN(W982));
  NOR2X1 G359 (.A1(W659), .A2(W53), .ZN(W3107));
  NOR2X1 G360 (.A1(W889), .A2(W529), .ZN(W980));
  NOR2X1 G361 (.A1(W1051), .A2(W709), .ZN(W3108));
  NOR2X1 G362 (.A1(W1136), .A2(W703), .ZN(O810));
  NOR2X1 G363 (.A1(W1581), .A2(W1802), .ZN(O797));
  NOR2X1 G364 (.A1(W779), .A2(W576), .ZN(W971));
  NOR2X1 G365 (.A1(W651), .A2(W363), .ZN(W970));
  NOR2X1 G366 (.A1(W149), .A2(W1502), .ZN(O816));
  NOR2X1 G367 (.A1(W61), .A2(W653), .ZN(W967));
  NOR2X1 G368 (.A1(W1856), .A2(W19), .ZN(O820));
  NOR2X1 G369 (.A1(W3117), .A2(W147), .ZN(W3123));
  NOR2X1 G370 (.A1(W481), .A2(I116), .ZN(W963));
  NOR2X1 G371 (.A1(W598), .A2(W279), .ZN(W962));
  NOR2X1 G372 (.A1(I111), .A2(W1957), .ZN(O823));
  NOR2X1 G373 (.A1(W650), .A2(W532), .ZN(W960));
  NOR2X1 G374 (.A1(I71), .A2(W215), .ZN(W959));
  NOR2X1 G375 (.A1(W291), .A2(W545), .ZN(W1014));
  NOR2X1 G376 (.A1(W1671), .A2(W1502), .ZN(W3050));
  NOR2X1 G377 (.A1(W638), .A2(W493), .ZN(O774));
  NOR2X1 G378 (.A1(W1417), .A2(W243), .ZN(W3052));
  NOR2X1 G379 (.A1(W1600), .A2(W1739), .ZN(W3053));
  NOR2X1 G380 (.A1(W537), .A2(W37), .ZN(W1024));
  NOR2X1 G381 (.A1(W1005), .A2(W518), .ZN(O776));
  NOR2X1 G382 (.A1(W389), .A2(W488), .ZN(W1022));
  NOR2X1 G383 (.A1(W289), .A2(W26), .ZN(O54));
  NOR2X1 G384 (.A1(W1128), .A2(W761), .ZN(W3060));
  NOR2X1 G385 (.A1(W877), .A2(W1852), .ZN(O777));
  NOR2X1 G386 (.A1(W49), .A2(W86), .ZN(O778));
  NOR2X1 G387 (.A1(W972), .A2(W707), .ZN(W1016));
  NOR2X1 G388 (.A1(W1119), .A2(W167), .ZN(O545));
  NOR2X1 G389 (.A1(W344), .A2(W958), .ZN(W1013));
  NOR2X1 G390 (.A1(W663), .A2(I110), .ZN(O785));
  NOR2X1 G391 (.A1(W302), .A2(W2802), .ZN(O786));
  NOR2X1 G392 (.A1(W209), .A2(W864), .ZN(W3077));
  NOR2X1 G393 (.A1(W1707), .A2(W2325), .ZN(W3080));
  NOR2X1 G394 (.A1(W1542), .A2(W1469), .ZN(O792));
  NOR2X1 G395 (.A1(W884), .A2(W598), .ZN(W1003));
  NOR2X1 G396 (.A1(W147), .A2(W51), .ZN(O51));
  NOR2X1 G397 (.A1(W2755), .A2(W2637), .ZN(O794));
  NOR2X1 G398 (.A1(W138), .A2(I194), .ZN(W998));
  NOR2X1 G399 (.A1(W777), .A2(W324), .ZN(W994));
  NOR2X1 G400 (.A1(W1560), .A2(W47), .ZN(O219));
  NOR2X1 G401 (.A1(W778), .A2(W890), .ZN(O345));
  NOR2X1 G402 (.A1(W957), .A2(W958), .ZN(W1848));
  NOR2X1 G403 (.A1(W1469), .A2(W1176), .ZN(W2212));
  NOR2X1 G404 (.A1(W242), .A2(W824), .ZN(O226));
  NOR2X1 G405 (.A1(W1207), .A2(W1698), .ZN(O225));
  NOR2X1 G406 (.A1(W1446), .A2(W1655), .ZN(O224));
  NOR2X1 G407 (.A1(W1253), .A2(W2001), .ZN(O349));
  NOR2X1 G408 (.A1(W586), .A2(W71), .ZN(W1838));
  NOR2X1 G409 (.A1(W890), .A2(W2064), .ZN(W2223));
  NOR2X1 G410 (.A1(W1512), .A2(W2032), .ZN(O353));
  NOR2X1 G411 (.A1(W1293), .A2(W665), .ZN(O354));
  NOR2X1 G412 (.A1(W1125), .A2(W1076), .ZN(O355));
  NOR2X1 G413 (.A1(W814), .A2(W1954), .ZN(W2210));
  NOR2X1 G414 (.A1(W89), .A2(W1524), .ZN(O218));
  NOR2X1 G415 (.A1(W885), .A2(W1217), .ZN(W1824));
  NOR2X1 G416 (.A1(W302), .A2(W485), .ZN(O357));
  NOR2X1 G417 (.A1(W241), .A2(W2048), .ZN(O359));
  NOR2X1 G418 (.A1(W1161), .A2(W1430), .ZN(W2238));
  NOR2X1 G419 (.A1(W1343), .A2(W593), .ZN(W2239));
  NOR2X1 G420 (.A1(W1538), .A2(I112), .ZN(O217));
  NOR2X1 G421 (.A1(W1622), .A2(W529), .ZN(O216));
  NOR2X1 G422 (.A1(W865), .A2(W712), .ZN(W2241));
  NOR2X1 G423 (.A1(W1449), .A2(W794), .ZN(W2242));
  NOR2X1 G424 (.A1(W1346), .A2(W1802), .ZN(W2246));
  NOR2X1 G425 (.A1(W1066), .A2(W1261), .ZN(W2185));
  NOR2X1 G426 (.A1(W1324), .A2(W557), .ZN(W1886));
  NOR2X1 G427 (.A1(W2097), .A2(W1665), .ZN(O330));
  NOR2X1 G428 (.A1(W449), .A2(W1517), .ZN(W1884));
  NOR2X1 G429 (.A1(W95), .A2(W1615), .ZN(W1883));
  NOR2X1 G430 (.A1(W920), .A2(W422), .ZN(O240));
  NOR2X1 G431 (.A1(W902), .A2(W1015), .ZN(W1881));
  NOR2X1 G432 (.A1(W1802), .A2(W757), .ZN(W1880));
  NOR2X1 G433 (.A1(W1623), .A2(W1085), .ZN(O239));
  NOR2X1 G434 (.A1(W546), .A2(W388), .ZN(O332));
  NOR2X1 G435 (.A1(W1845), .A2(W551), .ZN(W1877));
  NOR2X1 G436 (.A1(W452), .A2(W358), .ZN(O333));
  NOR2X1 G437 (.A1(W227), .A2(I175), .ZN(W1875));
  NOR2X1 G438 (.A1(W209), .A2(W1475), .ZN(W1810));
  NOR2X1 G439 (.A1(W1158), .A2(W185), .ZN(O337));
  NOR2X1 G440 (.A1(W205), .A2(W400), .ZN(W2195));
  NOR2X1 G441 (.A1(W349), .A2(W1537), .ZN(W1865));
  NOR2X1 G442 (.A1(W294), .A2(W686), .ZN(W1864));
  NOR2X1 G443 (.A1(W1373), .A2(W326), .ZN(W2196));
  NOR2X1 G444 (.A1(W9), .A2(W1299), .ZN(W2202));
  NOR2X1 G445 (.A1(W286), .A2(W451), .ZN(O342));
  NOR2X1 G446 (.A1(W909), .A2(W524), .ZN(W1856));
  NOR2X1 G447 (.A1(W840), .A2(W613), .ZN(W1855));
  NOR2X1 G448 (.A1(W258), .A2(W946), .ZN(W1854));
  NOR2X1 G449 (.A1(W754), .A2(W1728), .ZN(W2206));
  NOR2X1 G450 (.A1(W127), .A2(W390), .ZN(W2320));
  NOR2X1 G451 (.A1(W1407), .A2(I156), .ZN(O200));
  NOR2X1 G452 (.A1(W735), .A2(W1529), .ZN(W1759));
  NOR2X1 G453 (.A1(W248), .A2(W299), .ZN(W2304));
  NOR2X1 G454 (.A1(W1278), .A2(W1198), .ZN(W1757));
  NOR2X1 G455 (.A1(W649), .A2(W1181), .ZN(W2309));
  NOR2X1 G456 (.A1(W1480), .A2(W1569), .ZN(O199));
  NOR2X1 G457 (.A1(W1616), .A2(W1239), .ZN(W1752));
  NOR2X1 G458 (.A1(W271), .A2(W635), .ZN(W1751));
  NOR2X1 G459 (.A1(W1736), .A2(W1494), .ZN(O197));
  NOR2X1 G460 (.A1(W343), .A2(W2255), .ZN(W2317));
  NOR2X1 G461 (.A1(W183), .A2(W129), .ZN(W2318));
  NOR2X1 G462 (.A1(W1122), .A2(W895), .ZN(W1745));
  NOR2X1 G463 (.A1(W1279), .A2(W147), .ZN(O388));
  NOR2X1 G464 (.A1(W593), .A2(W1501), .ZN(O394));
  NOR2X1 G465 (.A1(I112), .A2(W1372), .ZN(W1742));
  NOR2X1 G466 (.A1(W1577), .A2(W969), .ZN(W1741));
  NOR2X1 G467 (.A1(W1246), .A2(W137), .ZN(W1740));
  NOR2X1 G468 (.A1(I12), .A2(W2080), .ZN(W2323));
  NOR2X1 G469 (.A1(W1451), .A2(W2031), .ZN(W2325));
  NOR2X1 G470 (.A1(W951), .A2(W753), .ZN(W1736));
  NOR2X1 G471 (.A1(W822), .A2(W1350), .ZN(O195));
  NOR2X1 G472 (.A1(W315), .A2(W1212), .ZN(W1734));
  NOR2X1 G473 (.A1(W680), .A2(W1629), .ZN(W1733));
  NOR2X1 G474 (.A1(W1448), .A2(W62), .ZN(O395));
  NOR2X1 G475 (.A1(W948), .A2(W354), .ZN(W1786));
  NOR2X1 G476 (.A1(W428), .A2(W577), .ZN(O213));
  NOR2X1 G477 (.A1(W1579), .A2(W675), .ZN(O364));
  NOR2X1 G478 (.A1(W1600), .A2(W1077), .ZN(W2257));
  NOR2X1 G479 (.A1(W1567), .A2(W292), .ZN(W1799));
  NOR2X1 G480 (.A1(W1143), .A2(W1285), .ZN(W1798));
  NOR2X1 G481 (.A1(W1769), .A2(W1512), .ZN(O210));
  NOR2X1 G482 (.A1(W1085), .A2(W1124), .ZN(O369));
  NOR2X1 G483 (.A1(W2257), .A2(W1069), .ZN(W2268));
  NOR2X1 G484 (.A1(W774), .A2(W449), .ZN(W1792));
  NOR2X1 G485 (.A1(W995), .A2(W258), .ZN(W1790));
  NOR2X1 G486 (.A1(W128), .A2(W1667), .ZN(W2271));
  NOR2X1 G487 (.A1(W1102), .A2(W1684), .ZN(W1788));
  NOR2X1 G488 (.A1(W139), .A2(W1636), .ZN(O241));
  NOR2X1 G489 (.A1(W844), .A2(W1691), .ZN(O206));
  NOR2X1 G490 (.A1(W354), .A2(W104), .ZN(W1783));
  NOR2X1 G491 (.A1(W1175), .A2(W470), .ZN(O205));
  NOR2X1 G492 (.A1(W776), .A2(W1335), .ZN(W1781));
  NOR2X1 G493 (.A1(W1762), .A2(W543), .ZN(W1780));
  NOR2X1 G494 (.A1(W633), .A2(W1007), .ZN(W1778));
  NOR2X1 G495 (.A1(W1484), .A2(W1783), .ZN(O375));
  NOR2X1 G496 (.A1(W1822), .A2(W1409), .ZN(O380));
  NOR2X1 G497 (.A1(W1349), .A2(W497), .ZN(W1767));
  NOR2X1 G498 (.A1(W690), .A2(W2251), .ZN(O385));
  NOR2X1 G499 (.A1(W446), .A2(W1238), .ZN(O387));
  NOR2X1 G500 (.A1(W1500), .A2(I157), .ZN(W1980));
  NOR2X1 G501 (.A1(W629), .A2(I91), .ZN(O292));
  NOR2X1 G502 (.A1(W768), .A2(W1281), .ZN(W2066));
  NOR2X1 G503 (.A1(W986), .A2(W1099), .ZN(O272));
  NOR2X1 G504 (.A1(I116), .A2(W415), .ZN(W2069));
  NOR2X1 G505 (.A1(I190), .A2(W297), .ZN(W1995));
  NOR2X1 G506 (.A1(W178), .A2(W1935), .ZN(W1993));
  NOR2X1 G507 (.A1(W1051), .A2(W537), .ZN(W2072));
  NOR2X1 G508 (.A1(W839), .A2(W950), .ZN(W2074));
  NOR2X1 G509 (.A1(W102), .A2(W639), .ZN(W1989));
  NOR2X1 G510 (.A1(W859), .A2(W767), .ZN(W2077));
  NOR2X1 G511 (.A1(W1104), .A2(W692), .ZN(W2081));
  NOR2X1 G512 (.A1(I124), .A2(W1507), .ZN(W1983));
  NOR2X1 G513 (.A1(W115), .A2(W559), .ZN(O291));
  NOR2X1 G514 (.A1(W53), .A2(W545), .ZN(W2087));
  NOR2X1 G515 (.A1(W1568), .A2(W2082), .ZN(O300));
  NOR2X1 G516 (.A1(W1476), .A2(W67), .ZN(W2091));
  NOR2X1 G517 (.A1(W781), .A2(W135), .ZN(W1975));
  NOR2X1 G518 (.A1(W1600), .A2(W1794), .ZN(W2092));
  NOR2X1 G519 (.A1(W654), .A2(W2060), .ZN(W2093));
  NOR2X1 G520 (.A1(W1260), .A2(W970), .ZN(W1970));
  NOR2X1 G521 (.A1(W1461), .A2(I14), .ZN(O303));
  NOR2X1 G522 (.A1(W488), .A2(W742), .ZN(W2100));
  NOR2X1 G523 (.A1(W691), .A2(W1664), .ZN(W2101));
  NOR2X1 G524 (.A1(W1498), .A2(W393), .ZN(W1966));
  NOR2X1 G525 (.A1(W273), .A2(W301), .ZN(W2018));
  NOR2X1 G526 (.A1(W1585), .A2(W1985), .ZN(W2034));
  NOR2X1 G527 (.A1(W255), .A2(W1124), .ZN(W2035));
  NOR2X1 G528 (.A1(I18), .A2(W589), .ZN(W2036));
  NOR2X1 G529 (.A1(W200), .A2(W1676), .ZN(W2031));
  NOR2X1 G530 (.A1(W1855), .A2(W1347), .ZN(O281));
  NOR2X1 G531 (.A1(W1222), .A2(W1048), .ZN(W2027));
  NOR2X1 G532 (.A1(W1097), .A2(W237), .ZN(W2044));
  NOR2X1 G533 (.A1(W955), .A2(W938), .ZN(W2025));
  NOR2X1 G534 (.A1(W327), .A2(W193), .ZN(O284));
  NOR2X1 G535 (.A1(W1406), .A2(W760), .ZN(W2023));
  NOR2X1 G536 (.A1(W1693), .A2(W580), .ZN(O276));
  NOR2X1 G537 (.A1(I86), .A2(W1543), .ZN(W2048));
  NOR2X1 G538 (.A1(W1672), .A2(W427), .ZN(W2104));
  NOR2X1 G539 (.A1(W578), .A2(I71), .ZN(W2017));
  NOR2X1 G540 (.A1(W566), .A2(W1710), .ZN(W2050));
  NOR2X1 G541 (.A1(W1869), .A2(W1048), .ZN(W2015));
  NOR2X1 G542 (.A1(I163), .A2(W1591), .ZN(W2014));
  NOR2X1 G543 (.A1(W1378), .A2(W248), .ZN(W2051));
  NOR2X1 G544 (.A1(W139), .A2(W1025), .ZN(W2054));
  NOR2X1 G545 (.A1(W767), .A2(W788), .ZN(W2056));
  NOR2X1 G546 (.A1(W1601), .A2(I161), .ZN(O289));
  NOR2X1 G547 (.A1(W1497), .A2(W1151), .ZN(O275));
  NOR2X1 G548 (.A1(W1634), .A2(W880), .ZN(O290));
  NOR2X1 G549 (.A1(W119), .A2(W74), .ZN(W2006));
  NOR2X1 G550 (.A1(W1822), .A2(W1732), .ZN(W1907));
  NOR2X1 G551 (.A1(W1169), .A2(W1072), .ZN(W2138));
  NOR2X1 G552 (.A1(I48), .A2(W763), .ZN(W1922));
  NOR2X1 G553 (.A1(W2145), .A2(W1214), .ZN(W2146));
  NOR2X1 G554 (.A1(W1350), .A2(W1715), .ZN(O249));
  NOR2X1 G555 (.A1(W1976), .A2(W177), .ZN(W2148));
  NOR2X1 G556 (.A1(W1290), .A2(W1544), .ZN(W2150));
  NOR2X1 G557 (.A1(W88), .A2(W1297), .ZN(O248));
  NOR2X1 G558 (.A1(W1871), .A2(W1883), .ZN(O320));
  NOR2X1 G559 (.A1(W1466), .A2(W1622), .ZN(O246));
  NOR2X1 G560 (.A1(W574), .A2(W800), .ZN(W2157));
  NOR2X1 G561 (.A1(W1540), .A2(W315), .ZN(W1909));
  NOR2X1 G562 (.A1(W1532), .A2(W735), .ZN(O322));
  NOR2X1 G563 (.A1(W1439), .A2(I84), .ZN(W1925));
  NOR2X1 G564 (.A1(W850), .A2(W1146), .ZN(W2159));
  NOR2X1 G565 (.A1(W109), .A2(W1651), .ZN(W1904));
  NOR2X1 G566 (.A1(W272), .A2(W313), .ZN(O244));
  NOR2X1 G567 (.A1(W1835), .A2(W360), .ZN(O324));
  NOR2X1 G568 (.A1(W1344), .A2(W877), .ZN(W2165));
  NOR2X1 G569 (.A1(W1114), .A2(W1168), .ZN(O325));
  NOR2X1 G570 (.A1(W578), .A2(W662), .ZN(W1894));
  NOR2X1 G571 (.A1(W585), .A2(W2010), .ZN(W2171));
  NOR2X1 G572 (.A1(W1369), .A2(W1194), .ZN(O326));
  NOR2X1 G573 (.A1(W1132), .A2(I169), .ZN(O327));
  NOR2X1 G574 (.A1(W726), .A2(W1829), .ZN(W1890));
  NOR2X1 G575 (.A1(W1047), .A2(W1252), .ZN(W1946));
  NOR2X1 G576 (.A1(W924), .A2(W630), .ZN(W2109));
  NOR2X1 G577 (.A1(W1048), .A2(W1264), .ZN(W2110));
  NOR2X1 G578 (.A1(W1022), .A2(W255), .ZN(O260));
  NOR2X1 G579 (.A1(W690), .A2(W611), .ZN(O307));
  NOR2X1 G580 (.A1(I179), .A2(W274), .ZN(W1956));
  NOR2X1 G581 (.A1(W824), .A2(W317), .ZN(W1955));
  NOR2X1 G582 (.A1(W82), .A2(W989), .ZN(W2117));
  NOR2X1 G583 (.A1(W958), .A2(W1369), .ZN(O309));
  NOR2X1 G584 (.A1(W1987), .A2(W1777), .ZN(W2119));
  NOR2X1 G585 (.A1(W368), .A2(W912), .ZN(O259));
  NOR2X1 G586 (.A1(W655), .A2(W1350), .ZN(O258));
  NOR2X1 G587 (.A1(W1447), .A2(W1484), .ZN(W2121));
  NOR2X1 G588 (.A1(W505), .A2(W309), .ZN(W1730));
  NOR2X1 G589 (.A1(W399), .A2(W182), .ZN(W2123));
  NOR2X1 G590 (.A1(W1609), .A2(W1842), .ZN(W1943));
  NOR2X1 G591 (.A1(W1799), .A2(W467), .ZN(O255));
  NOR2X1 G592 (.A1(W671), .A2(W1074), .ZN(W2129));
  NOR2X1 G593 (.A1(W520), .A2(W1282), .ZN(O253));
  NOR2X1 G594 (.A1(W1113), .A2(W535), .ZN(W1934));
  NOR2X1 G595 (.A1(W987), .A2(I142), .ZN(W1931));
  NOR2X1 G596 (.A1(W1474), .A2(W1162), .ZN(O315));
  NOR2X1 G597 (.A1(I4), .A2(W1523), .ZN(W2134));
  NOR2X1 G598 (.A1(W1526), .A2(W280), .ZN(O316));
  NOR2X1 G599 (.A1(W1166), .A2(W1428), .ZN(O317));
  NOR2X1 G600 (.A1(W51), .A2(W78), .ZN(O488));
  NOR2X1 G601 (.A1(W415), .A2(W1444), .ZN(W1541));
  NOR2X1 G602 (.A1(I117), .A2(W1153), .ZN(W2517));
  NOR2X1 G603 (.A1(W1498), .A2(W1330), .ZN(W1533));
  NOR2X1 G604 (.A1(I30), .A2(W1215), .ZN(W1531));
  NOR2X1 G605 (.A1(W2334), .A2(W906), .ZN(W2529));
  NOR2X1 G606 (.A1(W853), .A2(W829), .ZN(W1528));
  NOR2X1 G607 (.A1(W1022), .A2(W1694), .ZN(W2534));
  NOR2X1 G608 (.A1(W311), .A2(W297), .ZN(W1525));
  NOR2X1 G609 (.A1(W785), .A2(W470), .ZN(W1524));
  NOR2X1 G610 (.A1(W1036), .A2(W615), .ZN(W1523));
  NOR2X1 G611 (.A1(W1322), .A2(W1714), .ZN(O487));
  NOR2X1 G612 (.A1(W1098), .A2(W345), .ZN(W1519));
  NOR2X1 G613 (.A1(W526), .A2(W338), .ZN(O479));
  NOR2X1 G614 (.A1(W876), .A2(W347), .ZN(W1514));
  NOR2X1 G615 (.A1(W1363), .A2(W265), .ZN(W1513));
  NOR2X1 G616 (.A1(W2101), .A2(W955), .ZN(O494));
  NOR2X1 G617 (.A1(W2474), .A2(W244), .ZN(O496));
  NOR2X1 G618 (.A1(W982), .A2(W675), .ZN(W2555));
  NOR2X1 G619 (.A1(W1270), .A2(W325), .ZN(W1507));
  NOR2X1 G620 (.A1(W489), .A2(W1283), .ZN(W1506));
  NOR2X1 G621 (.A1(W579), .A2(W1194), .ZN(W1504));
  NOR2X1 G622 (.A1(W787), .A2(I166), .ZN(W2559));
  NOR2X1 G623 (.A1(W1592), .A2(W91), .ZN(W2560));
  NOR2X1 G624 (.A1(W1038), .A2(W1218), .ZN(W1501));
  NOR2X1 G625 (.A1(W1457), .A2(W1282), .ZN(W2496));
  NOR2X1 G626 (.A1(W550), .A2(W524), .ZN(W1576));
  NOR2X1 G627 (.A1(W1196), .A2(W700), .ZN(O147));
  NOR2X1 G628 (.A1(W1055), .A2(W1839), .ZN(O467));
  NOR2X1 G629 (.A1(W1268), .A2(W1020), .ZN(O146));
  NOR2X1 G630 (.A1(W2257), .A2(W69), .ZN(O468));
  NOR2X1 G631 (.A1(W376), .A2(W32), .ZN(W2491));
  NOR2X1 G632 (.A1(W410), .A2(W923), .ZN(W1568));
  NOR2X1 G633 (.A1(W2408), .A2(W244), .ZN(O469));
  NOR2X1 G634 (.A1(W167), .A2(W448), .ZN(O144));
  NOR2X1 G635 (.A1(W4), .A2(W326), .ZN(W2494));
  NOR2X1 G636 (.A1(I60), .A2(W627), .ZN(W2495));
  NOR2X1 G637 (.A1(W642), .A2(W1069), .ZN(W1562));
  NOR2X1 G638 (.A1(W617), .A2(W826), .ZN(W1500));
  NOR2X1 G639 (.A1(W450), .A2(I102), .ZN(W1560));
  NOR2X1 G640 (.A1(W912), .A2(W1203), .ZN(W1559));
  NOR2X1 G641 (.A1(W442), .A2(W1161), .ZN(O142));
  NOR2X1 G642 (.A1(W1479), .A2(W1988), .ZN(W2497));
  NOR2X1 G643 (.A1(I175), .A2(W1137), .ZN(O140));
  NOR2X1 G644 (.A1(I174), .A2(W1341), .ZN(W2500));
  NOR2X1 G645 (.A1(W309), .A2(W1480), .ZN(O473));
  NOR2X1 G646 (.A1(W855), .A2(W1226), .ZN(W1551));
  NOR2X1 G647 (.A1(W2472), .A2(W1644), .ZN(O474));
  NOR2X1 G648 (.A1(W2318), .A2(W1073), .ZN(W2507));
  NOR2X1 G649 (.A1(W1655), .A2(W856), .ZN(W2510));
  NOR2X1 G650 (.A1(W1056), .A2(W1388), .ZN(W1437));
  NOR2X1 G651 (.A1(W811), .A2(W977), .ZN(O531));
  NOR2X1 G652 (.A1(W877), .A2(W97), .ZN(O533));
  NOR2X1 G653 (.A1(W2612), .A2(W1335), .ZN(W2623));
  NOR2X1 G654 (.A1(W1161), .A2(W650), .ZN(W1448));
  NOR2X1 G655 (.A1(W571), .A2(W64), .ZN(W1447));
  NOR2X1 G656 (.A1(W291), .A2(W537), .ZN(W1445));
  NOR2X1 G657 (.A1(W1116), .A2(W538), .ZN(W1444));
  NOR2X1 G658 (.A1(W1495), .A2(W1499), .ZN(O536));
  NOR2X1 G659 (.A1(I78), .A2(W140), .ZN(W1442));
  NOR2X1 G660 (.A1(I10), .A2(W985), .ZN(W1440));
  NOR2X1 G661 (.A1(W1137), .A2(W434), .ZN(W1439));
  NOR2X1 G662 (.A1(W1406), .A2(W1219), .ZN(O124));
  NOR2X1 G663 (.A1(W331), .A2(W490), .ZN(O125));
  NOR2X1 G664 (.A1(W1916), .A2(I75), .ZN(W2633));
  NOR2X1 G665 (.A1(W1029), .A2(I27), .ZN(W1435));
  NOR2X1 G666 (.A1(W178), .A2(W589), .ZN(W1433));
  NOR2X1 G667 (.A1(W97), .A2(W288), .ZN(O120));
  NOR2X1 G668 (.A1(W629), .A2(W1010), .ZN(W1430));
  NOR2X1 G669 (.A1(W186), .A2(W260), .ZN(W1428));
  NOR2X1 G670 (.A1(W1185), .A2(W264), .ZN(W2639));
  NOR2X1 G671 (.A1(W787), .A2(W596), .ZN(W1426));
  NOR2X1 G672 (.A1(W742), .A2(W2495), .ZN(O542));
  NOR2X1 G673 (.A1(W432), .A2(W1263), .ZN(W2642));
  NOR2X1 G674 (.A1(W2482), .A2(W2575), .ZN(O544));
  NOR2X1 G675 (.A1(W900), .A2(W315), .ZN(W1482));
  NOR2X1 G676 (.A1(W211), .A2(W424), .ZN(W2561));
  NOR2X1 G677 (.A1(W963), .A2(W438), .ZN(W1498));
  NOR2X1 G678 (.A1(W236), .A2(W1937), .ZN(O502));
  NOR2X1 G679 (.A1(W1119), .A2(W1385), .ZN(W1495));
  NOR2X1 G680 (.A1(W585), .A2(W66), .ZN(W1491));
  NOR2X1 G681 (.A1(W93), .A2(W6), .ZN(W1490));
  NOR2X1 G682 (.A1(W914), .A2(W401), .ZN(W1488));
  NOR2X1 G683 (.A1(W541), .A2(W1474), .ZN(W1487));
  NOR2X1 G684 (.A1(W60), .A2(W2251), .ZN(O509));
  NOR2X1 G685 (.A1(W23), .A2(W148), .ZN(O128));
  NOR2X1 G686 (.A1(W1993), .A2(W1792), .ZN(W2577));
  NOR2X1 G687 (.A1(I75), .A2(W869), .ZN(W1483));
  NOR2X1 G688 (.A1(W1133), .A2(W894), .ZN(W1577));
  NOR2X1 G689 (.A1(W1899), .A2(W159), .ZN(W2583));
  NOR2X1 G690 (.A1(W166), .A2(W828), .ZN(W1479));
  NOR2X1 G691 (.A1(W748), .A2(I52), .ZN(O512));
  NOR2X1 G692 (.A1(W2472), .A2(W2104), .ZN(O514));
  NOR2X1 G693 (.A1(W1271), .A2(I126), .ZN(W1474));
  NOR2X1 G694 (.A1(W776), .A2(W2537), .ZN(O516));
  NOR2X1 G695 (.A1(W1223), .A2(W1046), .ZN(W2598));
  NOR2X1 G696 (.A1(W802), .A2(W2055), .ZN(W2601));
  NOR2X1 G697 (.A1(I112), .A2(W1149), .ZN(W1464));
  NOR2X1 G698 (.A1(W2081), .A2(W1958), .ZN(W2611));
  NOR2X1 G699 (.A1(W1369), .A2(W386), .ZN(W2612));
  NOR2X1 G700 (.A1(W359), .A2(W1288), .ZN(O424));
  NOR2X1 G701 (.A1(W712), .A2(W644), .ZN(O405));
  NOR2X1 G702 (.A1(W1638), .A2(W1250), .ZN(O408));
  NOR2X1 G703 (.A1(I88), .A2(W871), .ZN(W1691));
  NOR2X1 G704 (.A1(W444), .A2(W1118), .ZN(O413));
  NOR2X1 G705 (.A1(W450), .A2(W1028), .ZN(W1684));
  NOR2X1 G706 (.A1(W2295), .A2(W1161), .ZN(W2378));
  NOR2X1 G707 (.A1(W2023), .A2(W119), .ZN(W2384));
  NOR2X1 G708 (.A1(W456), .A2(W856), .ZN(W1677));
  NOR2X1 G709 (.A1(W393), .A2(W1278), .ZN(W1676));
  NOR2X1 G710 (.A1(W448), .A2(W1465), .ZN(O421));
  NOR2X1 G711 (.A1(W483), .A2(W1475), .ZN(W1671));
  NOR2X1 G712 (.A1(W2104), .A2(W818), .ZN(W2392));
  NOR2X1 G713 (.A1(W277), .A2(W1374), .ZN(W1698));
  NOR2X1 G714 (.A1(W1299), .A2(W795), .ZN(W1668));
  NOR2X1 G715 (.A1(W518), .A2(W871), .ZN(W1664));
  NOR2X1 G716 (.A1(W119), .A2(I135), .ZN(O426));
  NOR2X1 G717 (.A1(W1470), .A2(W850), .ZN(O175));
  NOR2X1 G718 (.A1(W2036), .A2(W431), .ZN(W2398));
  NOR2X1 G719 (.A1(W34), .A2(W212), .ZN(O427));
  NOR2X1 G720 (.A1(W96), .A2(W761), .ZN(W1659));
  NOR2X1 G721 (.A1(W1116), .A2(W340), .ZN(W1658));
  NOR2X1 G722 (.A1(W2015), .A2(W665), .ZN(W2400));
  NOR2X1 G723 (.A1(W373), .A2(W2240), .ZN(W2402));
  NOR2X1 G724 (.A1(W944), .A2(W733), .ZN(W1655));
  NOR2X1 G725 (.A1(W355), .A2(W1170), .ZN(O190));
  NOR2X1 G726 (.A1(W2146), .A2(W1361), .ZN(O397));
  NOR2X1 G727 (.A1(W175), .A2(W1513), .ZN(W1727));
  NOR2X1 G728 (.A1(W925), .A2(W881), .ZN(W2333));
  NOR2X1 G729 (.A1(W754), .A2(I36), .ZN(W2336));
  NOR2X1 G730 (.A1(W1578), .A2(W1166), .ZN(W1722));
  NOR2X1 G731 (.A1(W2065), .A2(W1559), .ZN(W2337));
  NOR2X1 G732 (.A1(W2195), .A2(W1587), .ZN(O399));
  NOR2X1 G733 (.A1(W1795), .A2(W1314), .ZN(W2339));
  NOR2X1 G734 (.A1(W649), .A2(W1126), .ZN(W1718));
  NOR2X1 G735 (.A1(W384), .A2(W1168), .ZN(O191));
  NOR2X1 G736 (.A1(W1329), .A2(W427), .ZN(W2340));
  NOR2X1 G737 (.A1(I4), .A2(W318), .ZN(W1714));
  NOR2X1 G738 (.A1(W291), .A2(W932), .ZN(W1653));
  NOR2X1 G739 (.A1(W2323), .A2(W185), .ZN(W2344));
  NOR2X1 G740 (.A1(W2149), .A2(W1953), .ZN(W2345));
  NOR2X1 G741 (.A1(W1331), .A2(W831), .ZN(O402));
  NOR2X1 G742 (.A1(W1589), .A2(W625), .ZN(O188));
  NOR2X1 G743 (.A1(W936), .A2(W1454), .ZN(W2348));
  NOR2X1 G744 (.A1(W415), .A2(W245), .ZN(W1706));
  NOR2X1 G745 (.A1(W607), .A2(W423), .ZN(O187));
  NOR2X1 G746 (.A1(I180), .A2(W1042), .ZN(O186));
  NOR2X1 G747 (.A1(W199), .A2(W1127), .ZN(W1702));
  NOR2X1 G748 (.A1(I146), .A2(W724), .ZN(W1701));
  NOR2X1 G749 (.A1(W737), .A2(W1196), .ZN(O184));
  NOR2X1 G750 (.A1(W2280), .A2(W572), .ZN(W2465));
  NOR2X1 G751 (.A1(W42), .A2(W189), .ZN(W1616));
  NOR2X1 G752 (.A1(W401), .A2(W924), .ZN(W1614));
  NOR2X1 G753 (.A1(W100), .A2(I24), .ZN(W2440));
  NOR2X1 G754 (.A1(W114), .A2(W113), .ZN(O154));
  NOR2X1 G755 (.A1(W514), .A2(I40), .ZN(O448));
  NOR2X1 G756 (.A1(W953), .A2(W1282), .ZN(O449));
  NOR2X1 G757 (.A1(W1952), .A2(W2262), .ZN(W2449));
  NOR2X1 G758 (.A1(W1600), .A2(W1200), .ZN(W2450));
  NOR2X1 G759 (.A1(W1946), .A2(W231), .ZN(W2451));
  NOR2X1 G760 (.A1(W668), .A2(W1255), .ZN(W1600));
  NOR2X1 G761 (.A1(W2446), .A2(W358), .ZN(W2460));
  NOR2X1 G762 (.A1(W2384), .A2(W2352), .ZN(W2462));
  NOR2X1 G763 (.A1(W966), .A2(W840), .ZN(O156));
  NOR2X1 G764 (.A1(W2217), .A2(W18), .ZN(W2466));
  NOR2X1 G765 (.A1(W1168), .A2(W1474), .ZN(O458));
  NOR2X1 G766 (.A1(W765), .A2(W273), .ZN(O150));
  NOR2X1 G767 (.A1(W351), .A2(W2006), .ZN(O460));
  NOR2X1 G768 (.A1(W1692), .A2(W1208), .ZN(O462));
  NOR2X1 G769 (.A1(W946), .A2(W853), .ZN(W1584));
  NOR2X1 G770 (.A1(W287), .A2(W1363), .ZN(W2482));
  NOR2X1 G771 (.A1(W1666), .A2(W2420), .ZN(O465));
  NOR2X1 G772 (.A1(W229), .A2(W84), .ZN(O148));
  NOR2X1 G773 (.A1(W115), .A2(W660), .ZN(O466));
  NOR2X1 G774 (.A1(W426), .A2(W700), .ZN(W1578));
  NOR2X1 G775 (.A1(W1137), .A2(W303), .ZN(O434));
  NOR2X1 G776 (.A1(W305), .A2(W1599), .ZN(W1650));
  NOR2X1 G777 (.A1(W1160), .A2(W2384), .ZN(W2408));
  NOR2X1 G778 (.A1(W417), .A2(W437), .ZN(W1645));
  NOR2X1 G779 (.A1(W528), .A2(W563), .ZN(W1644));
  NOR2X1 G780 (.A1(W120), .A2(W328), .ZN(O167));
  NOR2X1 G781 (.A1(W57), .A2(W2230), .ZN(W2412));
  NOR2X1 G782 (.A1(W1508), .A2(W881), .ZN(O165));
  NOR2X1 G783 (.A1(W749), .A2(W1255), .ZN(O164));
  NOR2X1 G784 (.A1(W1251), .A2(W1057), .ZN(O163));
  NOR2X1 G785 (.A1(W1074), .A2(W426), .ZN(O432));
  NOR2X1 G786 (.A1(W430), .A2(W2305), .ZN(O433));
  NOR2X1 G787 (.A1(W1277), .A2(W1581), .ZN(O779));
  NOR2X1 G788 (.A1(W2224), .A2(W1722), .ZN(O435));
  NOR2X1 G789 (.A1(W54), .A2(W58), .ZN(O436));
  NOR2X1 G790 (.A1(W1920), .A2(W1429), .ZN(W2421));
  NOR2X1 G791 (.A1(W864), .A2(W1451), .ZN(W1630));
  NOR2X1 G792 (.A1(W1105), .A2(W2107), .ZN(O440));
  NOR2X1 G793 (.A1(W1381), .A2(W1925), .ZN(W2424));
  NOR2X1 G794 (.A1(W1072), .A2(W994), .ZN(O159));
  NOR2X1 G795 (.A1(W1560), .A2(W563), .ZN(W2426));
  NOR2X1 G796 (.A1(I126), .A2(W289), .ZN(W1623));
  NOR2X1 G797 (.A1(W971), .A2(I137), .ZN(W1620));
  NOR2X1 G798 (.A1(W973), .A2(W611), .ZN(W2436));
  NOR2X1 G799 (.A1(W1512), .A2(W2830), .ZN(O1192));
  NOR2X1 G800 (.A1(I29), .A2(I52), .ZN(W184));
  NOR2X1 G801 (.A1(W375), .A2(I112), .ZN(W486));
  NOR2X1 G802 (.A1(W58), .A2(I185), .ZN(W185));
  NOR2X1 G803 (.A1(W3631), .A2(W1716), .ZN(O1447));
  NOR2X1 G804 (.A1(I98), .A2(I92), .ZN(W187));
  NOR2X1 G805 (.A1(I86), .A2(I21), .ZN(W483));
  NOR2X1 G806 (.A1(W33), .A2(I57), .ZN(W482));
  NOR2X1 G807 (.A1(W382), .A2(W344), .ZN(W481));
  NOR2X1 G808 (.A1(I55), .A2(I68), .ZN(W188));
  NOR2X1 G809 (.A1(W2931), .A2(I14), .ZN(O1191));
  NOR2X1 G810 (.A1(W1268), .A2(W152), .ZN(O1183));
  NOR2X1 G811 (.A1(W31), .A2(W77), .ZN(W189));
  NOR2X1 G812 (.A1(W1842), .A2(W3019), .ZN(O1446));
  NOR2X1 G813 (.A1(W177), .A2(W2340), .ZN(O1444));
  NOR2X1 G814 (.A1(I13), .A2(W594), .ZN(O1195));
  NOR2X1 G815 (.A1(W96), .A2(W142), .ZN(W194));
  NOR2X1 G816 (.A1(W3735), .A2(W2518), .ZN(O1440));
  NOR2X1 G817 (.A1(W29), .A2(W162), .ZN(W196));
  NOR2X1 G818 (.A1(W176), .A2(W75), .ZN(W197));
  NOR2X1 G819 (.A1(W2496), .A2(W3389), .ZN(W3634));
  NOR2X1 G820 (.A1(I194), .A2(I5), .ZN(W176));
  NOR2X1 G821 (.A1(W353), .A2(W323), .ZN(W505));
  NOR2X1 G822 (.A1(W115), .A2(W56), .ZN(W504));
  NOR2X1 G823 (.A1(W449), .A2(W427), .ZN(W503));
  NOR2X1 G824 (.A1(W1004), .A2(W543), .ZN(O1170));
  NOR2X1 G825 (.A1(I142), .A2(W72), .ZN(W173));
  NOR2X1 G826 (.A1(W329), .A2(W271), .ZN(W501));
  NOR2X1 G827 (.A1(W9), .A2(W352), .ZN(O1171));
  NOR2X1 G828 (.A1(I109), .A2(I26), .ZN(W174));
  NOR2X1 G829 (.A1(W498), .A2(W2654), .ZN(O1172));
  NOR2X1 G830 (.A1(W2465), .A2(W3562), .ZN(O1199));
  NOR2X1 G831 (.A1(W107), .A2(W112), .ZN(W178));
  NOR2X1 G832 (.A1(W3080), .A2(W2674), .ZN(W3603));
  NOR2X1 G833 (.A1(I54), .A2(W122), .ZN(W179));
  NOR2X1 G834 (.A1(W3193), .A2(W1535), .ZN(O1178));
  NOR2X1 G835 (.A1(W2489), .A2(W248), .ZN(O1180));
  NOR2X1 G836 (.A1(I79), .A2(I95), .ZN(W180));
  NOR2X1 G837 (.A1(W178), .A2(I109), .ZN(W490));
  NOR2X1 G838 (.A1(I123), .A2(W96), .ZN(W182));
  NOR2X1 G839 (.A1(I140), .A2(W4), .ZN(W183));
  NOR2X1 G840 (.A1(W577), .A2(W3458), .ZN(W3663));
  NOR2X1 G841 (.A1(W138), .A2(I188), .ZN(W205));
  NOR2X1 G842 (.A1(W1967), .A2(W2144), .ZN(O1221));
  NOR2X1 G843 (.A1(W159), .A2(I56), .ZN(W206));
  NOR2X1 G844 (.A1(W3020), .A2(W252), .ZN(W3893));
  NOR2X1 G845 (.A1(W59), .A2(W2), .ZN(W209));
  NOR2X1 G846 (.A1(W40), .A2(W174), .ZN(W453));
  NOR2X1 G847 (.A1(W66), .A2(W9), .ZN(W210));
  NOR2X1 G848 (.A1(W155), .A2(I158), .ZN(W451));
  NOR2X1 G849 (.A1(W3114), .A2(W2028), .ZN(O1223));
  NOR2X1 G850 (.A1(W2656), .A2(W1253), .ZN(O1220));
  NOR2X1 G851 (.A1(I64), .A2(W130), .ZN(W212));
  NOR2X1 G852 (.A1(W375), .A2(W305), .ZN(W448));
  NOR2X1 G853 (.A1(W167), .A2(W31), .ZN(W213));
  NOR2X1 G854 (.A1(W1203), .A2(W1884), .ZN(O1225));
  NOR2X1 G855 (.A1(W834), .A2(W1467), .ZN(W3666));
  NOR2X1 G856 (.A1(W3397), .A2(W2155), .ZN(O1428));
  NOR2X1 G857 (.A1(W695), .A2(W315), .ZN(O1226));
  NOR2X1 G858 (.A1(W1338), .A2(W3320), .ZN(O1229));
  NOR2X1 G859 (.A1(W3245), .A2(W1792), .ZN(O1230));
  NOR2X1 G860 (.A1(I121), .A2(W80), .ZN(W201));
  NOR2X1 G861 (.A1(W178), .A2(I140), .ZN(W472));
  NOR2X1 G862 (.A1(W2728), .A2(W1680), .ZN(O1201));
  NOR2X1 G863 (.A1(I132), .A2(W109), .ZN(W198));
  NOR2X1 G864 (.A1(W2278), .A2(W571), .ZN(O1205));
  NOR2X1 G865 (.A1(W402), .A2(W459), .ZN(W468));
  NOR2X1 G866 (.A1(W7), .A2(W331), .ZN(W467));
  NOR2X1 G867 (.A1(W353), .A2(I24), .ZN(W466));
  NOR2X1 G868 (.A1(W3668), .A2(W3436), .ZN(O1438));
  NOR2X1 G869 (.A1(W290), .A2(W438), .ZN(W465));
  NOR2X1 G870 (.A1(W2278), .A2(W1274), .ZN(O1169));
  NOR2X1 G871 (.A1(I24), .A2(I169), .ZN(W202));
  NOR2X1 G872 (.A1(W13), .A2(W196), .ZN(W463));
  NOR2X1 G873 (.A1(W1578), .A2(W3494), .ZN(O1207));
  NOR2X1 G874 (.A1(W736), .A2(W2392), .ZN(O1211));
  NOR2X1 G875 (.A1(W1738), .A2(W1215), .ZN(W3650));
  NOR2X1 G876 (.A1(W996), .A2(W1903), .ZN(O1214));
  NOR2X1 G877 (.A1(W3013), .A2(W2366), .ZN(O1215));
  NOR2X1 G878 (.A1(W3169), .A2(W1219), .ZN(O1435));
  NOR2X1 G879 (.A1(W449), .A2(W29), .ZN(W456));
  NOR2X1 G880 (.A1(W1325), .A2(W2885), .ZN(O1486));
  NOR2X1 G881 (.A1(I160), .A2(I50), .ZN(W142));
  NOR2X1 G882 (.A1(W3452), .A2(W3043), .ZN(W3537));
  NOR2X1 G883 (.A1(W992), .A2(W2774), .ZN(W3538));
  NOR2X1 G884 (.A1(W42), .A2(W77), .ZN(W144));
  NOR2X1 G885 (.A1(W41), .A2(I169), .ZN(O1489));
  NOR2X1 G886 (.A1(W2316), .A2(W861), .ZN(O1128));
  NOR2X1 G887 (.A1(W3356), .A2(I184), .ZN(O1129));
  NOR2X1 G888 (.A1(I13), .A2(W129), .ZN(W147));
  NOR2X1 G889 (.A1(I48), .A2(I136), .ZN(O1130));
  NOR2X1 G890 (.A1(W289), .A2(I64), .ZN(W568));
  NOR2X1 G891 (.A1(W2761), .A2(W1746), .ZN(O1485));
  NOR2X1 G892 (.A1(W1060), .A2(W297), .ZN(O1133));
  NOR2X1 G893 (.A1(I34), .A2(W344), .ZN(O1134));
  NOR2X1 G894 (.A1(W169), .A2(I112), .ZN(W554));
  NOR2X1 G895 (.A1(I163), .A2(W2508), .ZN(O1483));
  NOR2X1 G896 (.A1(W1897), .A2(W1551), .ZN(O1481));
  NOR2X1 G897 (.A1(W1978), .A2(W922), .ZN(O1137));
  NOR2X1 G898 (.A1(I117), .A2(I182), .ZN(W153));
  NOR2X1 G899 (.A1(W314), .A2(W0), .ZN(O1138));
  NOR2X1 G900 (.A1(W191), .A2(W285), .ZN(W578));
  NOR2X1 G901 (.A1(I71), .A2(W63), .ZN(W127));
  NOR2X1 G902 (.A1(W507), .A2(W56), .ZN(W586));
  NOR2X1 G903 (.A1(W1099), .A2(W2533), .ZN(O1102));
  NOR2X1 G904 (.A1(W738), .A2(W2559), .ZN(O1104));
  NOR2X1 G905 (.A1(I80), .A2(W217), .ZN(O14));
  NOR2X1 G906 (.A1(W2446), .A2(W1142), .ZN(O1107));
  NOR2X1 G907 (.A1(W3421), .A2(W3568), .ZN(O1505));
  NOR2X1 G908 (.A1(W3353), .A2(W752), .ZN(O1111));
  NOR2X1 G909 (.A1(W401), .A2(W477), .ZN(W579));
  NOR2X1 G910 (.A1(W2531), .A2(W2997), .ZN(O1143));
  NOR2X1 G911 (.A1(I191), .A2(W73), .ZN(W133));
  NOR2X1 G912 (.A1(W3066), .A2(W445), .ZN(O1113));
  NOR2X1 G913 (.A1(W55), .A2(W114), .ZN(W134));
  NOR2X1 G914 (.A1(I94), .A2(W2), .ZN(W135));
  NOR2X1 G915 (.A1(W1712), .A2(W2855), .ZN(O1498));
  NOR2X1 G916 (.A1(W129), .A2(I132), .ZN(W138));
  NOR2X1 G917 (.A1(W508), .A2(W88), .ZN(W571));
  NOR2X1 G918 (.A1(W442), .A2(W9), .ZN(O13));
  NOR2X1 G919 (.A1(W50), .A2(W23), .ZN(W140));
  NOR2X1 G920 (.A1(W2656), .A2(W490), .ZN(W3583));
  NOR2X1 G921 (.A1(W2375), .A2(W1428), .ZN(O1152));
  NOR2X1 G922 (.A1(W3392), .A2(W1114), .ZN(O1156));
  NOR2X1 G923 (.A1(W3417), .A2(W1697), .ZN(O1158));
  NOR2X1 G924 (.A1(W2974), .A2(W3054), .ZN(O1159));
  NOR2X1 G925 (.A1(I62), .A2(I184), .ZN(W523));
  NOR2X1 G926 (.A1(W1494), .A2(W2666), .ZN(O1455));
  NOR2X1 G927 (.A1(I6), .A2(W300), .ZN(W521));
  NOR2X1 G928 (.A1(W204), .A2(W444), .ZN(W520));
  NOR2X1 G929 (.A1(I190), .A2(W80), .ZN(W517));
  NOR2X1 G930 (.A1(W512), .A2(W4), .ZN(W530));
  NOR2X1 G931 (.A1(I66), .A2(W32), .ZN(W171));
  NOR2X1 G932 (.A1(W173), .A2(W353), .ZN(W514));
  NOR2X1 G933 (.A1(W232), .A2(W148), .ZN(O1162));
  NOR2X1 G934 (.A1(W195), .A2(W321), .ZN(W511));
  NOR2X1 G935 (.A1(I7), .A2(W406), .ZN(W510));
  NOR2X1 G936 (.A1(W2713), .A2(W29), .ZN(O1165));
  NOR2X1 G937 (.A1(W696), .A2(W2517), .ZN(O1166));
  NOR2X1 G938 (.A1(I121), .A2(I58), .ZN(W172));
  NOR2X1 G939 (.A1(W277), .A2(W391), .ZN(W507));
  NOR2X1 G940 (.A1(I96), .A2(I186), .ZN(W541));
  NOR2X1 G941 (.A1(W41), .A2(I0), .ZN(W154));
  NOR2X1 G942 (.A1(W61), .A2(I145), .ZN(W156));
  NOR2X1 G943 (.A1(W285), .A2(I92), .ZN(W544));
  NOR2X1 G944 (.A1(W1070), .A2(W3089), .ZN(O1473));
  NOR2X1 G945 (.A1(W141), .A2(W116), .ZN(W158));
  NOR2X1 G946 (.A1(W37), .A2(I169), .ZN(W159));
  NOR2X1 G947 (.A1(W1331), .A2(W390), .ZN(O1145));
  NOR2X1 G948 (.A1(I134), .A2(W114), .ZN(W160));
  NOR2X1 G949 (.A1(W2442), .A2(W1116), .ZN(O1146));
  NOR2X1 G950 (.A1(W158), .A2(I103), .ZN(W218));
  NOR2X1 G951 (.A1(W658), .A2(W351), .ZN(O1147));
  NOR2X1 G952 (.A1(I71), .A2(W187), .ZN(W539));
  NOR2X1 G953 (.A1(W359), .A2(I84), .ZN(W537));
  NOR2X1 G954 (.A1(W1305), .A2(W3198), .ZN(O1150));
  NOR2X1 G955 (.A1(W43), .A2(W493), .ZN(W534));
  NOR2X1 G956 (.A1(W3609), .A2(W1745), .ZN(O1466));
  NOR2X1 G957 (.A1(W2889), .A2(W3292), .ZN(O1464));
  NOR2X1 G958 (.A1(W11), .A2(W417), .ZN(W532));
  NOR2X1 G959 (.A1(W267), .A2(W160), .ZN(W531));
  NOR2X1 G960 (.A1(W3243), .A2(W1003), .ZN(O1380));
  NOR2X1 G961 (.A1(W68), .A2(W32), .ZN(W260));
  NOR2X1 G962 (.A1(W159), .A2(W2), .ZN(W346));
  NOR2X1 G963 (.A1(W1115), .A2(W1821), .ZN(O1394));
  NOR2X1 G964 (.A1(W2993), .A2(W1605), .ZN(O1316));
  NOR2X1 G965 (.A1(W2175), .A2(W1703), .ZN(O1318));
  NOR2X1 G966 (.A1(W2709), .A2(W1694), .ZN(O1319));
  NOR2X1 G967 (.A1(W96), .A2(W190), .ZN(W339));
  NOR2X1 G968 (.A1(W1531), .A2(W2009), .ZN(O1320));
  NOR2X1 G969 (.A1(W232), .A2(W212), .ZN(W268));
  NOR2X1 G970 (.A1(W3302), .A2(W1762), .ZN(O1322));
  NOR2X1 G971 (.A1(W2913), .A2(W2551), .ZN(O1307));
  NOR2X1 G972 (.A1(W1444), .A2(W3042), .ZN(O1326));
  NOR2X1 G973 (.A1(W3443), .A2(W18), .ZN(O1327));
  NOR2X1 G974 (.A1(W263), .A2(W149), .ZN(W271));
  NOR2X1 G975 (.A1(I81), .A2(I75), .ZN(W329));
  NOR2X1 G976 (.A1(W180), .A2(W269), .ZN(W272));
  NOR2X1 G977 (.A1(W363), .A2(W3654), .ZN(O1379));
  NOR2X1 G978 (.A1(W275), .A2(W1767), .ZN(O1332));
  NOR2X1 G979 (.A1(W147), .A2(I162), .ZN(W274));
  NOR2X1 G980 (.A1(I78), .A2(W225), .ZN(W275));
  NOR2X1 G981 (.A1(W147), .A2(I120), .ZN(W356));
  NOR2X1 G982 (.A1(W2909), .A2(W3107), .ZN(O1291));
  NOR2X1 G983 (.A1(W276), .A2(I68), .ZN(W366));
  NOR2X1 G984 (.A1(W599), .A2(W1786), .ZN(O1402));
  NOR2X1 G985 (.A1(W211), .A2(W357), .ZN(W365));
  NOR2X1 G986 (.A1(I130), .A2(W2705), .ZN(W3741));
  NOR2X1 G987 (.A1(W78), .A2(W321), .ZN(O1401));
  NOR2X1 G988 (.A1(W155), .A2(W3058), .ZN(O1295));
  NOR2X1 G989 (.A1(W2804), .A2(W3509), .ZN(O1296));
  NOR2X1 G990 (.A1(W729), .A2(W2767), .ZN(O1399));
  NOR2X1 G991 (.A1(W3184), .A2(W3500), .ZN(O1377));
  NOR2X1 G992 (.A1(W308), .A2(W298), .ZN(W355));
  NOR2X1 G993 (.A1(W1476), .A2(W1636), .ZN(O1301));
  NOR2X1 G994 (.A1(W68), .A2(W90), .ZN(O5));
  NOR2X1 G995 (.A1(I102), .A2(I76), .ZN(W254));
  NOR2X1 G996 (.A1(W112), .A2(W69), .ZN(W256));
  NOR2X1 G997 (.A1(I175), .A2(W98), .ZN(W257));
  NOR2X1 G998 (.A1(I112), .A2(W140), .ZN(W258));
  NOR2X1 G999 (.A1(W256), .A2(W1041), .ZN(O1305));
  NOR2X1 G1000 (.A1(I118), .A2(W115), .ZN(W350));
  NOR2X1 G1001 (.A1(W2721), .A2(W107), .ZN(O1358));
  NOR2X1 G1002 (.A1(W1217), .A2(W3451), .ZN(O1353));
  NOR2X1 G1003 (.A1(I157), .A2(I23), .ZN(W307));
  NOR2X1 G1004 (.A1(I162), .A2(I160), .ZN(W306));
  NOR2X1 G1005 (.A1(I144), .A2(I65), .ZN(W304));
  NOR2X1 G1006 (.A1(W219), .A2(W259), .ZN(W303));
  NOR2X1 G1007 (.A1(W84), .A2(I9), .ZN(W302));
  NOR2X1 G1008 (.A1(W2468), .A2(W328), .ZN(O1356));
  NOR2X1 G1009 (.A1(W1412), .A2(W1062), .ZN(O1370));
  NOR2X1 G1010 (.A1(W188), .A2(I193), .ZN(W300));
  NOR2X1 G1011 (.A1(W3650), .A2(W3117), .ZN(O1351));
  NOR2X1 G1012 (.A1(W30), .A2(W8), .ZN(W298));
  NOR2X1 G1013 (.A1(W1949), .A2(W1773), .ZN(O1359));
  NOR2X1 G1014 (.A1(W1546), .A2(W1551), .ZN(O1361));
  NOR2X1 G1015 (.A1(W43), .A2(I115), .ZN(W295));
  NOR2X1 G1016 (.A1(W139), .A2(W51), .ZN(W294));
  NOR2X1 G1017 (.A1(W438), .A2(W3104), .ZN(O1362));
  NOR2X1 G1018 (.A1(W1590), .A2(I58), .ZN(O1364));
  NOR2X1 G1019 (.A1(W1742), .A2(W1507), .ZN(O1368));
  NOR2X1 G1020 (.A1(W991), .A2(W2339), .ZN(O1367));
  NOR2X1 G1021 (.A1(I21), .A2(W686), .ZN(O1341));
  NOR2X1 G1022 (.A1(W2010), .A2(W1738), .ZN(O1333));
  NOR2X1 G1023 (.A1(W221), .A2(W1349), .ZN(O1376));
  NOR2X1 G1024 (.A1(W116), .A2(W87), .ZN(W324));
  NOR2X1 G1025 (.A1(W114), .A2(I168), .ZN(W323));
  NOR2X1 G1026 (.A1(I178), .A2(W84), .ZN(W279));
  NOR2X1 G1027 (.A1(I30), .A2(W86), .ZN(W280));
  NOR2X1 G1028 (.A1(W1117), .A2(W3291), .ZN(O1339));
  NOR2X1 G1029 (.A1(W1411), .A2(W958), .ZN(O1340));
  NOR2X1 G1030 (.A1(W21), .A2(W232), .ZN(W281));
  NOR2X1 G1031 (.A1(W2653), .A2(W228), .ZN(O1289));
  NOR2X1 G1032 (.A1(W75), .A2(W981), .ZN(O1374));
  NOR2X1 G1033 (.A1(W85), .A2(W12), .ZN(W283));
  NOR2X1 G1034 (.A1(W3702), .A2(W1414), .ZN(W3799));
  NOR2X1 G1035 (.A1(W290), .A2(W301), .ZN(W315));
  NOR2X1 G1036 (.A1(W3621), .A2(I7), .ZN(O1373));
  NOR2X1 G1037 (.A1(W611), .A2(W2373), .ZN(W3802));
  NOR2X1 G1038 (.A1(W189), .A2(W2139), .ZN(O1347));
  NOR2X1 G1039 (.A1(W2842), .A2(I164), .ZN(O1350));
  NOR2X1 G1040 (.A1(I110), .A2(W82), .ZN(W310));
  NOR2X1 G1041 (.A1(W21), .A2(W124), .ZN(W230));
  NOR2X1 G1042 (.A1(W3050), .A2(W3603), .ZN(O1258));
  NOR2X1 G1043 (.A1(W341), .A2(W3088), .ZN(O1417));
  NOR2X1 G1044 (.A1(I27), .A2(W1037), .ZN(W3704));
  NOR2X1 G1045 (.A1(W2747), .A2(W2589), .ZN(W3705));
  NOR2X1 G1046 (.A1(W3324), .A2(W2034), .ZN(O1260));
  NOR2X1 G1047 (.A1(W1819), .A2(W1069), .ZN(O1261));
  NOR2X1 G1048 (.A1(W16), .A2(W256), .ZN(W411));
  NOR2X1 G1049 (.A1(W228), .A2(I121), .ZN(W410));
  NOR2X1 G1050 (.A1(W307), .A2(I112), .ZN(W409));
  NOR2X1 G1051 (.A1(W2542), .A2(W2316), .ZN(O1256));
  NOR2X1 G1052 (.A1(W193), .A2(I194), .ZN(W408));
  NOR2X1 G1053 (.A1(W380), .A2(W41), .ZN(W406));
  NOR2X1 G1054 (.A1(W267), .A2(W232), .ZN(W405));
  NOR2X1 G1055 (.A1(W3583), .A2(I128), .ZN(O1264));
  NOR2X1 G1056 (.A1(W197), .A2(W86), .ZN(W403));
  NOR2X1 G1057 (.A1(W827), .A2(W1090), .ZN(O942));
  NOR2X1 G1058 (.A1(W2075), .A2(W1645), .ZN(O1265));
  NOR2X1 G1059 (.A1(W290), .A2(W319), .ZN(W401));
  NOR2X1 G1060 (.A1(W186), .A2(I102), .ZN(W231));
  NOR2X1 G1061 (.A1(W101), .A2(W361), .ZN(W430));
  NOR2X1 G1062 (.A1(W631), .A2(W861), .ZN(O1236));
  NOR2X1 G1063 (.A1(W379), .A2(W173), .ZN(W436));
  NOR2X1 G1064 (.A1(I45), .A2(W142), .ZN(W219));
  NOR2X1 G1065 (.A1(W1543), .A2(W1458), .ZN(O1237));
  NOR2X1 G1066 (.A1(W97), .A2(I118), .ZN(W220));
  NOR2X1 G1067 (.A1(W3400), .A2(W699), .ZN(O1238));
  NOR2X1 G1068 (.A1(I132), .A2(W112), .ZN(W221));
  NOR2X1 G1069 (.A1(W3580), .A2(W1178), .ZN(O1240));
  NOR2X1 G1070 (.A1(W287), .A2(W189), .ZN(W431));
  NOR2X1 G1071 (.A1(W255), .A2(W197), .ZN(W400));
  NOR2X1 G1072 (.A1(W121), .A2(W343), .ZN(W428));
  NOR2X1 G1073 (.A1(W195), .A2(W390), .ZN(W425));
  NOR2X1 G1074 (.A1(W2401), .A2(W2598), .ZN(O1249));
  NOR2X1 G1075 (.A1(I79), .A2(W1563), .ZN(O1250));
  NOR2X1 G1076 (.A1(I10), .A2(W254), .ZN(W422));
  NOR2X1 G1077 (.A1(W254), .A2(W308), .ZN(W421));
  NOR2X1 G1078 (.A1(W3196), .A2(W1372), .ZN(O1253));
  NOR2X1 G1079 (.A1(W783), .A2(W562), .ZN(O1419));
  NOR2X1 G1080 (.A1(W3242), .A2(W2542), .ZN(O1418));
  NOR2X1 G1081 (.A1(W28), .A2(W146), .ZN(W241));
  NOR2X1 G1082 (.A1(W912), .A2(W2957), .ZN(O1277));
  NOR2X1 G1083 (.A1(W1100), .A2(W2507), .ZN(O1410));
  NOR2X1 G1084 (.A1(W162), .A2(W21), .ZN(W237));
  NOR2X1 G1085 (.A1(W41), .A2(W157), .ZN(W238));
  NOR2X1 G1086 (.A1(W90), .A2(I58), .ZN(W377));
  NOR2X1 G1087 (.A1(W340), .A2(I134), .ZN(W376));
  NOR2X1 G1088 (.A1(I123), .A2(I122), .ZN(W375));
  NOR2X1 G1089 (.A1(I190), .A2(I70), .ZN(W374));
  NOR2X1 G1090 (.A1(W266), .A2(W350), .ZN(W372));
  NOR2X1 G1091 (.A1(I196), .A2(W145), .ZN(W379));
  NOR2X1 G1092 (.A1(W3034), .A2(W1858), .ZN(O1406));
  NOR2X1 G1093 (.A1(W3708), .A2(W1892), .ZN(O1283));
  NOR2X1 G1094 (.A1(W24), .A2(W1727), .ZN(O1405));
  NOR2X1 G1095 (.A1(W230), .A2(W175), .ZN(W244));
  NOR2X1 G1096 (.A1(W1213), .A2(W2887), .ZN(W3735));
  NOR2X1 G1097 (.A1(W7), .A2(I40), .ZN(W245));
  NOR2X1 G1098 (.A1(I24), .A2(I28), .ZN(W246));
  NOR2X1 G1099 (.A1(W3750), .A2(W2367), .ZN(O1404));
  NOR2X1 G1100 (.A1(I112), .A2(W176), .ZN(W248));
  NOR2X1 G1101 (.A1(W308), .A2(W184), .ZN(W388));
  NOR2X1 G1102 (.A1(I13), .A2(W314), .ZN(W399));
  NOR2X1 G1103 (.A1(W22), .A2(W318), .ZN(W398));
  NOR2X1 G1104 (.A1(W180), .A2(W125), .ZN(W397));
  NOR2X1 G1105 (.A1(I78), .A2(I157), .ZN(W396));
  NOR2X1 G1106 (.A1(W1181), .A2(W1825), .ZN(O1266));
  NOR2X1 G1107 (.A1(W1674), .A2(W2473), .ZN(O1414));
  NOR2X1 G1108 (.A1(W109), .A2(I161), .ZN(W233));
  NOR2X1 G1109 (.A1(W306), .A2(W315), .ZN(W390));
  NOR2X1 G1110 (.A1(W3314), .A2(W3590), .ZN(O1273));
  NOR2X1 G1111 (.A1(I45), .A2(W2317), .ZN(W3560));
  NOR2X1 G1112 (.A1(W3047), .A2(W616), .ZN(O1274));
  NOR2X1 G1113 (.A1(I195), .A2(I108), .ZN(W386));
  NOR2X1 G1114 (.A1(W204), .A2(W192), .ZN(O8));
  NOR2X1 G1115 (.A1(W143), .A2(I195), .ZN(W384));
  NOR2X1 G1116 (.A1(W1742), .A2(W675), .ZN(O1411));
  NOR2X1 G1117 (.A1(W242), .A2(W201), .ZN(O7));
  NOR2X1 G1118 (.A1(W146), .A2(W36), .ZN(W382));
  NOR2X1 G1119 (.A1(W274), .A2(W1401), .ZN(O1276));
  NOR2X1 G1120 (.A1(W0), .A2(W230), .ZN(W380));
  NOR2X1 G1121 (.A1(I162), .A2(W218), .ZN(W700));
  NOR2X1 G1122 (.A1(I114), .A2(I115), .ZN(W57));
  NOR2X1 G1123 (.A1(W3781), .A2(W1050), .ZN(O1572));
  NOR2X1 G1124 (.A1(I120), .A2(I121), .ZN(W60));
  NOR2X1 G1125 (.A1(I122), .A2(I123), .ZN(W61));
  NOR2X1 G1126 (.A1(W2246), .A2(W346), .ZN(O1005));
  NOR2X1 G1127 (.A1(W2547), .A2(W1881), .ZN(O1570));
  NOR2X1 G1128 (.A1(W794), .A2(W567), .ZN(O1568));
  NOR2X1 G1129 (.A1(W396), .A2(W301), .ZN(W702));
  NOR2X1 G1130 (.A1(W286), .A2(W246), .ZN(O21));
  NOR2X1 G1131 (.A1(W674), .A2(W507), .ZN(W709));
  NOR2X1 G1132 (.A1(W449), .A2(W1030), .ZN(O1567));
  NOR2X1 G1133 (.A1(W547), .A2(W450), .ZN(W698));
  NOR2X1 G1134 (.A1(W75), .A2(W129), .ZN(W696));
  NOR2X1 G1135 (.A1(W290), .A2(W415), .ZN(W694));
  NOR2X1 G1136 (.A1(W287), .A2(I104), .ZN(W692));
  NOR2X1 G1137 (.A1(W2802), .A2(W552), .ZN(W3392));
  NOR2X1 G1138 (.A1(W1589), .A2(W2239), .ZN(O1012));
  NOR2X1 G1139 (.A1(W618), .A2(I174), .ZN(W688));
  NOR2X1 G1140 (.A1(I22), .A2(W117), .ZN(W687));
  NOR2X1 G1141 (.A1(W1464), .A2(W323), .ZN(O1578));
  NOR2X1 G1142 (.A1(W2232), .A2(W1539), .ZN(W3360));
  NOR2X1 G1143 (.A1(W396), .A2(I163), .ZN(W724));
  NOR2X1 G1144 (.A1(W2926), .A2(W469), .ZN(O992));
  NOR2X1 G1145 (.A1(I90), .A2(I91), .ZN(W45));
  NOR2X1 G1146 (.A1(W160), .A2(W56), .ZN(W721));
  NOR2X1 G1147 (.A1(W3243), .A2(W2867), .ZN(W3365));
  NOR2X1 G1148 (.A1(W689), .A2(W244), .ZN(O24));
  NOR2X1 G1149 (.A1(W3272), .A2(W984), .ZN(O994));
  NOR2X1 G1150 (.A1(W1518), .A2(W337), .ZN(O995));
  NOR2X1 G1151 (.A1(W2050), .A2(W536), .ZN(O1562));
  NOR2X1 G1152 (.A1(W3359), .A2(W1235), .ZN(O1576));
  NOR2X1 G1153 (.A1(W2555), .A2(W3249), .ZN(W3372));
  NOR2X1 G1154 (.A1(W3498), .A2(W1514), .ZN(O1573));
  NOR2X1 G1155 (.A1(I110), .A2(I111), .ZN(W55));
  NOR2X1 G1156 (.A1(W615), .A2(I27), .ZN(W712));
  NOR2X1 G1157 (.A1(W2567), .A2(W3324), .ZN(W3375));
  NOR2X1 G1158 (.A1(W550), .A2(W686), .ZN(W710));
  NOR2X1 G1159 (.A1(I112), .A2(I113), .ZN(W56));
  NOR2X1 G1160 (.A1(I170), .A2(I171), .ZN(W85));
  NOR2X1 G1161 (.A1(W349), .A2(W437), .ZN(W668));
  NOR2X1 G1162 (.A1(I162), .A2(I163), .ZN(O0));
  NOR2X1 G1163 (.A1(W714), .A2(W932), .ZN(O1031));
  NOR2X1 G1164 (.A1(W375), .A2(W456), .ZN(W666));
  NOR2X1 G1165 (.A1(W322), .A2(W659), .ZN(W665));
  NOR2X1 G1166 (.A1(I168), .A2(I169), .ZN(W84));
  NOR2X1 G1167 (.A1(W838), .A2(W1512), .ZN(O1033));
  NOR2X1 G1168 (.A1(W1831), .A2(W772), .ZN(O1034));
  NOR2X1 G1169 (.A1(W326), .A2(W3144), .ZN(O1037));
  NOR2X1 G1170 (.A1(I160), .A2(I161), .ZN(W80));
  NOR2X1 G1171 (.A1(W2686), .A2(W3196), .ZN(O1038));
  NOR2X1 G1172 (.A1(W1057), .A2(W463), .ZN(O1040));
  NOR2X1 G1173 (.A1(W591), .A2(W133), .ZN(W658));
  NOR2X1 G1174 (.A1(W3226), .A2(W1144), .ZN(O1041));
  NOR2X1 G1175 (.A1(W2348), .A2(W3344), .ZN(O1547));
  NOR2X1 G1176 (.A1(W538), .A2(W572), .ZN(W655));
  NOR2X1 G1177 (.A1(W307), .A2(W539), .ZN(W654));
  NOR2X1 G1178 (.A1(I174), .A2(I175), .ZN(W87));
  NOR2X1 G1179 (.A1(W3981), .A2(W3741), .ZN(O1546));
  NOR2X1 G1180 (.A1(I79), .A2(W85), .ZN(O19));
  NOR2X1 G1181 (.A1(W3225), .A2(W2095), .ZN(O1559));
  NOR2X1 G1182 (.A1(W506), .A2(W686), .ZN(W3397));
  NOR2X1 G1183 (.A1(W2978), .A2(W2093), .ZN(O1556));
  NOR2X1 G1184 (.A1(W2766), .A2(W651), .ZN(O1555));
  NOR2X1 G1185 (.A1(W3200), .A2(W628), .ZN(O1018));
  NOR2X1 G1186 (.A1(W5), .A2(I150), .ZN(O20));
  NOR2X1 G1187 (.A1(W26), .A2(W193), .ZN(W680));
  NOR2X1 G1188 (.A1(W440), .A2(W1839), .ZN(O1554));
  NOR2X1 G1189 (.A1(W1812), .A2(W792), .ZN(O1020));
  NOR2X1 G1190 (.A1(W2182), .A2(W1304), .ZN(W3357));
  NOR2X1 G1191 (.A1(I146), .A2(I147), .ZN(W73));
  NOR2X1 G1192 (.A1(I34), .A2(I124), .ZN(O18));
  NOR2X1 G1193 (.A1(I150), .A2(I151), .ZN(W75));
  NOR2X1 G1194 (.A1(W63), .A2(W2341), .ZN(O1026));
  NOR2X1 G1195 (.A1(I152), .A2(I153), .ZN(W76));
  NOR2X1 G1196 (.A1(W1412), .A2(W1501), .ZN(O1551));
  NOR2X1 G1197 (.A1(W1146), .A2(W2086), .ZN(W3416));
  NOR2X1 G1198 (.A1(W139), .A2(W49), .ZN(W670));
  NOR2X1 G1199 (.A1(I195), .A2(W664), .ZN(W775));
  NOR2X1 G1200 (.A1(W752), .A2(I28), .ZN(W782));
  NOR2X1 G1201 (.A1(W301), .A2(W721), .ZN(W781));
  NOR2X1 G1202 (.A1(I20), .A2(I21), .ZN(W10));
  NOR2X1 G1203 (.A1(W173), .A2(W274), .ZN(O28));
  NOR2X1 G1204 (.A1(W513), .A2(W23), .ZN(W779));
  NOR2X1 G1205 (.A1(W2974), .A2(I123), .ZN(O1622));
  NOR2X1 G1206 (.A1(W2593), .A2(W3310), .ZN(O1621));
  NOR2X1 G1207 (.A1(I26), .A2(I27), .ZN(W13));
  NOR2X1 G1208 (.A1(W3286), .A2(W1581), .ZN(O953));
  NOR2X1 G1209 (.A1(W1810), .A2(W3584), .ZN(O1624));
  NOR2X1 G1210 (.A1(I30), .A2(I31), .ZN(W15));
  NOR2X1 G1211 (.A1(W361), .A2(W312), .ZN(W774));
  NOR2X1 G1212 (.A1(W430), .A2(I71), .ZN(W773));
  NOR2X1 G1213 (.A1(W647), .A2(W577), .ZN(W772));
  NOR2X1 G1214 (.A1(W3421), .A2(W3822), .ZN(O1614));
  NOR2X1 G1215 (.A1(W1723), .A2(W901), .ZN(O955));
  NOR2X1 G1216 (.A1(W149), .A2(W3341), .ZN(O1611));
  NOR2X1 G1217 (.A1(W133), .A2(W739), .ZN(W768));
  NOR2X1 G1218 (.A1(W248), .A2(W649), .ZN(O1610));
  NOR2X1 G1219 (.A1(W2967), .A2(W2689), .ZN(W3292));
  NOR2X1 G1220 (.A1(W157), .A2(W2509), .ZN(O1630));
  NOR2X1 G1221 (.A1(W1232), .A2(W3666), .ZN(O1629));
  NOR2X1 G1222 (.A1(I6), .A2(I7), .ZN(W3));
  NOR2X1 G1223 (.A1(I8), .A2(I9), .ZN(W4));
  NOR2X1 G1224 (.A1(W2864), .A2(W1234), .ZN(W3289));
  NOR2X1 G1225 (.A1(W480), .A2(W240), .ZN(W796));
  NOR2X1 G1226 (.A1(I10), .A2(I11), .ZN(W5));
  NOR2X1 G1227 (.A1(W2170), .A2(W39), .ZN(W3290));
  NOR2X1 G1228 (.A1(W808), .A2(W1728), .ZN(W3291));
  NOR2X1 G1229 (.A1(I42), .A2(I43), .ZN(W21));
  NOR2X1 G1230 (.A1(W156), .A2(W556), .ZN(W792));
  NOR2X1 G1231 (.A1(I80), .A2(W99), .ZN(W791));
  NOR2X1 G1232 (.A1(I100), .A2(W66), .ZN(O29));
  NOR2X1 G1233 (.A1(I138), .A2(W263), .ZN(W788));
  NOR2X1 G1234 (.A1(W1761), .A2(I12), .ZN(O945));
  NOR2X1 G1235 (.A1(W204), .A2(W135), .ZN(W785));
  NOR2X1 G1236 (.A1(W1325), .A2(W1552), .ZN(O948));
  NOR2X1 G1237 (.A1(W1146), .A2(W2834), .ZN(O949));
  NOR2X1 G1238 (.A1(I70), .A2(I71), .ZN(W35));
  NOR2X1 G1239 (.A1(I66), .A2(I182), .ZN(W748));
  NOR2X1 G1240 (.A1(W179), .A2(W68), .ZN(W747));
  NOR2X1 G1241 (.A1(W485), .A2(W2813), .ZN(O1602));
  NOR2X1 G1242 (.A1(I64), .A2(I65), .ZN(W32));
  NOR2X1 G1243 (.A1(I142), .A2(W815), .ZN(W3339));
  NOR2X1 G1244 (.A1(W106), .A2(W2773), .ZN(O1601));
  NOR2X1 G1245 (.A1(W2078), .A2(W43), .ZN(O980));
  NOR2X1 G1246 (.A1(W3221), .A2(W2168), .ZN(O981));
  NOR2X1 G1247 (.A1(W662), .A2(W125), .ZN(W738));
  NOR2X1 G1248 (.A1(W303), .A2(W595), .ZN(W750));
  NOR2X1 G1249 (.A1(W1848), .A2(W89), .ZN(O984));
  NOR2X1 G1250 (.A1(W2851), .A2(W1990), .ZN(O1597));
  NOR2X1 G1251 (.A1(W97), .A2(W532), .ZN(W733));
  NOR2X1 G1252 (.A1(I74), .A2(I75), .ZN(W37));
  NOR2X1 G1253 (.A1(I40), .A2(W391), .ZN(W731));
  NOR2X1 G1254 (.A1(W1771), .A2(W3031), .ZN(O988));
  NOR2X1 G1255 (.A1(I78), .A2(I79), .ZN(W39));
  NOR2X1 G1256 (.A1(I80), .A2(I81), .ZN(W40));
  NOR2X1 G1257 (.A1(W335), .A2(W3254), .ZN(W3356));
  NOR2X1 G1258 (.A1(I113), .A2(W272), .ZN(W757));
  NOR2X1 G1259 (.A1(W670), .A2(W2897), .ZN(W3310));
  NOR2X1 G1260 (.A1(W2123), .A2(W2990), .ZN(W3313));
  NOR2X1 G1261 (.A1(W3633), .A2(W2019), .ZN(O1608));
  NOR2X1 G1262 (.A1(W2786), .A2(W2544), .ZN(O963));
  NOR2X1 G1263 (.A1(I48), .A2(I49), .ZN(W24));
  NOR2X1 G1264 (.A1(W56), .A2(W78), .ZN(W761));
  NOR2X1 G1265 (.A1(W496), .A2(W65), .ZN(W760));
  NOR2X1 G1266 (.A1(W1351), .A2(W2639), .ZN(W3322));
  NOR2X1 G1267 (.A1(I50), .A2(I51), .ZN(W25));
  NOR2X1 G1268 (.A1(W555), .A2(W268), .ZN(W693));
  NOR2X1 G1269 (.A1(I80), .A2(W705), .ZN(W756));
  NOR2X1 G1270 (.A1(W1935), .A2(W576), .ZN(O967));
  NOR2X1 G1271 (.A1(W189), .A2(I10), .ZN(W754));
  NOR2X1 G1272 (.A1(W194), .A2(W1883), .ZN(O968));
  NOR2X1 G1273 (.A1(W1466), .A2(W2931), .ZN(O1605));
  NOR2X1 G1274 (.A1(I124), .A2(W2254), .ZN(O969));
  NOR2X1 G1275 (.A1(W2964), .A2(W1794), .ZN(W3332));
  NOR2X1 G1276 (.A1(I56), .A2(I57), .ZN(W28));
  NOR2X1 G1277 (.A1(I102), .A2(W27), .ZN(W119));
  NOR2X1 G1278 (.A1(I154), .A2(I46), .ZN(W107));
  NOR2X1 G1279 (.A1(W1988), .A2(W1636), .ZN(O1083));
  NOR2X1 G1280 (.A1(W3161), .A2(I43), .ZN(O1528));
  NOR2X1 G1281 (.A1(W697), .A2(W1775), .ZN(W3458));
  NOR2X1 G1282 (.A1(W2207), .A2(W2189), .ZN(O1057));
  NOR2X1 G1283 (.A1(W298), .A2(W3435), .ZN(W3489));
  NOR2X1 G1284 (.A1(W1659), .A2(W3978), .ZN(O1529));
  NOR2X1 G1285 (.A1(I45), .A2(W62), .ZN(W103));
  NOR2X1 G1286 (.A1(I51), .A2(W3633), .ZN(O1531));
  NOR2X1 G1287 (.A1(W3), .A2(W356), .ZN(W635));
  NOR2X1 G1288 (.A1(W342), .A2(W574), .ZN(W629));
  NOR2X1 G1289 (.A1(W774), .A2(W2390), .ZN(O1533));
  NOR2X1 G1290 (.A1(W334), .A2(W2599), .ZN(O1086));
  NOR2X1 G1291 (.A1(W886), .A2(W284), .ZN(W3494));
  NOR2X1 G1292 (.A1(W484), .A2(W35), .ZN(W600));
  NOR2X1 G1293 (.A1(W508), .A2(I166), .ZN(W599));
  NOR2X1 G1294 (.A1(W356), .A2(W142), .ZN(O1536));
  NOR2X1 G1295 (.A1(I192), .A2(I193), .ZN(W96));
  NOR2X1 G1296 (.A1(W3105), .A2(W2876), .ZN(O1513));
  NOR2X1 G1297 (.A1(W540), .A2(W497), .ZN(W639));
  NOR2X1 G1298 (.A1(W1732), .A2(W1692), .ZN(O1089));
  NOR2X1 G1299 (.A1(W596), .A2(W3289), .ZN(W3981));
  NOR2X1 G1300 (.A1(W504), .A2(W1751), .ZN(O1519));
  NOR2X1 G1301 (.A1(W39), .A2(W3190), .ZN(O1520));
  NOR2X1 G1302 (.A1(W395), .A2(W559), .ZN(W619));
  NOR2X1 G1303 (.A1(W197), .A2(W394), .ZN(O16));
  NOR2X1 G1304 (.A1(W3343), .A2(W1334), .ZN(O1517));
  NOR2X1 G1305 (.A1(I55), .A2(W80), .ZN(W110));
  NOR2X1 G1306 (.A1(W460), .A2(I145), .ZN(W621));
  NOR2X1 G1307 (.A1(W2491), .A2(W1612), .ZN(O1076));
  NOR2X1 G1308 (.A1(I148), .A2(W35), .ZN(W109));
  NOR2X1 G1309 (.A1(W1758), .A2(W2897), .ZN(O1069));
  NOR2X1 G1310 (.A1(W40), .A2(W520), .ZN(W589));
  NOR2X1 G1311 (.A1(W912), .A2(W764), .ZN(O1514));
  NOR2X1 G1312 (.A1(W653), .A2(W2366), .ZN(O1068));
  NOR2X1 G1313 (.A1(W1305), .A2(W1935), .ZN(O1080));
  NOR2X1 G1314 (.A1(W25), .A2(I58), .ZN(W625));
  NOR2X1 G1315 (.A1(W2382), .A2(W2756), .ZN(W3978));
  NOR2X1 G1316 (.A1(W3435), .A2(W317), .ZN(O1081));
  NOR2X1 G1317 (.A1(W2957), .A2(W2926), .ZN(O1067));
  NOR2X1 G1318 (.A1(W171), .A2(W453), .ZN(W3485));
  NOR2X1 G1319 (.A1(W441), .A2(W451), .ZN(W627));
  NOR2X1 G1320 (.A1(W3392), .A2(W3278), .ZN(O1066));
  NOR2X1 G1321 (.A1(W506), .A2(W466), .ZN(W590));
  NOR2X1 G1322 (.A1(W2832), .A2(W2946), .ZN(W3435));
  NOR2X1 G1323 (.A1(W552), .A2(W279), .ZN(W652));
  NOR2X1 G1324 (.A1(W263), .A2(I151), .ZN(O1092));
  NOR2X1 G1325 (.A1(I178), .A2(I179), .ZN(W89));
  NOR2X1 G1326 (.A1(W1831), .A2(W2708), .ZN(O1047));
  NOR2X1 G1327 (.A1(W2961), .A2(W1904), .ZN(W3442));
  NOR2X1 G1328 (.A1(I180), .A2(I181), .ZN(W90));
  NOR2X1 G1329 (.A1(W592), .A2(W370), .ZN(W653));
  NOR2X1 G1330 (.A1(W2608), .A2(W321), .ZN(W3438));
  NOR2X1 G1331 (.A1(I70), .A2(W65), .ZN(W122));
  NOR2X1 G1332 (.A1(W2205), .A2(W388), .ZN(O1090));
  NOR2X1 G1333 (.A1(W376), .A2(I109), .ZN(W651));
  NOR2X1 G1334 (.A1(I184), .A2(I185), .ZN(W92));
  NOR2X1 G1335 (.A1(I190), .A2(I191), .ZN(W95));
  NOR2X1 G1336 (.A1(I146), .A2(W74), .ZN(W124));
  NOR2X1 G1337 (.A1(W379), .A2(W350), .ZN(W593));
  NANDX1 G1338 (.A1(W1213), .A2(W2290), .ZN(W2411));
  NANDX1 G1339 (.A1(W854), .A2(W1594), .ZN(W2065));
  NANDX1 G1340 (.A1(W566), .A2(W1308), .ZN(O431));
  NANDX1 G1341 (.A1(W1973), .A2(W290), .ZN(W2409));
  NANDX1 G1342 (.A1(W1989), .A2(W1592), .ZN(O1515));
  NANDX1 G1343 (.A1(W1666), .A2(W29), .ZN(O279));
  NANDX1 G1344 (.A1(W329), .A2(W1534), .ZN(O363));
  NANDX1 G1345 (.A1(I95), .A2(W1332), .ZN(O294));
  NANDX1 G1346 (.A1(W106), .A2(W2306), .ZN(O429));
  NANDX1 G1347 (.A1(W1433), .A2(I142), .ZN(W2245));
  NANDX1 G1348 (.A1(W177), .A2(W915), .ZN(O456));
  NANDX1 G1349 (.A1(W2002), .A2(W1819), .ZN(O1506));
  NANDX1 G1350 (.A1(W816), .A2(W1755), .ZN(W2064));
  NANDX1 G1351 (.A1(W3705), .A2(W2956), .ZN(O1398));
  NANDX1 G1352 (.A1(W365), .A2(I191), .ZN(O1606));
  NANDX1 G1353 (.A1(W257), .A2(W1289), .ZN(O1487));
  NANDX1 G1354 (.A1(W900), .A2(I16), .ZN(O346));
  NANDX1 G1355 (.A1(W2050), .A2(W807), .ZN(W2214));
  NANDX1 G1356 (.A1(W1465), .A2(W2234), .ZN(W2240));
  NANDX1 G1357 (.A1(W691), .A2(W1104), .ZN(O344));
  NANDX1 G1358 (.A1(W2897), .A2(W1542), .ZN(O1395));
  NANDX1 G1359 (.A1(W1347), .A2(W1944), .ZN(O1600));
  NANDX1 G1360 (.A1(W1371), .A2(W567), .ZN(W2259));
  NANDX1 G1361 (.A1(W1631), .A2(W3432), .ZN(O1409));
  NANDX1 G1362 (.A1(W1473), .A2(W1905), .ZN(O334));
  NANDX1 G1363 (.A1(W1147), .A2(W369), .ZN(W2079));
  NANDX1 G1364 (.A1(W615), .A2(W1379), .ZN(W2394));
  NANDX1 G1365 (.A1(W1931), .A2(W1466), .ZN(O425));
  NANDX1 G1366 (.A1(W17), .A2(W818), .ZN(W2396));
  NANDX1 G1367 (.A1(W1946), .A2(W2182), .ZN(O1588));
  NANDX1 G1368 (.A1(W476), .A2(W1906), .ZN(O1407));
  NANDX1 G1369 (.A1(W1591), .A2(W1719), .ZN(W2258));
  NANDX1 G1370 (.A1(I197), .A2(W1202), .ZN(O335));
  NANDX1 G1371 (.A1(W2041), .A2(W1644), .ZN(O366));
  NANDX1 G1372 (.A1(I192), .A2(W1162), .ZN(W2075));
  NANDX1 G1373 (.A1(I70), .A2(W1079), .ZN(W2251));
  NANDX1 G1374 (.A1(W97), .A2(W2194), .ZN(O1509));
  NANDX1 G1375 (.A1(W279), .A2(W1564), .ZN(O428));
  NANDX1 G1376 (.A1(W863), .A2(W1890), .ZN(O365));
  NANDX1 G1377 (.A1(W539), .A2(W1055), .ZN(O296));
  NANDX1 G1378 (.A1(W1893), .A2(W2148), .ZN(O336));
  NANDX1 G1379 (.A1(W1732), .A2(W1224), .ZN(O338));
  NANDX1 G1380 (.A1(W611), .A2(W444), .ZN(O1403));
  NANDX1 G1381 (.A1(W2033), .A2(W1937), .ZN(O295));
  NANDX1 G1382 (.A1(W2534), .A2(W289), .ZN(O1603));
  NANDX1 G1383 (.A1(W2396), .A2(W2369), .ZN(W2403));
  NANDX1 G1384 (.A1(W3560), .A2(W525), .ZN(O1369));
  NANDX1 G1385 (.A1(W707), .A2(W1701), .ZN(W2070));
  NANDX1 G1386 (.A1(W193), .A2(W1516), .ZN(W2194));
  NANDX1 G1387 (.A1(W1872), .A2(W1536), .ZN(W3854));
  NANDX1 G1388 (.A1(W1957), .A2(W1482), .ZN(O457));
  NANDX1 G1389 (.A1(W1330), .A2(W999), .ZN(O1604));
  NANDX1 G1390 (.A1(W1796), .A2(W1335), .ZN(W2443));
  NANDX1 G1391 (.A1(I138), .A2(W902), .ZN(W2232));
  NANDX1 G1392 (.A1(W1740), .A2(W87), .ZN(W2217));
  NANDX1 G1393 (.A1(I84), .A2(W2935), .ZN(O1613));
  NANDX1 G1394 (.A1(W210), .A2(W1907), .ZN(O447));
  NANDX1 G1395 (.A1(W972), .A2(W474), .ZN(W2230));
  NANDX1 G1396 (.A1(W2207), .A2(W885), .ZN(O453));
  NANDX1 G1397 (.A1(W765), .A2(W3140), .ZN(O1493));
  NANDX1 G1398 (.A1(W1200), .A2(W1204), .ZN(O1627));
  NANDX1 G1399 (.A1(W2043), .A2(W1754), .ZN(W2438));
  NANDX1 G1400 (.A1(I8), .A2(W936), .ZN(W2439));
  NANDX1 G1401 (.A1(W3609), .A2(W257), .ZN(O1499));
  NANDX1 G1402 (.A1(W1398), .A2(W2122), .ZN(O356));
  NANDX1 G1403 (.A1(W1034), .A2(W1093), .ZN(W2441));
  NANDX1 G1404 (.A1(W1783), .A2(W26), .ZN(O1494));
  NANDX1 G1405 (.A1(W67), .A2(W114), .ZN(W2442));
  NANDX1 G1406 (.A1(W1546), .A2(W2134), .ZN(W2205));
  NANDX1 G1407 (.A1(W1047), .A2(W3088), .ZN(O1375));
  NANDX1 G1408 (.A1(W755), .A2(W245), .ZN(O1619));
  NANDX1 G1409 (.A1(W1687), .A2(W391), .ZN(O1626));
  NANDX1 G1410 (.A1(W800), .A2(W446), .ZN(W2445));
  NANDX1 G1411 (.A1(W958), .A2(I153), .ZN(W2446));
  NANDX1 G1412 (.A1(W232), .A2(W209), .ZN(W2226));
  NANDX1 G1413 (.A1(W1504), .A2(W1541), .ZN(O1511));
  NANDX1 G1414 (.A1(W1979), .A2(W771), .ZN(O286));
  NANDX1 G1415 (.A1(W2207), .A2(W1883), .ZN(O350));
  NANDX1 G1416 (.A1(W731), .A2(W1880), .ZN(O351));
  NANDX1 G1417 (.A1(W615), .A2(W1388), .ZN(W2224));
  NANDX1 G1418 (.A1(W2548), .A2(W2823), .ZN(O1512));
  NANDX1 G1419 (.A1(W555), .A2(W339), .ZN(O285));
  NANDX1 G1420 (.A1(W449), .A2(W30), .ZN(O352));
  NANDX1 G1421 (.A1(W3748), .A2(W1851), .ZN(O1389));
  NANDX1 G1422 (.A1(W3089), .A2(W1635), .ZN(O1488));
  NANDX1 G1423 (.A1(W2336), .A2(W3168), .ZN(O1504));
  NANDX1 G1424 (.A1(W902), .A2(W291), .ZN(O348));
  NANDX1 G1425 (.A1(W329), .A2(W3332), .ZN(O1392));
  NANDX1 G1426 (.A1(W1851), .A2(W2400), .ZN(O1501));
  NANDX1 G1427 (.A1(W2551), .A2(W2324), .ZN(O1391));
  NANDX1 G1428 (.A1(W2105), .A2(W1397), .ZN(O339));
  NANDX1 G1429 (.A1(W430), .A2(W1615), .ZN(O437));
  NANDX1 G1430 (.A1(W145), .A2(W1932), .ZN(W2043));
  NANDX1 G1431 (.A1(W1233), .A2(W922), .ZN(W2198));
  NANDX1 G1432 (.A1(W327), .A2(W107), .ZN(O438));
  NANDX1 G1433 (.A1(W1276), .A2(W557), .ZN(O1491));
  NANDX1 G1434 (.A1(W554), .A2(W3489), .ZN(O1607));
  NANDX1 G1435 (.A1(W1741), .A2(W489), .ZN(O455));
  NANDX1 G1436 (.A1(W2612), .A2(W597), .ZN(O1628));
  NANDX1 G1437 (.A1(W1710), .A2(W896), .ZN(W2059));
  NANDX1 G1438 (.A1(W610), .A2(W3290), .ZN(O1388));
  NANDX1 G1439 (.A1(W3039), .A2(W55), .ZN(O1386));
  NANDX1 G1440 (.A1(W66), .A2(W1995), .ZN(W2200));
  NANDX1 G1441 (.A1(W2109), .A2(W1563), .ZN(W2234));
  NANDX1 G1442 (.A1(W974), .A2(W2893), .ZN(O1383));
  NANDX1 G1443 (.A1(W155), .A2(W1897), .ZN(O341));
  NANDX1 G1444 (.A1(W209), .A2(W1677), .ZN(O442));
  NANDX1 G1445 (.A1(W2082), .A2(I122), .ZN(W2433));
  NANDX1 G1446 (.A1(W297), .A2(I135), .ZN(O1371));
  NANDX1 G1447 (.A1(W933), .A2(W3352), .ZN(O1609));
  NANDX1 G1448 (.A1(W1263), .A2(W2525), .ZN(O1492));
  NANDX1 G1449 (.A1(W129), .A2(W565), .ZN(O287));
  NANDX1 G1450 (.A1(W1759), .A2(W1340), .ZN(W2434));
  NANDX1 G1451 (.A1(W1103), .A2(W233), .ZN(O446));
  NANDX1 G1452 (.A1(W218), .A2(W2605), .ZN(O1431));
  NANDX1 G1453 (.A1(W353), .A2(W1752), .ZN(O313));
  NANDX1 G1454 (.A1(I120), .A2(W566), .ZN(O1430));
  NANDX1 G1455 (.A1(W125), .A2(I31), .ZN(O328));
  NANDX1 G1456 (.A1(I176), .A2(W1333), .ZN(O314));
  NANDX1 G1457 (.A1(W1181), .A2(W251), .ZN(O377));
  NANDX1 G1458 (.A1(W1532), .A2(W690), .ZN(W2132));
  NANDX1 G1459 (.A1(W1520), .A2(W1038), .ZN(O1534));
  NANDX1 G1460 (.A1(W2421), .A2(W2997), .ZN(O1535));
  NANDX1 G1461 (.A1(W3165), .A2(W496), .ZN(O1561));
  NANDX1 G1462 (.A1(W19), .A2(W2149), .ZN(O381));
  NANDX1 G1463 (.A1(W1975), .A2(W1877), .ZN(W2286));
  NANDX1 G1464 (.A1(W1922), .A2(W909), .ZN(W2331));
  NANDX1 G1465 (.A1(W1430), .A2(W300), .ZN(W2287));
  NANDX1 G1466 (.A1(I171), .A2(W505), .ZN(O382));
  NANDX1 G1467 (.A1(I182), .A2(W1809), .ZN(W2330));
  NANDX1 G1468 (.A1(W666), .A2(W3755), .ZN(O1553));
  NANDX1 G1469 (.A1(W1134), .A2(W112), .ZN(O318));
  NANDX1 G1470 (.A1(W1341), .A2(W1471), .ZN(O312));
  NANDX1 G1471 (.A1(W58), .A2(W1748), .ZN(O311));
  NANDX1 G1472 (.A1(W730), .A2(W559), .ZN(W3886));
  NANDX1 G1473 (.A1(W407), .A2(W933), .ZN(O1564));
  NANDX1 G1474 (.A1(W2979), .A2(W3886), .ZN(O1425));
  NANDX1 G1475 (.A1(W353), .A2(W517), .ZN(O1426));
  NANDX1 G1476 (.A1(W2924), .A2(W2260), .ZN(O1532));
  NANDX1 G1477 (.A1(W115), .A2(W1623), .ZN(O1508));
  NANDX1 G1478 (.A1(W635), .A2(W208), .ZN(W2126));
  NANDX1 G1479 (.A1(W1035), .A2(W1668), .ZN(O396));
  NANDX1 G1480 (.A1(W1205), .A2(W460), .ZN(W2128));
  NANDX1 G1481 (.A1(W710), .A2(W1397), .ZN(O329));
  NANDX1 G1482 (.A1(W1773), .A2(W663), .ZN(O1454));
  NANDX1 G1483 (.A1(I158), .A2(W291), .ZN(O401));
  NANDX1 G1484 (.A1(W107), .A2(W77), .ZN(O376));
  NANDX1 G1485 (.A1(W1613), .A2(W2636), .ZN(O1429));
  NANDX1 G1486 (.A1(W597), .A2(W988), .ZN(W2280));
  NANDX1 G1487 (.A1(W922), .A2(W914), .ZN(W2302));
  NANDX1 G1488 (.A1(W2594), .A2(W2081), .ZN(O1443));
  NANDX1 G1489 (.A1(W3999), .A2(W1555), .ZN(O1549));
  NANDX1 G1490 (.A1(W1377), .A2(W344), .ZN(O1542));
  NANDX1 G1491 (.A1(W1406), .A2(W1292), .ZN(O1548));
  NANDX1 G1492 (.A1(W588), .A2(W2121), .ZN(W2162));
  NANDX1 G1493 (.A1(W429), .A2(W1322), .ZN(O321));
  NANDX1 G1494 (.A1(W936), .A2(W1050), .ZN(W2161));
  NANDX1 G1495 (.A1(W1869), .A2(W593), .ZN(W2154));
  NANDX1 G1496 (.A1(W950), .A2(W925), .ZN(O1540));
  NANDX1 G1497 (.A1(W1883), .A2(I58), .ZN(O1453));
  NANDX1 G1498 (.A1(W1332), .A2(W726), .ZN(W2314));
  NANDX1 G1499 (.A1(W688), .A2(W961), .ZN(W2160));
  NANDX1 G1500 (.A1(W1190), .A2(W119), .ZN(O391));
  NANDX1 G1501 (.A1(W1265), .A2(W1940), .ZN(O1452));
  NANDX1 G1502 (.A1(W244), .A2(W530), .ZN(O1448));
  NANDX1 G1503 (.A1(W2294), .A2(W1894), .ZN(O389));
  NANDX1 G1504 (.A1(W161), .A2(W1961), .ZN(W2167));
  NANDX1 G1505 (.A1(I27), .A2(W317), .ZN(W2289));
  NANDX1 G1506 (.A1(W1614), .A2(W482), .ZN(W2327));
  NANDX1 G1507 (.A1(W472), .A2(I55), .ZN(O1539));
  NANDX1 G1508 (.A1(W3404), .A2(W482), .ZN(O1439));
  NANDX1 G1509 (.A1(W1083), .A2(W978), .ZN(W2168));
  NANDX1 G1510 (.A1(W1934), .A2(I49), .ZN(W2141));
  NANDX1 G1511 (.A1(W2077), .A2(W1674), .ZN(O1552));
  NANDX1 G1512 (.A1(W1389), .A2(W926), .ZN(W2143));
  NANDX1 G1513 (.A1(W1869), .A2(W2019), .ZN(W2352));
  NANDX1 G1514 (.A1(W1029), .A2(W1837), .ZN(W2166));
  NANDX1 G1515 (.A1(W929), .A2(W1889), .ZN(W2290));
  NANDX1 G1516 (.A1(I21), .A2(W924), .ZN(W2147));
  NANDX1 G1517 (.A1(W3214), .A2(W2320), .ZN(O1550));
  NANDX1 G1518 (.A1(I3), .A2(W386), .ZN(O383));
  NANDX1 G1519 (.A1(W3614), .A2(W2846), .ZN(O1442));
  NANDX1 G1520 (.A1(W511), .A2(W1775), .ZN(W2322));
  NANDX1 G1521 (.A1(W1192), .A2(W1979), .ZN(O1585));
  NANDX1 G1522 (.A1(W3802), .A2(W3196), .ZN(O1587));
  NANDX1 G1523 (.A1(W634), .A2(W1405), .ZN(W2094));
  NANDX1 G1524 (.A1(W549), .A2(W2132), .ZN(W2382));
  NANDX1 G1525 (.A1(W1030), .A2(I169), .ZN(W2380));
  NANDX1 G1526 (.A1(W2210), .A2(W1389), .ZN(O1521));
  NANDX1 G1527 (.A1(W1079), .A2(W1534), .ZN(O302));
  NANDX1 G1528 (.A1(W1371), .A2(W468), .ZN(W2269));
  NANDX1 G1529 (.A1(W242), .A2(W3056), .ZN(O1586));
  NANDX1 G1530 (.A1(W197), .A2(W2091), .ZN(O1413));
  NANDX1 G1531 (.A1(W1686), .A2(W3382), .ZN(O1583));
  NANDX1 G1532 (.A1(W1759), .A2(W2259), .ZN(O1582));
  NANDX1 G1533 (.A1(W2822), .A2(W2548), .ZN(O1527));
  NANDX1 G1534 (.A1(W3978), .A2(W2089), .ZN(O1581));
  NANDX1 G1535 (.A1(W1917), .A2(W702), .ZN(W2105));
  NANDX1 G1536 (.A1(W1357), .A2(W1667), .ZN(W2376));
  NANDX1 G1537 (.A1(W789), .A2(W2294), .ZN(W2375));
  NANDX1 G1538 (.A1(W1669), .A2(W1210), .ZN(W2106));
  NANDX1 G1539 (.A1(W1719), .A2(W59), .ZN(W2089));
  NANDX1 G1540 (.A1(W522), .A2(W1441), .ZN(W2260));
  NANDX1 G1541 (.A1(W1321), .A2(W1942), .ZN(W2186));
  NANDX1 G1542 (.A1(W1348), .A2(W845), .ZN(O298));
  NANDX1 G1543 (.A1(W1454), .A2(W512), .ZN(O299));
  NANDX1 G1544 (.A1(W1111), .A2(W543), .ZN(W2653));
  NANDX1 G1545 (.A1(W1421), .A2(W1134), .ZN(W2390));
  NANDX1 G1546 (.A1(W3854), .A2(W359), .ZN(O1594));
  NANDX1 G1547 (.A1(W3379), .A2(W936), .ZN(O1475));
  NANDX1 G1548 (.A1(W2559), .A2(W2650), .ZN(O1472));
  NANDX1 G1549 (.A1(W52), .A2(W2200), .ZN(W2261));
  NANDX1 G1550 (.A1(W1696), .A2(W942), .ZN(O368));
  NANDX1 G1551 (.A1(W3380), .A2(W3123), .ZN(O1591));
  NANDX1 G1552 (.A1(W4044), .A2(W22), .ZN(O1589));
  NANDX1 G1553 (.A1(W867), .A2(W513), .ZN(O420));
  NANDX1 G1554 (.A1(W1824), .A2(W879), .ZN(O390));
  NANDX1 G1555 (.A1(W2067), .A2(W1092), .ZN(W2385));
  NANDX1 G1556 (.A1(W596), .A2(W2226), .ZN(O404));
  NANDX1 G1557 (.A1(W1930), .A2(W381), .ZN(O1571));
  NANDX1 G1558 (.A1(W1433), .A2(W876), .ZN(O1420));
  NANDX1 G1559 (.A1(W3704), .A2(W3414), .ZN(O1462));
  NANDX1 G1560 (.A1(W867), .A2(W2933), .ZN(O1421));
  NANDX1 G1561 (.A1(W324), .A2(I176), .ZN(W2354));
  NANDX1 G1562 (.A1(W2167), .A2(W3214), .ZN(O1422));
  NANDX1 G1563 (.A1(W508), .A2(W2921), .ZN(O1423));
  NANDX1 G1564 (.A1(W1120), .A2(W1796), .ZN(W2120));
  NANDX1 G1565 (.A1(W2257), .A2(W399), .ZN(O373));
  NANDX1 G1566 (.A1(I78), .A2(W1032), .ZN(W2122));
  NANDX1 G1567 (.A1(W433), .A2(W1655), .ZN(O1461));
  NANDX1 G1568 (.A1(W3279), .A2(W1377), .ZN(O1456));
  NANDX1 G1569 (.A1(W493), .A2(W1095), .ZN(O374));
  NANDX1 G1570 (.A1(W2842), .A2(W3952), .ZN(O1530));
  NANDX1 G1571 (.A1(W380), .A2(W1562), .ZN(O310));
  NANDX1 G1572 (.A1(W1216), .A2(W3622), .ZN(O1566));
  NANDX1 G1573 (.A1(W833), .A2(W3731), .ZN(O1416));
  NANDX1 G1574 (.A1(W803), .A2(W1141), .ZN(W2369));
  NANDX1 G1575 (.A1(W1460), .A2(W328), .ZN(O1471));
  NANDX1 G1576 (.A1(W783), .A2(W483), .ZN(W2367));
  NANDX1 G1577 (.A1(W167), .A2(W44), .ZN(O305));
  NANDX1 G1578 (.A1(W3105), .A2(W175), .ZN(O1575));
  NANDX1 G1579 (.A1(W473), .A2(W2094), .ZN(O306));
  NANDX1 G1580 (.A1(W213), .A2(W1714), .ZN(W2366));
  NANDX1 G1581 (.A1(W727), .A2(W1089), .ZN(W2272));
  NANDX1 G1582 (.A1(W1183), .A2(W1842), .ZN(W2082));
  NANDX1 G1583 (.A1(W1253), .A2(W1169), .ZN(O411));
  NANDX1 G1584 (.A1(W367), .A2(W1180), .ZN(O410));
  NANDX1 G1585 (.A1(W1944), .A2(W1538), .ZN(W2360));
  NANDX1 G1586 (.A1(W3334), .A2(W3128), .ZN(O1470));
  NANDX1 G1587 (.A1(W910), .A2(W1150), .ZN(O407));
  NANDX1 G1588 (.A1(W1676), .A2(W151), .ZN(W2357));
  NANDX1 G1589 (.A1(W2147), .A2(W1382), .ZN(O406));
  NANDX1 G1590 (.A1(W2150), .A2(W2214), .ZN(O757));
  NANDX1 G1591 (.A1(W1192), .A2(W252), .ZN(W3037));
  NANDX1 G1592 (.A1(W2482), .A2(W1330), .ZN(W3035));
  NANDX1 G1593 (.A1(W2580), .A2(W1730), .ZN(O766));
  NANDX1 G1594 (.A1(W993), .A2(W46), .ZN(O1051));
  NANDX1 G1595 (.A1(W1401), .A2(W2657), .ZN(W3031));
  NANDX1 G1596 (.A1(W97), .A2(W2825), .ZN(O1053));
  NANDX1 G1597 (.A1(W998), .A2(W2826), .ZN(O1054));
  NANDX1 G1598 (.A1(W287), .A2(W1002), .ZN(W3027));
  NANDX1 G1599 (.A1(W1282), .A2(W2286), .ZN(O761));
  NANDX1 G1600 (.A1(W1286), .A2(W2245), .ZN(O759));
  NANDX1 G1601 (.A1(W2152), .A2(W2081), .ZN(W3451));
  NANDX1 G1602 (.A1(W2632), .A2(W643), .ZN(O1056));
  NANDX1 G1603 (.A1(W163), .A2(W2327), .ZN(W3022));
  NANDX1 G1604 (.A1(W3089), .A2(W2632), .ZN(O1048));
  NANDX1 G1605 (.A1(W1897), .A2(W1668), .ZN(W3015));
  NANDX1 G1606 (.A1(W325), .A2(W1135), .ZN(O1063));
  NANDX1 G1607 (.A1(W2466), .A2(W2737), .ZN(O1070));
  NANDX1 G1608 (.A1(W779), .A2(W2322), .ZN(O750));
  NANDX1 G1609 (.A1(W238), .A2(W739), .ZN(O744));
  NANDX1 G1610 (.A1(W1148), .A2(W1307), .ZN(O743));
  NANDX1 G1611 (.A1(W902), .A2(W1459), .ZN(W3472));
  NANDX1 G1612 (.A1(W1380), .A2(W1086), .ZN(W2992));
  NANDX1 G1613 (.A1(W1810), .A2(W361), .ZN(O739));
  NANDX1 G1614 (.A1(W1545), .A2(W2272), .ZN(W2990));
  NANDX1 G1615 (.A1(W2084), .A2(W2827), .ZN(O1072));
  NANDX1 G1616 (.A1(W2939), .A2(W592), .ZN(W2986));
  NANDX1 G1617 (.A1(W2544), .A2(W331), .ZN(O1074));
  NANDX1 G1618 (.A1(W1379), .A2(W1515), .ZN(O1633));
  NANDX1 G1619 (.A1(W2494), .A2(W1889), .ZN(O796));
  NANDX1 G1620 (.A1(W1030), .A2(W665), .ZN(W3088));
  NANDX1 G1621 (.A1(W2154), .A2(W2764), .ZN(O795));
  NANDX1 G1622 (.A1(I20), .A2(W304), .ZN(O1028));
  NANDX1 G1623 (.A1(W2160), .A2(W358), .ZN(W3085));
  NANDX1 G1624 (.A1(W1573), .A2(W1223), .ZN(O793));
  NANDX1 G1625 (.A1(W2583), .A2(W1429), .ZN(O1030));
  NANDX1 G1626 (.A1(W148), .A2(W2606), .ZN(W3081));
  NANDX1 G1627 (.A1(W1772), .A2(W529), .ZN(W3072));
  NANDX1 G1628 (.A1(W2624), .A2(W2402), .ZN(W3421));
  NANDX1 G1629 (.A1(W2385), .A2(W2360), .ZN(O782));
  NANDX1 G1630 (.A1(W3015), .A2(W2986), .ZN(W3066));
  NANDX1 G1631 (.A1(W2481), .A2(W2560), .ZN(O780));
  NANDX1 G1632 (.A1(W1596), .A2(W1183), .ZN(O736));
  NANDX1 G1633 (.A1(I102), .A2(W1601), .ZN(W3432));
  NANDX1 G1634 (.A1(W40), .A2(W1604), .ZN(W3058));
  NANDX1 G1635 (.A1(W384), .A2(W408), .ZN(W3054));
  NANDX1 G1636 (.A1(W3339), .A2(W2339), .ZN(O1042));
  NANDX1 G1637 (.A1(W511), .A2(W2985), .ZN(O773));
  NANDX1 G1638 (.A1(W1043), .A2(W3404), .ZN(O1043));
  NANDX1 G1639 (.A1(W3313), .A2(W965), .ZN(O1044));
  NANDX1 G1640 (.A1(W1348), .A2(W1518), .ZN(W3047));
  NANDX1 G1641 (.A1(W1575), .A2(W1255), .ZN(O772));
  NANDX1 G1642 (.A1(W176), .A2(W800), .ZN(O1045));
  NANDX1 G1643 (.A1(W3084), .A2(W1733), .ZN(O1046));
  NANDX1 G1644 (.A1(W3407), .A2(W944), .ZN(W3443));
  NANDX1 G1645 (.A1(W522), .A2(W1831), .ZN(W3039));
  NANDX1 G1646 (.A1(W2373), .A2(W2455), .ZN(W2909));
  NANDX1 G1647 (.A1(W2253), .A2(W1294), .ZN(W2922));
  NANDX1 G1648 (.A1(W2044), .A2(W908), .ZN(W2919));
  NANDX1 G1649 (.A1(W1157), .A2(W2724), .ZN(W2918));
  NANDX1 G1650 (.A1(W3128), .A2(W1690), .ZN(W3525));
  NANDX1 G1651 (.A1(W1931), .A2(W2105), .ZN(O1114));
  NANDX1 G1652 (.A1(W2185), .A2(W1262), .ZN(O704));
  NANDX1 G1653 (.A1(W260), .A2(W709), .ZN(O703));
  NANDX1 G1654 (.A1(I182), .A2(W942), .ZN(W3528));
  NANDX1 G1655 (.A1(I56), .A2(W1896), .ZN(W2915));
  NANDX1 G1656 (.A1(W413), .A2(W2520), .ZN(O1115));
  NANDX1 G1657 (.A1(W225), .A2(W2823), .ZN(O702));
  NANDX1 G1658 (.A1(W2945), .A2(W3053), .ZN(O1116));
  NANDX1 G1659 (.A1(W2497), .A2(W2051), .ZN(O701));
  NANDX1 G1660 (.A1(W227), .A2(W2763), .ZN(W2926));
  NANDX1 G1661 (.A1(W1422), .A2(W2011), .ZN(W2907));
  NANDX1 G1662 (.A1(W2331), .A2(W2266), .ZN(W2906));
  NANDX1 G1663 (.A1(W484), .A2(W810), .ZN(O698));
  NANDX1 G1664 (.A1(W1325), .A2(W27), .ZN(O1118));
  NANDX1 G1665 (.A1(W796), .A2(I110), .ZN(O1121));
  NANDX1 G1666 (.A1(W2070), .A2(W1884), .ZN(O696));
  NANDX1 G1667 (.A1(W1784), .A2(W1957), .ZN(W2902));
  NANDX1 G1668 (.A1(W1834), .A2(W392), .ZN(O1123));
  NANDX1 G1669 (.A1(W398), .A2(W1650), .ZN(O1126));
  NANDX1 G1670 (.A1(W1980), .A2(W1478), .ZN(O1127));
  NANDX1 G1671 (.A1(W2881), .A2(W549), .ZN(W2900));
  NANDX1 G1672 (.A1(W1885), .A2(W2860), .ZN(O694));
  NANDX1 G1673 (.A1(W2162), .A2(W791), .ZN(O693));
  NANDX1 G1674 (.A1(W1081), .A2(W293), .ZN(O718));
  NANDX1 G1675 (.A1(W388), .A2(W1927), .ZN(O1075));
  NANDX1 G1676 (.A1(W1970), .A2(W1582), .ZN(O1077));
  NANDX1 G1677 (.A1(W360), .A2(W184), .ZN(O1078));
  NANDX1 G1678 (.A1(W3367), .A2(W1865), .ZN(O1079));
  NANDX1 G1679 (.A1(W2403), .A2(W2772), .ZN(W2967));
  NANDX1 G1680 (.A1(W2128), .A2(W2510), .ZN(W3487));
  NANDX1 G1681 (.A1(W1228), .A2(W2446), .ZN(O722));
  NANDX1 G1682 (.A1(W2074), .A2(W123), .ZN(O721));
  NANDX1 G1683 (.A1(W2394), .A2(W2295), .ZN(O1085));
  NANDX1 G1684 (.A1(W3292), .A2(W2657), .ZN(W3492));
  NANDX1 G1685 (.A1(W1150), .A2(W1040), .ZN(O1087));
  NANDX1 G1686 (.A1(W1086), .A2(W669), .ZN(O1088));
  NANDX1 G1687 (.A1(W2223), .A2(W1225), .ZN(O719));
  NANDX1 G1688 (.A1(W1100), .A2(W1300), .ZN(W3414));
  NANDX1 G1689 (.A1(W2026), .A2(W160), .ZN(W3500));
  NANDX1 G1690 (.A1(W1424), .A2(W138), .ZN(W2946));
  NANDX1 G1691 (.A1(W3099), .A2(W723), .ZN(O1091));
  NANDX1 G1692 (.A1(W1010), .A2(W573), .ZN(O713));
  NANDX1 G1693 (.A1(W2195), .A2(W1571), .ZN(O1096));
  NANDX1 G1694 (.A1(W3049), .A2(W1559), .ZN(O1100));
  NANDX1 G1695 (.A1(W2388), .A2(W236), .ZN(W2938));
  NANDX1 G1696 (.A1(W594), .A2(W1747), .ZN(O710));
  NANDX1 G1697 (.A1(W603), .A2(W664), .ZN(W2934));
  NANDX1 G1698 (.A1(W193), .A2(W2337), .ZN(O709));
  NANDX1 G1699 (.A1(W534), .A2(W1776), .ZN(W2931));
  NANDX1 G1700 (.A1(W1744), .A2(W1378), .ZN(W2930));
  NANDX1 G1701 (.A1(W982), .A2(W799), .ZN(O1109));
  NANDX1 G1702 (.A1(W2370), .A2(W416), .ZN(O886));
  NANDX1 G1703 (.A1(W1969), .A2(W1773), .ZN(O966));
  NANDX1 G1704 (.A1(W2702), .A2(W1475), .ZN(W3323));
  NANDX1 G1705 (.A1(W606), .A2(W2608), .ZN(O898));
  NANDX1 G1706 (.A1(W1515), .A2(W2007), .ZN(W3230));
  NANDX1 G1707 (.A1(W2333), .A2(W3089), .ZN(O897));
  NANDX1 G1708 (.A1(W395), .A2(W388), .ZN(O896));
  NANDX1 G1709 (.A1(W624), .A2(W1522), .ZN(W3226));
  NANDX1 G1710 (.A1(W2502), .A2(W688), .ZN(O894));
  NANDX1 G1711 (.A1(W187), .A2(W860), .ZN(O890));
  NANDX1 G1712 (.A1(W2335), .A2(W2791), .ZN(O974));
  NANDX1 G1713 (.A1(W2589), .A2(W1355), .ZN(W3334));
  NANDX1 G1714 (.A1(W578), .A2(W2722), .ZN(O887));
  NANDX1 G1715 (.A1(W2927), .A2(W551), .ZN(O976));
  NANDX1 G1716 (.A1(W3187), .A2(W2830), .ZN(O905));
  NANDX1 G1717 (.A1(W118), .A2(W2937), .ZN(O977));
  NANDX1 G1718 (.A1(W421), .A2(W1664), .ZN(W3341));
  NANDX1 G1719 (.A1(W2728), .A2(W3060), .ZN(O882));
  NANDX1 G1720 (.A1(W1435), .A2(I28), .ZN(O877));
  NANDX1 G1721 (.A1(W1304), .A2(W508), .ZN(W3344));
  NANDX1 G1722 (.A1(W3341), .A2(W489), .ZN(O982));
  NANDX1 G1723 (.A1(W2945), .A2(W1652), .ZN(O983));
  NANDX1 G1724 (.A1(W753), .A2(W410), .ZN(O872));
  NANDX1 G1725 (.A1(W415), .A2(W1045), .ZN(O985));
  NANDX1 G1726 (.A1(W320), .A2(I154), .ZN(W3193));
  NANDX1 G1727 (.A1(W2178), .A2(W3088), .ZN(O870));
  NANDX1 G1728 (.A1(W379), .A2(W17), .ZN(O987));
  NANDX1 G1729 (.A1(W389), .A2(W2501), .ZN(W3353));
  NANDX1 G1730 (.A1(W2659), .A2(W479), .ZN(O921));
  NANDX1 G1731 (.A1(W2304), .A2(W563), .ZN(O940));
  NANDX1 G1732 (.A1(W504), .A2(W2165), .ZN(O939));
  NANDX1 G1733 (.A1(W2434), .A2(W1669), .ZN(O938));
  NANDX1 G1734 (.A1(W1223), .A2(W2625), .ZN(O943));
  NANDX1 G1735 (.A1(W504), .A2(W1740), .ZN(O936));
  NANDX1 G1736 (.A1(W2448), .A2(W2496), .ZN(O935));
  NANDX1 G1737 (.A1(W362), .A2(W837), .ZN(O929));
  NANDX1 G1738 (.A1(W638), .A2(W469), .ZN(O944));
  NANDX1 G1739 (.A1(W1744), .A2(W2404), .ZN(O946));
  NANDX1 G1740 (.A1(W87), .A2(W430), .ZN(O924));
  NANDX1 G1741 (.A1(W1658), .A2(W934), .ZN(W3264));
  NANDX1 G1742 (.A1(W909), .A2(W562), .ZN(O923));
  NANDX1 G1743 (.A1(W984), .A2(W2821), .ZN(O922));
  NANDX1 G1744 (.A1(W2650), .A2(W698), .ZN(W3188));
  NANDX1 G1745 (.A1(W171), .A2(W222), .ZN(W3299));
  NANDX1 G1746 (.A1(W219), .A2(W1366), .ZN(O951));
  NANDX1 G1747 (.A1(I96), .A2(W200), .ZN(O919));
  NANDX1 G1748 (.A1(W3053), .A2(W1063), .ZN(O916));
  NANDX1 G1749 (.A1(W1684), .A2(W2677), .ZN(O914));
  NANDX1 G1750 (.A1(W2468), .A2(W727), .ZN(O954));
  NANDX1 G1751 (.A1(W3170), .A2(W1120), .ZN(O957));
  NANDX1 G1752 (.A1(W577), .A2(I60), .ZN(O912));
  NANDX1 G1753 (.A1(W1469), .A2(W2677), .ZN(O958));
  NANDX1 G1754 (.A1(W1688), .A2(W3085), .ZN(O909));
  NANDX1 G1755 (.A1(W3124), .A2(W534), .ZN(W3245));
  NANDX1 G1756 (.A1(W596), .A2(W2537), .ZN(O908));
  NANDX1 G1757 (.A1(W3052), .A2(W640), .ZN(O961));
  NANDX1 G1758 (.A1(W2469), .A2(I137), .ZN(W3117));
  NANDX1 G1759 (.A1(W422), .A2(W2829), .ZN(O1003));
  NANDX1 G1760 (.A1(W3129), .A2(W3239), .ZN(W3382));
  NANDX1 G1761 (.A1(W3263), .A2(W368), .ZN(O1006));
  NANDX1 G1762 (.A1(W812), .A2(W1262), .ZN(W3139));
  NANDX1 G1763 (.A1(W1119), .A2(W3081), .ZN(O830));
  NANDX1 G1764 (.A1(W137), .A2(W170), .ZN(O828));
  NANDX1 G1765 (.A1(W1658), .A2(W2871), .ZN(O825));
  NANDX1 G1766 (.A1(W971), .A2(W982), .ZN(O824));
  NANDX1 G1767 (.A1(W2787), .A2(W2906), .ZN(O1007));
  NANDX1 G1768 (.A1(W246), .A2(W2327), .ZN(O1008));
  NANDX1 G1769 (.A1(W449), .A2(W1503), .ZN(W3389));
  NANDX1 G1770 (.A1(W699), .A2(W1491), .ZN(O818));
  NANDX1 G1771 (.A1(W327), .A2(W598), .ZN(O1009));
  NANDX1 G1772 (.A1(W2022), .A2(W1133), .ZN(O1002));
  NANDX1 G1773 (.A1(W1800), .A2(W2639), .ZN(O815));
  NANDX1 G1774 (.A1(W645), .A2(W2143), .ZN(O814));
  NANDX1 G1775 (.A1(W317), .A2(W860), .ZN(O813));
  NANDX1 G1776 (.A1(W2818), .A2(W120), .ZN(O812));
  NANDX1 G1777 (.A1(W2290), .A2(W2206), .ZN(O811));
  NANDX1 G1778 (.A1(W2069), .A2(W3299), .ZN(O1015));
  NANDX1 G1779 (.A1(W1628), .A2(W837), .ZN(W3400));
  NANDX1 G1780 (.A1(W3), .A2(W2958), .ZN(O1017));
  NANDX1 G1781 (.A1(W2424), .A2(W2411), .ZN(O805));
  NANDX1 G1782 (.A1(W1781), .A2(W1534), .ZN(O1021));
  NANDX1 G1783 (.A1(W749), .A2(W1105), .ZN(O802));
  NANDX1 G1784 (.A1(W524), .A2(W344), .ZN(O801));
  NANDX1 G1785 (.A1(I7), .A2(W2498), .ZN(O1025));
  NANDX1 G1786 (.A1(W1623), .A2(W2293), .ZN(O851));
  NANDX1 G1787 (.A1(W51), .A2(W858), .ZN(W3187));
  NANDX1 G1788 (.A1(W2119), .A2(W264), .ZN(O867));
  NANDX1 G1789 (.A1(W580), .A2(W2054), .ZN(O990));
  NANDX1 G1790 (.A1(W1076), .A2(W1823), .ZN(O864));
  NANDX1 G1791 (.A1(W1584), .A2(W3022), .ZN(W3179));
  NANDX1 G1792 (.A1(W2628), .A2(W363), .ZN(O991));
  NANDX1 G1793 (.A1(W2311), .A2(W1236), .ZN(O860));
  NANDX1 G1794 (.A1(W2134), .A2(W78), .ZN(O858));
  NANDX1 G1795 (.A1(W1435), .A2(W1157), .ZN(O857));
  NANDX1 G1796 (.A1(W1066), .A2(W1980), .ZN(O856));
  NANDX1 G1797 (.A1(W2628), .A2(W2443), .ZN(W3367));
  NANDX1 G1798 (.A1(W236), .A2(W1515), .ZN(O854));
  NANDX1 G1799 (.A1(W2603), .A2(W2861), .ZN(O853));
  NANDX1 G1800 (.A1(W3472), .A2(W1567), .ZN(O1131));
  NANDX1 G1801 (.A1(W1377), .A2(W2020), .ZN(W3162));
  NANDX1 G1802 (.A1(W1357), .A2(W710), .ZN(O997));
  NANDX1 G1803 (.A1(W793), .A2(W3054), .ZN(O848));
  NANDX1 G1804 (.A1(W2394), .A2(W1779), .ZN(O846));
  NANDX1 G1805 (.A1(W2959), .A2(W721), .ZN(O999));
  NANDX1 G1806 (.A1(W2934), .A2(W121), .ZN(O841));
  NANDX1 G1807 (.A1(W2487), .A2(W363), .ZN(O840));
  NANDX1 G1808 (.A1(W2930), .A2(W1410), .ZN(O839));
  NANDX1 G1809 (.A1(W468), .A2(W2421), .ZN(O838));
  NANDX1 G1810 (.A1(W2764), .A2(W2525), .ZN(O836));
  NANDX1 G1811 (.A1(W1963), .A2(W693), .ZN(O1001));
  NANDX1 G1812 (.A1(I70), .A2(W1708), .ZN(O834));
  NANDX1 G1813 (.A1(W1714), .A2(W402), .ZN(W2599));
  NANDX1 G1814 (.A1(W186), .A2(W824), .ZN(O535));
  NANDX1 G1815 (.A1(W1168), .A2(W1376), .ZN(W2627));
  NANDX1 G1816 (.A1(W1341), .A2(W1305), .ZN(O534));
  NANDX1 G1817 (.A1(W1346), .A2(W128), .ZN(W2624));
  NANDX1 G1818 (.A1(W1748), .A2(W908), .ZN(W2620));
  NANDX1 G1819 (.A1(W1726), .A2(W2453), .ZN(O530));
  NANDX1 G1820 (.A1(W1363), .A2(W2510), .ZN(O529));
  NANDX1 G1821 (.A1(W75), .A2(W433), .ZN(W2615));
  NANDX1 G1822 (.A1(W1405), .A2(W1479), .ZN(O1278));
  NANDX1 G1823 (.A1(W164), .A2(W1232), .ZN(O523));
  NANDX1 G1824 (.A1(W2601), .A2(W565), .ZN(W2606));
  NANDX1 G1825 (.A1(W981), .A2(W2323), .ZN(O522));
  NANDX1 G1826 (.A1(W1792), .A2(W738), .ZN(O521));
  NANDX1 G1827 (.A1(W1345), .A2(W1960), .ZN(O537));
  NANDX1 G1828 (.A1(W1256), .A2(W1024), .ZN(O1287));
  NANDX1 G1829 (.A1(W179), .A2(W1062), .ZN(W2597));
  NANDX1 G1830 (.A1(W2116), .A2(W1741), .ZN(W2594));
  NANDX1 G1831 (.A1(W635), .A2(W838), .ZN(O517));
  NANDX1 G1832 (.A1(W1156), .A2(W60), .ZN(W2588));
  NANDX1 G1833 (.A1(W1127), .A2(W786), .ZN(O513));
  NANDX1 G1834 (.A1(W1027), .A2(W168), .ZN(O1292));
  NANDX1 G1835 (.A1(W2123), .A2(W1163), .ZN(W2581));
  NANDX1 G1836 (.A1(W1292), .A2(W3451), .ZN(O1293));
  NANDX1 G1837 (.A1(W997), .A2(W3034), .ZN(O1298));
  NANDX1 G1838 (.A1(W1857), .A2(W120), .ZN(W3750));
  NANDX1 G1839 (.A1(W2292), .A2(W31), .ZN(O1299));
  NANDX1 G1840 (.A1(W770), .A2(W2487), .ZN(W2575));
  NANDX1 G1841 (.A1(W2310), .A2(W2128), .ZN(O560));
  NANDX1 G1842 (.A1(W1117), .A2(W1625), .ZN(O578));
  NANDX1 G1843 (.A1(W2253), .A2(I10), .ZN(W2700));
  NANDX1 G1844 (.A1(W1497), .A2(W532), .ZN(O572));
  NANDX1 G1845 (.A1(W3323), .A2(W579), .ZN(O1255));
  NANDX1 G1846 (.A1(W2538), .A2(W1418), .ZN(O569));
  NANDX1 G1847 (.A1(W1773), .A2(W1017), .ZN(O568));
  NANDX1 G1848 (.A1(W2009), .A2(W1168), .ZN(W2686));
  NANDX1 G1849 (.A1(W2097), .A2(W821), .ZN(O567));
  NANDX1 G1850 (.A1(W2452), .A2(W485), .ZN(O566));
  NANDX1 G1851 (.A1(W795), .A2(W702), .ZN(O564));
  NANDX1 G1852 (.A1(W1027), .A2(W2179), .ZN(O1259));
  NANDX1 G1853 (.A1(W801), .A2(W2012), .ZN(O563));
  NANDX1 G1854 (.A1(W1216), .A2(W1589), .ZN(O562));
  NANDX1 G1855 (.A1(W684), .A2(W2518), .ZN(O508));
  NANDX1 G1856 (.A1(W582), .A2(W1775), .ZN(O553));
  NANDX1 G1857 (.A1(W213), .A2(W562), .ZN(W2662));
  NANDX1 G1858 (.A1(W993), .A2(W1126), .ZN(O551));
  NANDX1 G1859 (.A1(W330), .A2(W1239), .ZN(O1263));
  NANDX1 G1860 (.A1(W2027), .A2(W519), .ZN(O550));
  NANDX1 G1861 (.A1(W666), .A2(W1273), .ZN(O546));
  NANDX1 G1862 (.A1(W752), .A2(W2973), .ZN(O1267));
  NANDX1 G1863 (.A1(W1889), .A2(W1738), .ZN(O1268));
  NANDX1 G1864 (.A1(W1525), .A2(W1356), .ZN(W2637));
  NANDX1 G1865 (.A1(W759), .A2(W1925), .ZN(O1269));
  NANDX1 G1866 (.A1(W1067), .A2(W2462), .ZN(O1270));
  NANDX1 G1867 (.A1(W1938), .A2(W1631), .ZN(W2636));
  NANDX1 G1868 (.A1(W1742), .A2(W857), .ZN(O538));
  NANDX1 G1869 (.A1(W363), .A2(W943), .ZN(W2505));
  NANDX1 G1870 (.A1(W877), .A2(W649), .ZN(O482));
  NANDX1 G1871 (.A1(I154), .A2(W1982), .ZN(W2523));
  NANDX1 G1872 (.A1(W1271), .A2(W2429), .ZN(O480));
  NANDX1 G1873 (.A1(W1528), .A2(W2007), .ZN(W2519));
  NANDX1 G1874 (.A1(W2079), .A2(W1466), .ZN(W2518));
  NANDX1 G1875 (.A1(W1440), .A2(W1855), .ZN(W2516));
  NANDX1 G1876 (.A1(W2311), .A2(I122), .ZN(O1335));
  NANDX1 G1877 (.A1(W1017), .A2(W1676), .ZN(O477));
  NANDX1 G1878 (.A1(W1307), .A2(W1652), .ZN(O476));
  NANDX1 G1879 (.A1(I176), .A2(W1382), .ZN(O475));
  NANDX1 G1880 (.A1(W925), .A2(W646), .ZN(W2509));
  NANDX1 G1881 (.A1(W2240), .A2(W502), .ZN(W3793));
  NANDX1 G1882 (.A1(W3538), .A2(W1375), .ZN(O1338));
  NANDX1 G1883 (.A1(W1366), .A2(W1812), .ZN(W2525));
  NANDX1 G1884 (.A1(W2450), .A2(W691), .ZN(W2502));
  NANDX1 G1885 (.A1(W1613), .A2(W2100), .ZN(O471));
  NANDX1 G1886 (.A1(W670), .A2(W3357), .ZN(O1342));
  NANDX1 G1887 (.A1(W2252), .A2(W1695), .ZN(O1344));
  NANDX1 G1888 (.A1(W152), .A2(W2309), .ZN(O470));
  NANDX1 G1889 (.A1(W432), .A2(W157), .ZN(O1355));
  NANDX1 G1890 (.A1(W906), .A2(W1798), .ZN(W2489));
  NANDX1 G1891 (.A1(W1815), .A2(W1114), .ZN(W2487));
  NANDX1 G1892 (.A1(W1923), .A2(I112), .ZN(W2483));
  NANDX1 G1893 (.A1(W1603), .A2(W1483), .ZN(O1363));
  NANDX1 G1894 (.A1(W15), .A2(W542), .ZN(W2471));
  NANDX1 G1895 (.A1(W2958), .A2(W2850), .ZN(O1365));
  NANDX1 G1896 (.A1(W986), .A2(W346), .ZN(W2469));
  NANDX1 G1897 (.A1(W2465), .A2(W2186), .ZN(O493));
  NANDX1 G1898 (.A1(W323), .A2(W102), .ZN(O505));
  NANDX1 G1899 (.A1(W1718), .A2(W1164), .ZN(W2567));
  NANDX1 G1900 (.A1(W3661), .A2(W2753), .ZN(O1302));
  NANDX1 G1901 (.A1(W2231), .A2(W839), .ZN(W3755));
  NANDX1 G1902 (.A1(W395), .A2(W661), .ZN(O501));
  NANDX1 G1903 (.A1(I122), .A2(W1754), .ZN(O1308));
  NANDX1 G1904 (.A1(W3485), .A2(W1387), .ZN(O1309));
  NANDX1 G1905 (.A1(W773), .A2(W3537), .ZN(O1310));
  NANDX1 G1906 (.A1(W1495), .A2(W1619), .ZN(O499));
  NANDX1 G1907 (.A1(W96), .A2(W1298), .ZN(O1311));
  NANDX1 G1908 (.A1(W2106), .A2(W1148), .ZN(O1315));
  NANDX1 G1909 (.A1(W1468), .A2(W2245), .ZN(O497));
  NANDX1 G1910 (.A1(W1389), .A2(W497), .ZN(W2551));
  NANDX1 G1911 (.A1(W2779), .A2(W2082), .ZN(O1247));
  NANDX1 G1912 (.A1(W2017), .A2(W1305), .ZN(W2544));
  NANDX1 G1913 (.A1(W1488), .A2(W495), .ZN(W2542));
  NANDX1 G1914 (.A1(W3438), .A2(W1933), .ZN(W3774));
  NANDX1 G1915 (.A1(W2507), .A2(W1040), .ZN(W2537));
  NANDX1 G1916 (.A1(W688), .A2(W2697), .ZN(O1324));
  NANDX1 G1917 (.A1(W1135), .A2(W1230), .ZN(W2535));
  NANDX1 G1918 (.A1(W1087), .A2(W1375), .ZN(O1325));
  NANDX1 G1919 (.A1(W1331), .A2(W175), .ZN(O1328));
  NANDX1 G1920 (.A1(W2241), .A2(W2508), .ZN(W2531));
  NANDX1 G1921 (.A1(W764), .A2(W48), .ZN(O1330));
  NANDX1 G1922 (.A1(W416), .A2(W91), .ZN(O483));
  NANDX1 G1923 (.A1(W339), .A2(W2996), .ZN(O1331));
  NANDX1 G1924 (.A1(W2384), .A2(W233), .ZN(O1164));
  NANDX1 G1925 (.A1(W1585), .A2(W1478), .ZN(O666));
  NANDX1 G1926 (.A1(W1448), .A2(W1159), .ZN(O665));
  NANDX1 G1927 (.A1(W2988), .A2(W2480), .ZN(O1154));
  NANDX1 G1928 (.A1(W2580), .A2(W82), .ZN(O1155));
  NANDX1 G1929 (.A1(W2402), .A2(W2082), .ZN(O656));
  NANDX1 G1930 (.A1(W1359), .A2(W815), .ZN(W3579));
  NANDX1 G1931 (.A1(W441), .A2(W2258), .ZN(O652));
  NANDX1 G1932 (.A1(W682), .A2(W1688), .ZN(W3580));
  NANDX1 G1933 (.A1(W581), .A2(W962), .ZN(W3582));
  NANDX1 G1934 (.A1(W2123), .A2(W2420), .ZN(W2828));
  NANDX1 G1935 (.A1(W1103), .A2(W1267), .ZN(W2827));
  NANDX1 G1936 (.A1(W283), .A2(W1014), .ZN(W2825));
  NANDX1 G1937 (.A1(W3579), .A2(W281), .ZN(W3584));
  NANDX1 G1938 (.A1(W2673), .A2(W1925), .ZN(O1151));
  NANDX1 G1939 (.A1(W2650), .A2(W236), .ZN(W2822));
  NANDX1 G1940 (.A1(W2305), .A2(W964), .ZN(W2820));
  NANDX1 G1941 (.A1(W1272), .A2(W2335), .ZN(W2819));
  NANDX1 G1942 (.A1(I188), .A2(W1460), .ZN(W2818));
  NANDX1 G1943 (.A1(W2302), .A2(W505), .ZN(O649));
  NANDX1 G1944 (.A1(I185), .A2(W2287), .ZN(O644));
  NANDX1 G1945 (.A1(W1716), .A2(W469), .ZN(W2808));
  NANDX1 G1946 (.A1(W321), .A2(W1278), .ZN(O641));
  NANDX1 G1947 (.A1(W2939), .A2(W1227), .ZN(W3599));
  NANDX1 G1948 (.A1(W2519), .A2(W2577), .ZN(W2804));
  NANDX1 G1949 (.A1(W2084), .A2(W779), .ZN(O1173));
  NANDX1 G1950 (.A1(W2855), .A2(W3249), .ZN(O1175));
  NANDX1 G1951 (.A1(W2615), .A2(W1891), .ZN(O639));
  NANDX1 G1952 (.A1(W2600), .A2(W1470), .ZN(W2876));
  NANDX1 G1953 (.A1(W1318), .A2(W66), .ZN(W2897));
  NANDX1 G1954 (.A1(W2252), .A2(W2556), .ZN(O1132));
  NANDX1 G1955 (.A1(W553), .A2(W1773), .ZN(O690));
  NANDX1 G1956 (.A1(W1172), .A2(W1650), .ZN(O1135));
  NANDX1 G1957 (.A1(W2957), .A2(W1376), .ZN(O1136));
  NANDX1 G1958 (.A1(W1233), .A2(W2441), .ZN(W2891));
  NANDX1 G1959 (.A1(I65), .A2(W882), .ZN(O688));
  NANDX1 G1960 (.A1(W1598), .A2(W1360), .ZN(W2889));
  NANDX1 G1961 (.A1(W1852), .A2(W622), .ZN(W2887));
  NANDX1 G1962 (.A1(W468), .A2(W351), .ZN(O686));
  NANDX1 G1963 (.A1(W2167), .A2(W1979), .ZN(O1139));
  NANDX1 G1964 (.A1(W2952), .A2(W3120), .ZN(O1142));
  NANDX1 G1965 (.A1(W2489), .A2(W916), .ZN(O683));
  NANDX1 G1966 (.A1(W10), .A2(W1344), .ZN(O1179));
  NANDX1 G1967 (.A1(W960), .A2(W936), .ZN(O679));
  NANDX1 G1968 (.A1(W135), .A2(I46), .ZN(O678));
  NANDX1 G1969 (.A1(W2938), .A2(W2289), .ZN(W3562));
  NANDX1 G1970 (.A1(I193), .A2(W65), .ZN(O675));
  NANDX1 G1971 (.A1(W263), .A2(W509), .ZN(W2868));
  NANDX1 G1972 (.A1(W1037), .A2(W927), .ZN(W2867));
  NANDX1 G1973 (.A1(W2439), .A2(W112), .ZN(O673));
  NANDX1 G1974 (.A1(W2535), .A2(W2051), .ZN(W2864));
  NANDX1 G1975 (.A1(W1538), .A2(W1504), .ZN(O672));
  NANDX1 G1976 (.A1(W1030), .A2(W2433), .ZN(O671));
  NANDX1 G1977 (.A1(W2974), .A2(W944), .ZN(O1148));
  NANDX1 G1978 (.A1(W2385), .A2(W541), .ZN(W3568));
  NANDX1 G1979 (.A1(W175), .A2(W1192), .ZN(W2853));
  NANDX1 G1980 (.A1(W2443), .A2(W2398), .ZN(W2724));
  NANDX1 G1981 (.A1(W1458), .A2(W989), .ZN(O605));
  NANDX1 G1982 (.A1(W1117), .A2(I81), .ZN(O604));
  NANDX1 G1983 (.A1(W2119), .A2(W2857), .ZN(O1206));
  NANDX1 G1984 (.A1(W1059), .A2(W2117), .ZN(O599));
  NANDX1 G1985 (.A1(W2271), .A2(W1934), .ZN(O1216));
  NANDX1 G1986 (.A1(W982), .A2(W1734), .ZN(O598));
  NANDX1 G1987 (.A1(W46), .A2(I109), .ZN(W2736));
  NANDX1 G1988 (.A1(W1795), .A2(W870), .ZN(W2733));
  NANDX1 G1989 (.A1(W195), .A2(W1934), .ZN(O594));
  NANDX1 G1990 (.A1(W2462), .A2(I134), .ZN(O593));
  NANDX1 G1991 (.A1(W1121), .A2(W2722), .ZN(W2728));
  NANDX1 G1992 (.A1(W806), .A2(W1731), .ZN(O1222));
  NANDX1 G1993 (.A1(W733), .A2(W2120), .ZN(O590));
  NANDX1 G1994 (.A1(W2345), .A2(W2072), .ZN(O606));
  NANDX1 G1995 (.A1(W2594), .A2(W2545), .ZN(W2722));
  NANDX1 G1996 (.A1(W2339), .A2(W3365), .ZN(O1224));
  NANDX1 G1997 (.A1(I104), .A2(W67), .ZN(W2720));
  NANDX1 G1998 (.A1(W2926), .A2(W498), .ZN(W3668));
  NANDX1 G1999 (.A1(W154), .A2(W1348), .ZN(W2719));
  NANDX1 G2000 (.A1(I147), .A2(W1706), .ZN(O1232));
  NANDX1 G2001 (.A1(I22), .A2(W1378), .ZN(O1234));
  NANDX1 G2002 (.A1(W2069), .A2(W2939), .ZN(O1235));
  NANDX1 G2003 (.A1(W972), .A2(W2263), .ZN(W2708));
  NANDX1 G2004 (.A1(W494), .A2(W737), .ZN(O581));
  NANDX1 G2005 (.A1(W602), .A2(W3607), .ZN(O1239));
  NANDX1 G2006 (.A1(W465), .A2(W2238), .ZN(O1244));
  NANDX1 G2007 (.A1(W364), .A2(W3372), .ZN(O1245));
  NANDX1 G2008 (.A1(W1710), .A2(W2317), .ZN(O619));
  NANDX1 G2009 (.A1(W1815), .A2(W3590), .ZN(W3609));
  NANDX1 G2010 (.A1(W717), .A2(W818), .ZN(O636));
  NANDX1 G2011 (.A1(I20), .A2(W1469), .ZN(O630));
  NANDX1 G2012 (.A1(W2691), .A2(W203), .ZN(O629));
  NANDX1 G2013 (.A1(W1540), .A2(W2138), .ZN(O1182));
  NANDX1 G2014 (.A1(W1316), .A2(W1355), .ZN(O628));
  NANDX1 G2015 (.A1(W1364), .A2(W2196), .ZN(O627));
  NANDX1 G2016 (.A1(W157), .A2(W1770), .ZN(O1186));
  NANDX1 G2017 (.A1(W1462), .A2(W35), .ZN(O625));
  NANDX1 G2018 (.A1(W3323), .A2(W2825), .ZN(O1187));
  NANDX1 G2019 (.A1(W2974), .A2(W2730), .ZN(O1188));
  NANDX1 G2020 (.A1(W1433), .A2(W1341), .ZN(O621));
  NANDX1 G2021 (.A1(W1378), .A2(W892), .ZN(O620));
  NANDX1 G2022 (.A1(W2380), .A2(W935), .ZN(W2468));
  NANDX1 G2023 (.A1(W1696), .A2(W1006), .ZN(O618));
  NANDX1 G2024 (.A1(I111), .A2(W269), .ZN(O617));
  NANDX1 G2025 (.A1(W372), .A2(W632), .ZN(W2772));
  NANDX1 G2026 (.A1(W1053), .A2(W440), .ZN(O615));
  NANDX1 G2027 (.A1(W1325), .A2(W2268), .ZN(O1196));
  NANDX1 G2028 (.A1(W2984), .A2(W328), .ZN(O1198));
  NANDX1 G2029 (.A1(W2141), .A2(W1990), .ZN(W3633));
  NANDX1 G2030 (.A1(W1392), .A2(W415), .ZN(O613));
  NANDX1 G2031 (.A1(W1926), .A2(W509), .ZN(O1202));
  NANDX1 G2032 (.A1(W152), .A2(W1032), .ZN(W2754));
  NANDX1 G2033 (.A1(W80), .A2(W2110), .ZN(W2752));
  NANDX1 G2034 (.A1(W782), .A2(W2000), .ZN(O607));
  NANDX1 G2035 (.A1(W334), .A2(W114), .ZN(W474));
  NANDX1 G2036 (.A1(W343), .A2(W734), .ZN(W1335));
  NANDX1 G2037 (.A1(W59), .A2(I114), .ZN(W459));
  NANDX1 G2038 (.A1(W1128), .A2(I182), .ZN(O105));
  NANDX1 G2039 (.A1(I2), .A2(W191), .ZN(W462));
  NANDX1 G2040 (.A1(W0), .A2(W352), .ZN(W464));
  NANDX1 G2041 (.A1(W69), .A2(W97), .ZN(W469));
  NANDX1 G2042 (.A1(W142), .A2(W604), .ZN(W1320));
  NANDX1 G2043 (.A1(I138), .A2(W1258), .ZN(O103));
  NANDX1 G2044 (.A1(W961), .A2(W624), .ZN(O102));
  NANDX1 G2045 (.A1(W139), .A2(W108), .ZN(W470));
  NANDX1 G2046 (.A1(I81), .A2(I58), .ZN(W471));
  NANDX1 G2047 (.A1(W641), .A2(W289), .ZN(W1316));
  NANDX1 G2048 (.A1(W37), .A2(W1180), .ZN(W1315));
  NANDX1 G2049 (.A1(W1303), .A2(W1213), .ZN(W1338));
  NANDX1 G2050 (.A1(I26), .A2(W3), .ZN(W476));
  NANDX1 G2051 (.A1(W93), .A2(W71), .ZN(W1311));
  NANDX1 G2052 (.A1(W86), .A2(W164), .ZN(W477));
  NANDX1 G2053 (.A1(W472), .A2(W14), .ZN(W478));
  NANDX1 G2054 (.A1(I109), .A2(I185), .ZN(W479));
  NANDX1 G2055 (.A1(W1094), .A2(W763), .ZN(W1303));
  NANDX1 G2056 (.A1(I102), .A2(W1053), .ZN(W1301));
  NANDX1 G2057 (.A1(W981), .A2(I81), .ZN(W1300));
  NANDX1 G2058 (.A1(W1168), .A2(W1262), .ZN(W1297));
  NANDX1 G2059 (.A1(W527), .A2(I9), .ZN(O96));
  NANDX1 G2060 (.A1(W99), .A2(I24), .ZN(W485));
  NANDX1 G2061 (.A1(W333), .A2(W5), .ZN(W487));
  NANDX1 G2062 (.A1(W973), .A2(I56), .ZN(O94));
  NANDX1 G2063 (.A1(W333), .A2(W42), .ZN(W447));
  NANDX1 G2064 (.A1(W407), .A2(I168), .ZN(O10));
  NANDX1 G2065 (.A1(W1157), .A2(W941), .ZN(W1383));
  NANDX1 G2066 (.A1(W298), .A2(W1381), .ZN(W1382));
  NANDX1 G2067 (.A1(I65), .A2(W185), .ZN(W1381));
  NANDX1 G2068 (.A1(W328), .A2(I26), .ZN(W440));
  NANDX1 G2069 (.A1(I192), .A2(W271), .ZN(W1376));
  NANDX1 G2070 (.A1(I4), .A2(W842), .ZN(W1373));
  NANDX1 G2071 (.A1(W960), .A2(W144), .ZN(O110));
  NANDX1 G2072 (.A1(W575), .A2(W1335), .ZN(W1367));
  NANDX1 G2073 (.A1(W1292), .A2(W611), .ZN(W1366));
  NANDX1 G2074 (.A1(I184), .A2(W245), .ZN(W444));
  NANDX1 G2075 (.A1(W120), .A2(W221), .ZN(W445));
  NANDX1 G2076 (.A1(W124), .A2(I92), .ZN(W446));
  NANDX1 G2077 (.A1(W337), .A2(W142), .ZN(W488));
  NANDX1 G2078 (.A1(W1292), .A2(W1249), .ZN(W1360));
  NANDX1 G2079 (.A1(W160), .A2(W7), .ZN(W450));
  NANDX1 G2080 (.A1(W326), .A2(W666), .ZN(O108));
  NANDX1 G2081 (.A1(W1080), .A2(W1030), .ZN(W1355));
  NANDX1 G2082 (.A1(W54), .A2(W437), .ZN(W452));
  NANDX1 G2083 (.A1(W248), .A2(W28), .ZN(W455));
  NANDX1 G2084 (.A1(W1261), .A2(W503), .ZN(W1345));
  NANDX1 G2085 (.A1(I135), .A2(W107), .ZN(W1343));
  NANDX1 G2086 (.A1(W934), .A2(W1232), .ZN(O107));
  NANDX1 G2087 (.A1(I8), .A2(W386), .ZN(W1341));
  NANDX1 G2088 (.A1(W1232), .A2(W493), .ZN(W1340));
  NANDX1 G2089 (.A1(W367), .A2(W20), .ZN(W1339));
  NANDX1 G2090 (.A1(W45), .A2(W84), .ZN(W457));
  NANDX1 G2091 (.A1(W3), .A2(W514), .ZN(W1209));
  NANDX1 G2092 (.A1(W16), .A2(I138), .ZN(W525));
  NANDX1 G2093 (.A1(W1100), .A2(W666), .ZN(W1226));
  NANDX1 G2094 (.A1(W357), .A2(W139), .ZN(W526));
  NANDX1 G2095 (.A1(I62), .A2(W96), .ZN(W527));
  NANDX1 G2096 (.A1(W1150), .A2(W890), .ZN(W1223));
  NANDX1 G2097 (.A1(W149), .A2(I60), .ZN(W528));
  NANDX1 G2098 (.A1(W195), .A2(W403), .ZN(W535));
  NANDX1 G2099 (.A1(I76), .A2(W414), .ZN(W536));
  NANDX1 G2100 (.A1(I30), .A2(W191), .ZN(W1217));
  NANDX1 G2101 (.A1(W1042), .A2(W740), .ZN(W1216));
  NANDX1 G2102 (.A1(W512), .A2(W516), .ZN(O80));
  NANDX1 G2103 (.A1(W391), .A2(W39), .ZN(W543));
  NANDX1 G2104 (.A1(W459), .A2(I68), .ZN(W545));
  NANDX1 G2105 (.A1(W299), .A2(W463), .ZN(W524));
  NANDX1 G2106 (.A1(I158), .A2(W512), .ZN(W1208));
  NANDX1 G2107 (.A1(I21), .A2(W542), .ZN(O79));
  NANDX1 G2108 (.A1(W173), .A2(W479), .ZN(W1205));
  NANDX1 G2109 (.A1(I164), .A2(W785), .ZN(W1204));
  NANDX1 G2110 (.A1(W967), .A2(W1194), .ZN(W1203));
  NANDX1 G2111 (.A1(W161), .A2(W319), .ZN(W546));
  NANDX1 G2112 (.A1(W752), .A2(W320), .ZN(O78));
  NANDX1 G2113 (.A1(W1081), .A2(I54), .ZN(W1198));
  NANDX1 G2114 (.A1(W368), .A2(W1158), .ZN(W1196));
  NANDX1 G2115 (.A1(W462), .A2(W433), .ZN(W549));
  NANDX1 G2116 (.A1(W147), .A2(W509), .ZN(W551));
  NANDX1 G2117 (.A1(W240), .A2(W92), .ZN(W552));
  NANDX1 G2118 (.A1(I92), .A2(W201), .ZN(W553));
  NANDX1 G2119 (.A1(W1102), .A2(I153), .ZN(W1261));
  NANDX1 G2120 (.A1(W463), .A2(W325), .ZN(W489));
  NANDX1 G2121 (.A1(W1083), .A2(W487), .ZN(W1281));
  NANDX1 G2122 (.A1(W401), .A2(W448), .ZN(W1280));
  NANDX1 G2123 (.A1(W217), .A2(W51), .ZN(W494));
  NANDX1 G2124 (.A1(W31), .A2(I28), .ZN(W1278));
  NANDX1 G2125 (.A1(W921), .A2(W989), .ZN(W1277));
  NANDX1 G2126 (.A1(W118), .A2(W861), .ZN(W1276));
  NANDX1 G2127 (.A1(W670), .A2(W308), .ZN(W1274));
  NANDX1 G2128 (.A1(I92), .A2(I196), .ZN(W496));
  NANDX1 G2129 (.A1(W11), .A2(W1119), .ZN(O92));
  NANDX1 G2130 (.A1(W122), .A2(W466), .ZN(W1265));
  NANDX1 G2131 (.A1(W80), .A2(W239), .ZN(W497));
  NANDX1 G2132 (.A1(I19), .A2(W473), .ZN(W498));
  NANDX1 G2133 (.A1(W757), .A2(W387), .ZN(W1384));
  NANDX1 G2134 (.A1(W156), .A2(W694), .ZN(W1260));
  NANDX1 G2135 (.A1(I122), .A2(W1072), .ZN(W1258));
  NANDX1 G2136 (.A1(W169), .A2(W292), .ZN(W502));
  NANDX1 G2137 (.A1(I56), .A2(W872), .ZN(W1256));
  NANDX1 G2138 (.A1(W496), .A2(W199), .ZN(W508));
  NANDX1 G2139 (.A1(I172), .A2(W272), .ZN(W509));
  NANDX1 G2140 (.A1(W95), .A2(W101), .ZN(W512));
  NANDX1 G2141 (.A1(W309), .A2(W106), .ZN(W513));
  NANDX1 G2142 (.A1(I80), .A2(W1221), .ZN(W1239));
  NANDX1 G2143 (.A1(I86), .A2(W208), .ZN(W1235));
  NANDX1 G2144 (.A1(I165), .A2(I196), .ZN(W516));
  NANDX1 G2145 (.A1(W390), .A2(W1016), .ZN(W1233));
  NANDX1 G2146 (.A1(W1132), .A2(W1070), .ZN(W1232));
  NANDX1 G2147 (.A1(W646), .A2(W309), .ZN(W1508));
  NANDX1 G2148 (.A1(I68), .A2(W183), .ZN(W325));
  NANDX1 G2149 (.A1(I88), .A2(W12), .ZN(W327));
  NANDX1 G2150 (.A1(W789), .A2(W332), .ZN(W1526));
  NANDX1 G2151 (.A1(W98), .A2(I146), .ZN(W328));
  NANDX1 G2152 (.A1(W1179), .A2(W735), .ZN(O135));
  NANDX1 G2153 (.A1(W353), .A2(W1460), .ZN(W1520));
  NANDX1 G2154 (.A1(I116), .A2(W702), .ZN(W1518));
  NANDX1 G2155 (.A1(I19), .A2(W273), .ZN(W331));
  NANDX1 G2156 (.A1(W171), .A2(I190), .ZN(W336));
  NANDX1 G2157 (.A1(W291), .A2(W70), .ZN(W1515));
  NANDX1 G2158 (.A1(W456), .A2(W1318), .ZN(W1511));
  NANDX1 G2159 (.A1(W823), .A2(W756), .ZN(O134));
  NANDX1 G2160 (.A1(W641), .A2(W490), .ZN(O133));
  NANDX1 G2161 (.A1(I36), .A2(W382), .ZN(W1529));
  NANDX1 G2162 (.A1(W161), .A2(W67), .ZN(W341));
  NANDX1 G2163 (.A1(W171), .A2(W994), .ZN(W1502));
  NANDX1 G2164 (.A1(W758), .A2(W132), .ZN(O132));
  NANDX1 G2165 (.A1(W474), .A2(W1330), .ZN(W1494));
  NANDX1 G2166 (.A1(W143), .A2(W16), .ZN(W344));
  NANDX1 G2167 (.A1(W146), .A2(I96), .ZN(W347));
  NANDX1 G2168 (.A1(I198), .A2(W268), .ZN(W349));
  NANDX1 G2169 (.A1(W1391), .A2(I104), .ZN(O130));
  NANDX1 G2170 (.A1(W749), .A2(W3), .ZN(W1489));
  NANDX1 G2171 (.A1(W58), .A2(W12), .ZN(W351));
  NANDX1 G2172 (.A1(I195), .A2(I138), .ZN(W352));
  NANDX1 G2173 (.A1(W127), .A2(W287), .ZN(W354));
  NANDX1 G2174 (.A1(I32), .A2(I170), .ZN(W358));
  NANDX1 G2175 (.A1(W1), .A2(W409), .ZN(W1552));
  NANDX1 G2176 (.A1(W795), .A2(W938), .ZN(O149));
  NANDX1 G2177 (.A1(W136), .A2(I22), .ZN(W297));
  NANDX1 G2178 (.A1(W68), .A2(W1060), .ZN(W1579));
  NANDX1 G2179 (.A1(I144), .A2(W1099), .ZN(W1573));
  NANDX1 G2180 (.A1(W1530), .A2(W1491), .ZN(W1571));
  NANDX1 G2181 (.A1(I194), .A2(W1465), .ZN(W1570));
  NANDX1 G2182 (.A1(W196), .A2(W52), .ZN(W301));
  NANDX1 G2183 (.A1(I116), .A2(W728), .ZN(W1567));
  NANDX1 G2184 (.A1(W93), .A2(W1533), .ZN(O143));
  NANDX1 G2185 (.A1(W951), .A2(W89), .ZN(O141));
  NANDX1 G2186 (.A1(W306), .A2(W157), .ZN(W309));
  NANDX1 G2187 (.A1(W1448), .A2(W784), .ZN(O139));
  NANDX1 G2188 (.A1(W861), .A2(W1205), .ZN(W1553));
  NANDX1 G2189 (.A1(W117), .A2(I134), .ZN(W360));
  NANDX1 G2190 (.A1(W724), .A2(W461), .ZN(O138));
  NANDX1 G2191 (.A1(W22), .A2(I92), .ZN(W312));
  NANDX1 G2192 (.A1(W972), .A2(W1453), .ZN(O136));
  NANDX1 G2193 (.A1(W872), .A2(W1484), .ZN(W1544));
  NANDX1 G2194 (.A1(W652), .A2(W549), .ZN(W1543));
  NANDX1 G2195 (.A1(I95), .A2(W1516), .ZN(W1542));
  NANDX1 G2196 (.A1(W107), .A2(W1322), .ZN(W1539));
  NANDX1 G2197 (.A1(W1267), .A2(W185), .ZN(W1538));
  NANDX1 G2198 (.A1(W46), .A2(W92), .ZN(W317));
  NANDX1 G2199 (.A1(W1387), .A2(W1177), .ZN(W1535));
  NANDX1 G2200 (.A1(W96), .A2(W312), .ZN(W320));
  NANDX1 G2201 (.A1(W124), .A2(W26), .ZN(W321));
  NANDX1 G2202 (.A1(W266), .A2(I55), .ZN(W322));
  NANDX1 G2203 (.A1(W842), .A2(W751), .ZN(W1406));
  NANDX1 G2204 (.A1(W134), .A2(W317), .ZN(W412));
  NANDX1 G2205 (.A1(W1278), .A2(W261), .ZN(O118));
  NANDX1 G2206 (.A1(W754), .A2(W411), .ZN(W1422));
  NANDX1 G2207 (.A1(W79), .A2(W274), .ZN(W1419));
  NANDX1 G2208 (.A1(W227), .A2(W180), .ZN(W415));
  NANDX1 G2209 (.A1(W272), .A2(W36), .ZN(W416));
  NANDX1 G2210 (.A1(W1146), .A2(W1353), .ZN(W1418));
  NANDX1 G2211 (.A1(W245), .A2(W1079), .ZN(W1417));
  NANDX1 G2212 (.A1(W349), .A2(W766), .ZN(W1414));
  NANDX1 G2213 (.A1(W16), .A2(W273), .ZN(W418));
  NANDX1 G2214 (.A1(W28), .A2(I130), .ZN(W419));
  NANDX1 G2215 (.A1(W410), .A2(W294), .ZN(O9));
  NANDX1 G2216 (.A1(W836), .A2(W951), .ZN(W1408));
  NANDX1 G2217 (.A1(W257), .A2(W197), .ZN(W1424));
  NANDX1 G2218 (.A1(W1218), .A2(W801), .ZN(W1403));
  NANDX1 G2219 (.A1(W75), .A2(W226), .ZN(W426));
  NANDX1 G2220 (.A1(W1329), .A2(W80), .ZN(W1401));
  NANDX1 G2221 (.A1(W109), .A2(I146), .ZN(W427));
  NANDX1 G2222 (.A1(W1339), .A2(W1121), .ZN(O113));
  NANDX1 G2223 (.A1(W1279), .A2(I193), .ZN(W1397));
  NANDX1 G2224 (.A1(W931), .A2(W86), .ZN(W1396));
  NANDX1 G2225 (.A1(W487), .A2(W979), .ZN(W1395));
  NANDX1 G2226 (.A1(W902), .A2(W513), .ZN(W1394));
  NANDX1 G2227 (.A1(W227), .A2(I19), .ZN(W1392));
  NANDX1 G2228 (.A1(W192), .A2(W241), .ZN(W1391));
  NANDX1 G2229 (.A1(W726), .A2(W684), .ZN(W1390));
  NANDX1 G2230 (.A1(W456), .A2(W654), .ZN(W1388));
  NANDX1 G2231 (.A1(W883), .A2(W1329), .ZN(W1455));
  NANDX1 G2232 (.A1(W212), .A2(W136), .ZN(W361));
  NANDX1 G2233 (.A1(W1452), .A2(W795), .ZN(W1473));
  NANDX1 G2234 (.A1(I102), .A2(I175), .ZN(W362));
  NANDX1 G2235 (.A1(W816), .A2(W1076), .ZN(W1470));
  NANDX1 G2236 (.A1(W103), .A2(W328), .ZN(W368));
  NANDX1 G2237 (.A1(W345), .A2(W312), .ZN(W1468));
  NANDX1 G2238 (.A1(W1171), .A2(W225), .ZN(O126));
  NANDX1 G2239 (.A1(W566), .A2(I84), .ZN(W1461));
  NANDX1 G2240 (.A1(W1238), .A2(W367), .ZN(W1460));
  NANDX1 G2241 (.A1(W805), .A2(W163), .ZN(W1459));
  NANDX1 G2242 (.A1(I43), .A2(I85), .ZN(W373));
  NANDX1 G2243 (.A1(I185), .A2(W1101), .ZN(W1458));
  NANDX1 G2244 (.A1(W837), .A2(W300), .ZN(W1457));
  NANDX1 G2245 (.A1(I74), .A2(W381), .ZN(W1194));
  NANDX1 G2246 (.A1(W380), .A2(W1216), .ZN(W1454));
  NANDX1 G2247 (.A1(W77), .A2(I24), .ZN(W381));
  NANDX1 G2248 (.A1(W55), .A2(W211), .ZN(W387));
  NANDX1 G2249 (.A1(W307), .A2(I111), .ZN(W389));
  NANDX1 G2250 (.A1(W1), .A2(I13), .ZN(W391));
  NANDX1 G2251 (.A1(W1018), .A2(W195), .ZN(W1446));
  NANDX1 G2252 (.A1(I198), .A2(W316), .ZN(W392));
  NANDX1 G2253 (.A1(W1108), .A2(W1024), .ZN(W1441));
  NANDX1 G2254 (.A1(I198), .A2(W1112), .ZN(O121));
  NANDX1 G2255 (.A1(I196), .A2(W1040), .ZN(W1429));
  NANDX1 G2256 (.A1(W284), .A2(W29), .ZN(W404));
  NANDX1 G2257 (.A1(W117), .A2(W246), .ZN(W407));
  NANDX1 G2258 (.A1(W15), .A2(W747), .ZN(W931));
  NANDX1 G2259 (.A1(W444), .A2(W307), .ZN(W705));
  NANDX1 G2260 (.A1(I191), .A2(I61), .ZN(W706));
  NANDX1 G2261 (.A1(W455), .A2(W203), .ZN(W949));
  NANDX1 G2262 (.A1(W413), .A2(I24), .ZN(W708));
  NANDX1 G2263 (.A1(I178), .A2(W671), .ZN(O22));
  NANDX1 G2264 (.A1(W679), .A2(I40), .ZN(W941));
  NANDX1 G2265 (.A1(W20), .A2(W685), .ZN(W938));
  NANDX1 G2266 (.A1(W447), .A2(W656), .ZN(W936));
  NANDX1 G2267 (.A1(W255), .A2(I182), .ZN(W715));
  NANDX1 G2268 (.A1(W887), .A2(W358), .ZN(W934));
  NANDX1 G2269 (.A1(W737), .A2(W743), .ZN(W933));
  NANDX1 G2270 (.A1(W596), .A2(I68), .ZN(W716));
  NANDX1 G2271 (.A1(I134), .A2(W246), .ZN(W932));
  NANDX1 G2272 (.A1(W105), .A2(W151), .ZN(W953));
  NANDX1 G2273 (.A1(W77), .A2(W254), .ZN(W717));
  NANDX1 G2274 (.A1(I137), .A2(W221), .ZN(W930));
  NANDX1 G2275 (.A1(W471), .A2(W666), .ZN(W929));
  NANDX1 G2276 (.A1(W456), .A2(I151), .ZN(W722));
  NANDX1 G2277 (.A1(W139), .A2(W48), .ZN(W723));
  NANDX1 G2278 (.A1(W123), .A2(W656), .ZN(W727));
  NANDX1 G2279 (.A1(W896), .A2(W835), .ZN(W921));
  NANDX1 G2280 (.A1(W352), .A2(W573), .ZN(W920));
  NANDX1 G2281 (.A1(W333), .A2(W146), .ZN(W728));
  NANDX1 G2282 (.A1(W490), .A2(W74), .ZN(W916));
  NANDX1 G2283 (.A1(W362), .A2(W108), .ZN(W730));
  NANDX1 G2284 (.A1(I46), .A2(W224), .ZN(W912));
  NANDX1 G2285 (.A1(W255), .A2(W759), .ZN(W908));
  NANDX1 G2286 (.A1(W289), .A2(I154), .ZN(W683));
  NANDX1 G2287 (.A1(W205), .A2(W406), .ZN(W995));
  NANDX1 G2288 (.A1(W857), .A2(I11), .ZN(W993));
  NANDX1 G2289 (.A1(W11), .A2(W618), .ZN(W991));
  NANDX1 G2290 (.A1(W150), .A2(W332), .ZN(W673));
  NANDX1 G2291 (.A1(W402), .A2(W34), .ZN(W675));
  NANDX1 G2292 (.A1(I142), .A2(W416), .ZN(W987));
  NANDX1 G2293 (.A1(W313), .A2(W67), .ZN(W985));
  NANDX1 G2294 (.A1(W155), .A2(W293), .ZN(W677));
  NANDX1 G2295 (.A1(W603), .A2(W535), .ZN(W679));
  NANDX1 G2296 (.A1(W782), .A2(W531), .ZN(W981));
  NANDX1 G2297 (.A1(I44), .A2(W31), .ZN(W682));
  NANDX1 G2298 (.A1(W24), .A2(W176), .ZN(W978));
  NANDX1 G2299 (.A1(W363), .A2(W703), .ZN(W977));
  NANDX1 G2300 (.A1(W282), .A2(W448), .ZN(W734));
  NANDX1 G2301 (.A1(W480), .A2(W300), .ZN(W974));
  NANDX1 G2302 (.A1(W131), .A2(W272), .ZN(W685));
  NANDX1 G2303 (.A1(W30), .A2(W562), .ZN(W686));
  NANDX1 G2304 (.A1(W145), .A2(W48), .ZN(W689));
  NANDX1 G2305 (.A1(W112), .A2(I10), .ZN(W690));
  NANDX1 G2306 (.A1(W131), .A2(W650), .ZN(W965));
  NANDX1 G2307 (.A1(W779), .A2(W760), .ZN(W964));
  NANDX1 G2308 (.A1(I58), .A2(W90), .ZN(W695));
  NANDX1 G2309 (.A1(W955), .A2(W886), .ZN(W961));
  NANDX1 G2310 (.A1(W238), .A2(W626), .ZN(W697));
  NANDX1 G2311 (.A1(I34), .A2(W474), .ZN(W699));
  NANDX1 G2312 (.A1(W79), .A2(W619), .ZN(W703));
  NANDX1 G2313 (.A1(W266), .A2(I136), .ZN(W954));
  NANDX1 G2314 (.A1(W409), .A2(W292), .ZN(W784));
  NANDX1 G2315 (.A1(W572), .A2(W552), .ZN(W765));
  NANDX1 G2316 (.A1(W80), .A2(W402), .ZN(W850));
  NANDX1 G2317 (.A1(W751), .A2(I76), .ZN(W766));
  NANDX1 G2318 (.A1(W565), .A2(W707), .ZN(O34));
  NANDX1 G2319 (.A1(W595), .A2(I6), .ZN(W847));
  NANDX1 G2320 (.A1(W712), .A2(W224), .ZN(O27));
  NANDX1 G2321 (.A1(W261), .A2(W109), .ZN(W846));
  NANDX1 G2322 (.A1(W490), .A2(I195), .ZN(W776));
  NANDX1 G2323 (.A1(W87), .A2(W587), .ZN(W835));
  NANDX1 G2324 (.A1(I174), .A2(W621), .ZN(W834));
  NANDX1 G2325 (.A1(I150), .A2(W282), .ZN(W778));
  NANDX1 G2326 (.A1(W291), .A2(W280), .ZN(W828));
  NANDX1 G2327 (.A1(W487), .A2(W663), .ZN(W826));
  NANDX1 G2328 (.A1(I50), .A2(W539), .ZN(W854));
  NANDX1 G2329 (.A1(W259), .A2(W807), .ZN(W823));
  NANDX1 G2330 (.A1(W86), .A2(W634), .ZN(W787));
  NANDX1 G2331 (.A1(W361), .A2(W629), .ZN(W815));
  NANDX1 G2332 (.A1(W418), .A2(W476), .ZN(W794));
  NANDX1 G2333 (.A1(I195), .A2(W487), .ZN(W795));
  NANDX1 G2334 (.A1(I36), .A2(W333), .ZN(W797));
  NANDX1 G2335 (.A1(W778), .A2(W110), .ZN(O30));
  NANDX1 G2336 (.A1(W50), .A2(W128), .ZN(W799));
  NANDX1 G2337 (.A1(W93), .A2(W15), .ZN(W810));
  NANDX1 G2338 (.A1(W438), .A2(W113), .ZN(W807));
  NANDX1 G2339 (.A1(W588), .A2(W436), .ZN(W806));
  NANDX1 G2340 (.A1(W741), .A2(W328), .ZN(W804));
  NANDX1 G2341 (.A1(I110), .A2(W201), .ZN(W800));
  NANDX1 G2342 (.A1(W706), .A2(W344), .ZN(O25));
  NANDX1 G2343 (.A1(I164), .A2(W92), .ZN(W907));
  NANDX1 G2344 (.A1(I142), .A2(I170), .ZN(W739));
  NANDX1 G2345 (.A1(W401), .A2(W208), .ZN(W902));
  NANDX1 G2346 (.A1(W193), .A2(I39), .ZN(W900));
  NANDX1 G2347 (.A1(W320), .A2(I45), .ZN(O40));
  NANDX1 G2348 (.A1(W794), .A2(W320), .ZN(W897));
  NANDX1 G2349 (.A1(W726), .A2(W162), .ZN(W894));
  NANDX1 G2350 (.A1(I43), .A2(W38), .ZN(W891));
  NANDX1 G2351 (.A1(W688), .A2(W44), .ZN(W741));
  NANDX1 G2352 (.A1(W15), .A2(W582), .ZN(W890));
  NANDX1 G2353 (.A1(W218), .A2(W737), .ZN(W742));
  NANDX1 G2354 (.A1(I156), .A2(I46), .ZN(W889));
  NANDX1 G2355 (.A1(W236), .A2(I75), .ZN(O39));
  NANDX1 G2356 (.A1(W599), .A2(W286), .ZN(O17));
  NANDX1 G2357 (.A1(W758), .A2(I147), .ZN(W885));
  NANDX1 G2358 (.A1(W359), .A2(I106), .ZN(W749));
  NANDX1 G2359 (.A1(W523), .A2(W465), .ZN(W751));
  NANDX1 G2360 (.A1(W617), .A2(W623), .ZN(W883));
  NANDX1 G2361 (.A1(W756), .A2(I176), .ZN(W879));
  NANDX1 G2362 (.A1(W259), .A2(W39), .ZN(O37));
  NANDX1 G2363 (.A1(W616), .A2(W692), .ZN(W755));
  NANDX1 G2364 (.A1(W482), .A2(I196), .ZN(W872));
  NANDX1 G2365 (.A1(W231), .A2(W32), .ZN(W871));
  NANDX1 G2366 (.A1(W683), .A2(W199), .ZN(W758));
  NANDX1 G2367 (.A1(W809), .A2(W786), .ZN(W866));
  NANDX1 G2368 (.A1(W242), .A2(W574), .ZN(W860));
  NANDX1 G2369 (.A1(W522), .A2(I145), .ZN(W764));
  NANDX1 G2370 (.A1(I111), .A2(W835), .ZN(W1111));
  NANDX1 G2371 (.A1(I40), .A2(W68), .ZN(W573));
  NANDX1 G2372 (.A1(W358), .A2(W414), .ZN(W574));
  NANDX1 G2373 (.A1(W433), .A2(W136), .ZN(W1135));
  NANDX1 G2374 (.A1(W339), .A2(W534), .ZN(W577));
  NANDX1 G2375 (.A1(W370), .A2(W541), .ZN(W1132));
  NANDX1 G2376 (.A1(W233), .A2(W467), .ZN(W1128));
  NANDX1 G2377 (.A1(W539), .A2(W553), .ZN(W581));
  NANDX1 G2378 (.A1(I146), .A2(W21), .ZN(W1126));
  NANDX1 G2379 (.A1(W910), .A2(W512), .ZN(O64));
  NANDX1 G2380 (.A1(W521), .A2(W124), .ZN(W582));
  NANDX1 G2381 (.A1(W1034), .A2(W108), .ZN(W1120));
  NANDX1 G2382 (.A1(W454), .A2(W320), .ZN(W587));
  NANDX1 G2383 (.A1(W613), .A2(W535), .ZN(W1113));
  NANDX1 G2384 (.A1(W1103), .A2(W976), .ZN(O67));
  NANDX1 G2385 (.A1(W561), .A2(W704), .ZN(W1110));
  NANDX1 G2386 (.A1(W95), .A2(W1020), .ZN(W1109));
  NANDX1 G2387 (.A1(W64), .A2(W108), .ZN(O63));
  NANDX1 G2388 (.A1(W415), .A2(I126), .ZN(W588));
  NANDX1 G2389 (.A1(W508), .A2(W1098), .ZN(W1103));
  NANDX1 G2390 (.A1(W510), .A2(W124), .ZN(W592));
  NANDX1 G2391 (.A1(W422), .A2(W720), .ZN(W1095));
  NANDX1 G2392 (.A1(W404), .A2(W1062), .ZN(W1093));
  NANDX1 G2393 (.A1(W486), .A2(W52), .ZN(W595));
  NANDX1 G2394 (.A1(W1090), .A2(W853), .ZN(W1091));
  NANDX1 G2395 (.A1(W908), .A2(W311), .ZN(W1090));
  NANDX1 G2396 (.A1(W683), .A2(W705), .ZN(O62));
  NANDX1 G2397 (.A1(W587), .A2(W247), .ZN(W1087));
  NANDX1 G2398 (.A1(W1134), .A2(I140), .ZN(O70));
  NANDX1 G2399 (.A1(W106), .A2(W80), .ZN(W555));
  NANDX1 G2400 (.A1(W358), .A2(I109), .ZN(W1190));
  NANDX1 G2401 (.A1(W2), .A2(W365), .ZN(O75));
  NANDX1 G2402 (.A1(W712), .A2(W1121), .ZN(O74));
  NANDX1 G2403 (.A1(W216), .A2(W349), .ZN(W557));
  NANDX1 G2404 (.A1(W149), .A2(W840), .ZN(O73));
  NANDX1 G2405 (.A1(I138), .A2(W336), .ZN(W1186));
  NANDX1 G2406 (.A1(W781), .A2(W1168), .ZN(O72));
  NANDX1 G2407 (.A1(W277), .A2(I13), .ZN(W559));
  NANDX1 G2408 (.A1(W232), .A2(W949), .ZN(W1179));
  NANDX1 G2409 (.A1(W490), .A2(I130), .ZN(O12));
  NANDX1 G2410 (.A1(I32), .A2(W507), .ZN(W561));
  NANDX1 G2411 (.A1(W69), .A2(W308), .ZN(W562));
  NANDX1 G2412 (.A1(W310), .A2(W143), .ZN(W605));
  NANDX1 G2413 (.A1(I36), .A2(W517), .ZN(W1168));
  NANDX1 G2414 (.A1(W41), .A2(W36), .ZN(W1164));
  NANDX1 G2415 (.A1(I56), .A2(I38), .ZN(W564));
  NANDX1 G2416 (.A1(W1057), .A2(W913), .ZN(W1158));
  NANDX1 G2417 (.A1(W318), .A2(W472), .ZN(W565));
  NANDX1 G2418 (.A1(I57), .A2(W550), .ZN(W1156));
  NANDX1 G2419 (.A1(W310), .A2(W927), .ZN(W1154));
  NANDX1 G2420 (.A1(W902), .A2(W863), .ZN(O68));
  NANDX1 G2421 (.A1(W757), .A2(W727), .ZN(W1150));
  NANDX1 G2422 (.A1(W351), .A2(W127), .ZN(W1148));
  NANDX1 G2423 (.A1(W1105), .A2(W336), .ZN(W1146));
  NANDX1 G2424 (.A1(W199), .A2(W127), .ZN(W1145));
  NANDX1 G2425 (.A1(W972), .A2(W309), .ZN(W1141));
  NANDX1 G2426 (.A1(W362), .A2(W182), .ZN(W656));
  NANDX1 G2427 (.A1(W464), .A2(I161), .ZN(W633));
  NANDX1 G2428 (.A1(W746), .A2(W153), .ZN(W1043));
  NANDX1 G2429 (.A1(W625), .A2(W561), .ZN(W636));
  NANDX1 G2430 (.A1(W533), .A2(W397), .ZN(W640));
  NANDX1 G2431 (.A1(W394), .A2(W276), .ZN(W1030));
  NANDX1 G2432 (.A1(W263), .A2(W381), .ZN(W644));
  NANDX1 G2433 (.A1(W114), .A2(W93), .ZN(W1028));
  NANDX1 G2434 (.A1(W1017), .A2(I147), .ZN(W1027));
  NANDX1 G2435 (.A1(W86), .A2(I148), .ZN(W1026));
  NANDX1 G2436 (.A1(W597), .A2(I170), .ZN(W645));
  NANDX1 G2437 (.A1(W318), .A2(W628), .ZN(W647));
  NANDX1 G2438 (.A1(W31), .A2(W216), .ZN(W648));
  NANDX1 G2439 (.A1(W0), .A2(W857), .ZN(W1020));
  NANDX1 G2440 (.A1(W9), .A2(W348), .ZN(W632));
  NANDX1 G2441 (.A1(I91), .A2(W379), .ZN(W1015));
  NANDX1 G2442 (.A1(I50), .A2(I90), .ZN(W657));
  NANDX1 G2443 (.A1(W741), .A2(I128), .ZN(O53));
  NANDX1 G2444 (.A1(I190), .A2(W609), .ZN(W1010));
  NANDX1 G2445 (.A1(W124), .A2(W887), .ZN(W1009));
  NANDX1 G2446 (.A1(I170), .A2(I79), .ZN(W661));
  NANDX1 G2447 (.A1(W188), .A2(W136), .ZN(W663));
  NANDX1 G2448 (.A1(W573), .A2(I6), .ZN(W667));
  NANDX1 G2449 (.A1(W273), .A2(W846), .ZN(W1005));
  NANDX1 G2450 (.A1(W367), .A2(W497), .ZN(W1001));
  NANDX1 G2451 (.A1(I66), .A2(W38), .ZN(W999));
  NANDX1 G2452 (.A1(W915), .A2(W172), .ZN(W997));
  NANDX1 G2453 (.A1(W238), .A2(W315), .ZN(W996));
  NANDX1 G2454 (.A1(W497), .A2(W189), .ZN(W615));
  NANDX1 G2455 (.A1(W639), .A2(W210), .ZN(W1086));
  NANDX1 G2456 (.A1(W537), .A2(W38), .ZN(W606));
  NANDX1 G2457 (.A1(W431), .A2(W268), .ZN(W1084));
  NANDX1 G2458 (.A1(I108), .A2(W518), .ZN(W607));
  NANDX1 G2459 (.A1(W296), .A2(W75), .ZN(O61));
  NANDX1 G2460 (.A1(W209), .A2(W637), .ZN(W1081));
  NANDX1 G2461 (.A1(W211), .A2(W531), .ZN(W1080));
  NANDX1 G2462 (.A1(W298), .A2(W1037), .ZN(W1079));
  NANDX1 G2463 (.A1(W499), .A2(W457), .ZN(W610));
  NANDX1 G2464 (.A1(W459), .A2(W955), .ZN(W1077));
  NANDX1 G2465 (.A1(I50), .A2(W782), .ZN(W1076));
  NANDX1 G2466 (.A1(W291), .A2(W533), .ZN(W613));
  NANDX1 G2467 (.A1(W349), .A2(W96), .ZN(W614));
  NANDX1 G2468 (.A1(W604), .A2(W982), .ZN(W2032));
  NANDX1 G2469 (.A1(W543), .A2(W835), .ZN(W1074));
  NANDX1 G2470 (.A1(W1047), .A2(W899), .ZN(W1073));
  NANDX1 G2471 (.A1(W95), .A2(W284), .ZN(W624));
  NANDX1 G2472 (.A1(W839), .A2(W22), .ZN(W1064));
  NANDX1 G2473 (.A1(W927), .A2(W695), .ZN(W1060));
  NANDX1 G2474 (.A1(W360), .A2(W263), .ZN(W1059));
  NANDX1 G2475 (.A1(W252), .A2(W655), .ZN(W1056));
  NANDX1 G2476 (.A1(W191), .A2(W609), .ZN(W1055));
  NANDX1 G2477 (.A1(W909), .A2(W1024), .ZN(W1054));
  NANDX1 G2478 (.A1(W618), .A2(W360), .ZN(W631));
  NANDX1 G2479 (.A1(W725), .A2(W78), .ZN(W1050));
  NANDX1 G2480 (.A1(W257), .A2(W202), .ZN(W1048));
  NANDX1 G2481 (.A1(W1306), .A2(W1629), .ZN(W1773));
  NANDX1 G2482 (.A1(I17), .A2(I91), .ZN(W1801));
  NANDX1 G2483 (.A1(W104), .A2(W1238), .ZN(W1796));
  NANDX1 G2484 (.A1(W41), .A2(I78), .ZN(W139));
  NANDX1 G2485 (.A1(W881), .A2(W633), .ZN(W1794));
  NANDX1 G2486 (.A1(W605), .A2(W1236), .ZN(O208));
  NANDX1 G2487 (.A1(W1470), .A2(W1344), .ZN(O207));
  NANDX1 G2488 (.A1(W20), .A2(W94), .ZN(W146));
  NANDX1 G2489 (.A1(W24), .A2(W71), .ZN(W148));
  NANDX1 G2490 (.A1(I186), .A2(W59), .ZN(W150));
  NANDX1 G2491 (.A1(I65), .A2(W1320), .ZN(W1777));
  NANDX1 G2492 (.A1(W7), .A2(I115), .ZN(W151));
  NANDX1 G2493 (.A1(I116), .A2(I156), .ZN(W1802));
  NANDX1 G2494 (.A1(W1490), .A2(W1586), .ZN(W1771));
  NANDX1 G2495 (.A1(W549), .A2(W1043), .ZN(W1769));
  NANDX1 G2496 (.A1(W758), .A2(W407), .ZN(O204));
  NANDX1 G2497 (.A1(W28), .A2(W49), .ZN(W155));
  NANDX1 G2498 (.A1(I175), .A2(I48), .ZN(W162));
  NANDX1 G2499 (.A1(W60), .A2(W111), .ZN(W163));
  NANDX1 G2500 (.A1(W511), .A2(W21), .ZN(O203));
  NANDX1 G2501 (.A1(W1300), .A2(I2), .ZN(O201));
  NANDX1 G2502 (.A1(W150), .A2(I86), .ZN(W164));
  NANDX1 G2503 (.A1(W806), .A2(W931), .ZN(W1762));
  NANDX1 G2504 (.A1(W251), .A2(W632), .ZN(W1758));
  NANDX1 G2505 (.A1(W1130), .A2(W1788), .ZN(W1821));
  NANDX1 G2506 (.A1(W1204), .A2(W627), .ZN(W1846));
  NANDX1 G2507 (.A1(W126), .A2(W1487), .ZN(W1845));
  NANDX1 G2508 (.A1(W56), .A2(I29), .ZN(W111));
  NANDX1 G2509 (.A1(W1714), .A2(W364), .ZN(W1837));
  NANDX1 G2510 (.A1(W1783), .A2(W541), .ZN(W1831));
  NANDX1 G2511 (.A1(I22), .A2(W1770), .ZN(W1830));
  NANDX1 G2512 (.A1(W106), .A2(I72), .ZN(W116));
  NANDX1 G2513 (.A1(I44), .A2(W88), .ZN(W117));
  NANDX1 G2514 (.A1(I100), .A2(I79), .ZN(W120));
  NANDX1 G2515 (.A1(W79), .A2(I134), .ZN(W121));
  NANDX1 G2516 (.A1(W1407), .A2(W708), .ZN(W1822));
  NANDX1 G2517 (.A1(W1045), .A2(W765), .ZN(W1756));
  NANDX1 G2518 (.A1(I52), .A2(I96), .ZN(W125));
  NANDX1 G2519 (.A1(W692), .A2(W520), .ZN(W1818));
  NANDX1 G2520 (.A1(W862), .A2(W1321), .ZN(W1815));
  NANDX1 G2521 (.A1(W1543), .A2(W1371), .ZN(O215));
  NANDX1 G2522 (.A1(W0), .A2(I39), .ZN(W128));
  NANDX1 G2523 (.A1(W1616), .A2(W1614), .ZN(O214));
  NANDX1 G2524 (.A1(W1766), .A2(W112), .ZN(W1809));
  NANDX1 G2525 (.A1(W1223), .A2(W129), .ZN(W1806));
  NANDX1 G2526 (.A1(W103), .A2(W7), .ZN(W131));
  NANDX1 G2527 (.A1(W54), .A2(W492), .ZN(W1803));
  NANDX1 G2528 (.A1(W127), .A2(W120), .ZN(W204));
  NANDX1 G2529 (.A1(W177), .A2(I31), .ZN(W199));
  NANDX1 G2530 (.A1(W861), .A2(W1408), .ZN(W1708));
  NANDX1 G2531 (.A1(W1610), .A2(W1253), .ZN(W1707));
  NANDX1 G2532 (.A1(W419), .A2(W657), .ZN(W1703));
  NANDX1 G2533 (.A1(W1048), .A2(W657), .ZN(O185));
  NANDX1 G2534 (.A1(I48), .A2(W47), .ZN(W203));
  NANDX1 G2535 (.A1(W1405), .A2(W229), .ZN(W1696));
  NANDX1 G2536 (.A1(W289), .A2(W875), .ZN(W1694));
  NANDX1 G2537 (.A1(I61), .A2(W324), .ZN(W1693));
  NANDX1 G2538 (.A1(W1006), .A2(W1403), .ZN(W1690));
  NANDX1 G2539 (.A1(I114), .A2(W1130), .ZN(O183));
  NANDX1 G2540 (.A1(W300), .A2(W1452), .ZN(W1710));
  NANDX1 G2541 (.A1(W203), .A2(W45), .ZN(O2));
  NANDX1 G2542 (.A1(W170), .A2(I126), .ZN(W215));
  NANDX1 G2543 (.A1(W46), .A2(W204), .ZN(W217));
  NANDX1 G2544 (.A1(W197), .A2(W1137), .ZN(O182));
  NANDX1 G2545 (.A1(W1481), .A2(W388), .ZN(O181));
  NANDX1 G2546 (.A1(I118), .A2(W182), .ZN(W223));
  NANDX1 G2547 (.A1(W195), .A2(W123), .ZN(W224));
  NANDX1 G2548 (.A1(W196), .A2(I61), .ZN(W225));
  NANDX1 G2549 (.A1(W336), .A2(W1441), .ZN(W1680));
  NANDX1 G2550 (.A1(W52), .A2(I114), .ZN(W227));
  NANDX1 G2551 (.A1(I88), .A2(W1408), .ZN(W1731));
  NANDX1 G2552 (.A1(W509), .A2(W1527), .ZN(W1754));
  NANDX1 G2553 (.A1(W119), .A2(I134), .ZN(W167));
  NANDX1 G2554 (.A1(W1385), .A2(W1406), .ZN(O198));
  NANDX1 G2555 (.A1(W1278), .A2(W963), .ZN(W1748));
  NANDX1 G2556 (.A1(W1447), .A2(W674), .ZN(W1747));
  NANDX1 G2557 (.A1(W256), .A2(W1629), .ZN(W1744));
  NANDX1 G2558 (.A1(W206), .A2(W1054), .ZN(O196));
  NANDX1 G2559 (.A1(I39), .A2(W991), .ZN(W1739));
  NANDX1 G2560 (.A1(I180), .A2(W144), .ZN(W170));
  NANDX1 G2561 (.A1(W364), .A2(W485), .ZN(W1737));
  NANDX1 G2562 (.A1(W61), .A2(W1190), .ZN(W1732));
  NANDX1 G2563 (.A1(W922), .A2(W1282), .ZN(O227));
  NANDX1 G2564 (.A1(W1007), .A2(W145), .ZN(W1729));
  NANDX1 G2565 (.A1(W1534), .A2(W32), .ZN(W1728));
  NANDX1 G2566 (.A1(I65), .A2(I82), .ZN(W177));
  NANDX1 G2567 (.A1(W932), .A2(W833), .ZN(W1725));
  NANDX1 G2568 (.A1(I120), .A2(W139), .ZN(W186));
  NANDX1 G2569 (.A1(I186), .A2(W2), .ZN(W190));
  NANDX1 G2570 (.A1(W660), .A2(W272), .ZN(O192));
  NANDX1 G2571 (.A1(W100), .A2(W51), .ZN(W192));
  NANDX1 G2572 (.A1(W104), .A2(W11), .ZN(W195));
  NANDX1 G2573 (.A1(W1080), .A2(W1232), .ZN(O189));
  NANDX1 G2574 (.A1(I84), .A2(I85), .ZN(W42));
  NANDX1 G2575 (.A1(W363), .A2(W825), .ZN(W1988));
  NANDX1 G2576 (.A1(W1702), .A2(W1483), .ZN(W1987));
  NANDX1 G2577 (.A1(I38), .A2(I39), .ZN(W19));
  NANDX1 G2578 (.A1(I44), .A2(I45), .ZN(W22));
  NANDX1 G2579 (.A1(W1260), .A2(W994), .ZN(W1985));
  NANDX1 G2580 (.A1(I54), .A2(I55), .ZN(W27));
  NANDX1 G2581 (.A1(I60), .A2(I61), .ZN(W30));
  NANDX1 G2582 (.A1(W1638), .A2(W1027), .ZN(O266));
  NANDX1 G2583 (.A1(W771), .A2(W982), .ZN(W1974));
  NANDX1 G2584 (.A1(W1824), .A2(W330), .ZN(O264));
  NANDX1 G2585 (.A1(W335), .A2(W1137), .ZN(W1969));
  NANDX1 G2586 (.A1(W1286), .A2(W1982), .ZN(W1990));
  NANDX1 G2587 (.A1(W218), .A2(W797), .ZN(W1963));
  NANDX1 G2588 (.A1(W766), .A2(W1023), .ZN(O261));
  NANDX1 G2589 (.A1(I94), .A2(I95), .ZN(W47));
  NANDX1 G2590 (.A1(W1629), .A2(W775), .ZN(W1954));
  NANDX1 G2591 (.A1(W161), .A2(W895), .ZN(W1953));
  NANDX1 G2592 (.A1(W1354), .A2(W1367), .ZN(W1952));
  NANDX1 G2593 (.A1(W257), .A2(W1352), .ZN(W1949));
  NANDX1 G2594 (.A1(I102), .A2(I103), .ZN(W51));
  NANDX1 G2595 (.A1(W1497), .A2(W1321), .ZN(O257));
  NANDX1 G2596 (.A1(W928), .A2(I13), .ZN(O256));
  NANDX1 G2597 (.A1(W1805), .A2(W1369), .ZN(W1940));
  NANDX1 G2598 (.A1(W988), .A2(W587), .ZN(W2011));
  NANDX1 G2599 (.A1(I2), .A2(I3), .ZN(W1));
  NANDX1 G2600 (.A1(I4), .A2(I5), .ZN(W2));
  NANDX1 G2601 (.A1(I12), .A2(I13), .ZN(W6));
  NANDX1 G2602 (.A1(I161), .A2(W548), .ZN(W2028));
  NANDX1 G2603 (.A1(I16), .A2(I17), .ZN(W8));
  NANDX1 G2604 (.A1(W2), .A2(W1606), .ZN(O277));
  NANDX1 G2605 (.A1(W135), .A2(W4), .ZN(W2020));
  NANDX1 G2606 (.A1(W382), .A2(W1218), .ZN(W2019));
  NANDX1 G2607 (.A1(I18), .A2(I19), .ZN(W9));
  NANDX1 G2608 (.A1(W1349), .A2(W826), .ZN(W2012));
  NANDX1 G2609 (.A1(I22), .A2(I23), .ZN(W11));
  NANDX1 G2610 (.A1(W783), .A2(W332), .ZN(W1938));
  NANDX1 G2611 (.A1(W479), .A2(W1250), .ZN(W2009));
  NANDX1 G2612 (.A1(W1990), .A2(W585), .ZN(W2007));
  NANDX1 G2613 (.A1(W651), .A2(W451), .ZN(O274));
  NANDX1 G2614 (.A1(I28), .A2(I29), .ZN(W14));
  NANDX1 G2615 (.A1(W1835), .A2(W1325), .ZN(O273));
  NANDX1 G2616 (.A1(W49), .A2(W357), .ZN(W2000));
  NANDX1 G2617 (.A1(W1178), .A2(W1937), .ZN(W1998));
  NANDX1 G2618 (.A1(W834), .A2(I134), .ZN(O271));
  NANDX1 G2619 (.A1(W564), .A2(W580), .ZN(O269));
  NANDX1 G2620 (.A1(W184), .A2(W1790), .ZN(W1991));
  NANDX1 G2621 (.A1(W745), .A2(W113), .ZN(O232));
  NANDX1 G2622 (.A1(W1093), .A2(W335), .ZN(O238));
  NANDX1 G2623 (.A1(W581), .A2(W602), .ZN(W1874));
  NANDX1 G2624 (.A1(I194), .A2(I195), .ZN(W97));
  NANDX1 G2625 (.A1(W942), .A2(W1186), .ZN(W1872));
  NANDX1 G2626 (.A1(W83), .A2(W1678), .ZN(W1871));
  NANDX1 G2627 (.A1(I196), .A2(I197), .ZN(W98));
  NANDX1 G2628 (.A1(W1135), .A2(W1526), .ZN(W1870));
  NANDX1 G2629 (.A1(W233), .A2(W99), .ZN(W1869));
  NANDX1 G2630 (.A1(W1311), .A2(W445), .ZN(O236));
  NANDX1 G2631 (.A1(W336), .A2(W502), .ZN(O233));
  NANDX1 G2632 (.A1(I29), .A2(I31), .ZN(W101));
  NANDX1 G2633 (.A1(W1593), .A2(I120), .ZN(W1889));
  NANDX1 G2634 (.A1(I40), .A2(I65), .ZN(W102));
  NANDX1 G2635 (.A1(I174), .A2(W526), .ZN(O231));
  NANDX1 G2636 (.A1(W58), .A2(I111), .ZN(W104));
  NANDX1 G2637 (.A1(W1360), .A2(W968), .ZN(W1858));
  NANDX1 G2638 (.A1(I166), .A2(I90), .ZN(W105));
  NANDX1 G2639 (.A1(W376), .A2(I9), .ZN(W1857));
  NANDX1 G2640 (.A1(W717), .A2(W216), .ZN(O229));
  NANDX1 G2641 (.A1(W454), .A2(W1403), .ZN(W1852));
  NANDX1 G2642 (.A1(I111), .A2(I116), .ZN(W106));
  NANDX1 G2643 (.A1(W62), .A2(W333), .ZN(W1851));
  NANDX1 G2644 (.A1(W1555), .A2(W568), .ZN(O247));
  NANDX1 G2645 (.A1(W149), .A2(W607), .ZN(W1937));
  NANDX1 G2646 (.A1(W1107), .A2(W761), .ZN(W1932));
  NANDX1 G2647 (.A1(W764), .A2(W331), .ZN(W1930));
  NANDX1 G2648 (.A1(W1824), .A2(W1575), .ZN(O252));
  NANDX1 G2649 (.A1(W1712), .A2(I30), .ZN(O251));
  NANDX1 G2650 (.A1(I108), .A2(I109), .ZN(W54));
  NANDX1 G2651 (.A1(I116), .A2(I117), .ZN(W58));
  NANDX1 G2652 (.A1(W1790), .A2(W1138), .ZN(W1921));
  NANDX1 G2653 (.A1(I134), .A2(I135), .ZN(W67));
  NANDX1 G2654 (.A1(I136), .A2(I137), .ZN(W68));
  NANDX1 G2655 (.A1(W1209), .A2(W1487), .ZN(W1916));
  NANDX1 G2656 (.A1(I100), .A2(I85), .ZN(W293));
  NANDX1 G2657 (.A1(W1201), .A2(W130), .ZN(W1910));
  NANDX1 G2658 (.A1(W1316), .A2(W1407), .ZN(O245));
  NANDX1 G2659 (.A1(W653), .A2(W1411), .ZN(W1905));
  NANDX1 G2660 (.A1(I144), .A2(I145), .ZN(W72));
  NANDX1 G2661 (.A1(W1701), .A2(W257), .ZN(W1902));
  NANDX1 G2662 (.A1(W303), .A2(I85), .ZN(O243));
  NANDX1 G2663 (.A1(I156), .A2(I157), .ZN(W78));
  NANDX1 G2664 (.A1(I164), .A2(I165), .ZN(W82));
  NANDX1 G2665 (.A1(I165), .A2(W995), .ZN(W1893));
  NANDX1 G2666 (.A1(W1324), .A2(W1029), .ZN(W1891));
  NANDX1 G2667 (.A1(W238), .A2(W370), .ZN(W1636));
  NANDX1 G2668 (.A1(W1113), .A2(I65), .ZN(W1631));
  NANDX1 G2669 (.A1(W33), .A2(W220), .ZN(O153));
  NANDX1 G2670 (.A1(I56), .A2(I20), .ZN(W252));
  NANDX1 G2671 (.A1(W404), .A2(W455), .ZN(O160));
  NANDX1 G2672 (.A1(W1443), .A2(W677), .ZN(O171));
  NANDX1 G2673 (.A1(W68), .A2(W129), .ZN(O6));
  NANDX1 G2674 (.A1(W164), .A2(W194), .ZN(W262));
  NANDX1 G2675 (.A1(W1411), .A2(W394), .ZN(W1667));
  NANDX1 G2676 (.A1(W27), .A2(I109), .ZN(W284));
  NANDX1 G2677 (.A1(I138), .A2(I160), .ZN(W235));
  NANDX1 G2678 (.A1(W1381), .A2(W942), .ZN(W1670));
  NANDX1 G2679 (.A1(I152), .A2(W51), .ZN(W263));
  NANDX1 G2680 (.A1(W1498), .A2(W152), .ZN(W1587));
  NANDX1 G2681 (.A1(W1341), .A2(W1085), .ZN(W1625));
  NANDX1 G2682 (.A1(W128), .A2(I39), .ZN(W288));
  NANDX1 G2683 (.A1(W544), .A2(I190), .ZN(W1593));
  NANDX1 G2684 (.A1(I40), .A2(I184), .ZN(W232));
  NANDX1 G2685 (.A1(I36), .A2(W321), .ZN(W1589));
  NANDX1 G2686 (.A1(W1224), .A2(W1537), .ZN(O173));
  NANDX1 G2687 (.A1(I191), .A2(W236), .ZN(W286));
  NANDX1 G2688 (.A1(W1363), .A2(W1020), .ZN(W1605));
  NANDX1 G2689 (.A1(I175), .A2(I98), .ZN(W269));
  NANDX1 G2690 (.A1(W39), .A2(W889), .ZN(W1591));
  NANDX1 G2691 (.A1(W99), .A2(W480), .ZN(W1592));
  NANDX1 G2692 (.A1(W1435), .A2(W628), .ZN(W1646));
  NANDX1 G2693 (.A1(W1240), .A2(W789), .ZN(O166));
  NANDX1 G2694 (.A1(I75), .A2(W52), .ZN(W242));
  NANDX1 G2695 (.A1(I109), .A2(W1420), .ZN(W1638));
  NANDX1 G2696 (.A1(W1210), .A2(W517), .ZN(O169));
  NANDX1 G2697 (.A1(W1210), .A2(W1180), .ZN(W1610));
  NANDX1 G2698 (.A1(W485), .A2(W1420), .ZN(O174));
  NANDX1 G2699 (.A1(W141), .A2(W19), .ZN(W287));
  NANDX1 G2700 (.A1(W1508), .A2(W856), .ZN(O176));
  NANDX1 G2701 (.A1(I180), .A2(W156), .ZN(W236));
  NANDX1 G2702 (.A1(W1372), .A2(W1391), .ZN(W1666));
  NANDX1 G2703 (.A1(W695), .A2(I71), .ZN(W1586));
  NANDX1 G2704 (.A1(W33), .A2(W1112), .ZN(W1615));
  NANDX1 G2705 (.A1(W83), .A2(W97), .ZN(W292));
  NANDX1 G2706 (.A1(W100), .A2(W1193), .ZN(W1651));
  NANDX1 G2707 (.A1(W221), .A2(W92), .ZN(W276));
  NANDX1 G2708 (.A1(W109), .A2(I174), .ZN(W229));
  NANDX1 G2709 (.A1(I150), .A2(W231), .ZN(W266));
  NANDX1 G2710 (.A1(I111), .A2(W249), .ZN(W265));
  NANDX1 G2711 (.A1(W344), .A2(W492), .ZN(W1678));
  NANDX1 G2712 (.A1(W621), .A2(W99), .ZN(W1674));
  NANDX1 G2713 (.A1(W232), .A2(W204), .ZN(W277));
  NANDX1 G2714 (.A1(W274), .A2(W1138), .ZN(W1612));
  NANDX1 G2715 (.A1(W1511), .A2(I31), .ZN(W1652));
  NANDX1 G2716 (.A1(I160), .A2(W4), .ZN(W259));
  NANDX1 G2717 (.A1(W889), .A2(W124), .ZN(O177));
  NANDX1 G2718 (.A1(W109), .A2(W92), .ZN(W290));
  NANDX1 G2719 (.A1(W1620), .A2(W1195), .ZN(W1654));
  NANDX1 G2720 (.A1(W826), .A2(W1181), .ZN(W1599));
  NANDX1 G2721 (.A1(W10), .A2(W191), .ZN(W240));
  NANDX1 G2722 (.A1(W835), .A2(W925), .ZN(W1618));
  NANDX1 G2723 (.A1(W866), .A2(W803), .ZN(W1603));
  NANDX1 G2724 (.A1(I31), .A2(W132), .ZN(W255));
  NANDX1 G2725 (.A1(W627), .A2(W514), .ZN(W1595));
  NANDX1 G2726 (.A1(I103), .A2(W31), .ZN(O4));
  NANDX1 G2727 (.A1(W567), .A2(W223), .ZN(W1624));
  NANDX1 G2728 (.A1(W177), .A2(I14), .ZN(W289));
  NANDX1 G2729 (.A1(W773), .A2(W1494), .ZN(W1601));
  NANDX1 G2730 (.A1(W456), .A2(W477), .ZN(O152));
  NANDX1 G2731 (.A1(W209), .A2(W222), .ZN(W264));
  INVX1 G2732 (.I(W92), .ZN(O1036));
  INVX1 G2733 (.I(I140), .ZN(W70));
  INVX1 G2734 (.I(W432), .ZN(W671));
  INVX1 G2735 (.I(W682), .ZN(W3417));
  INVX1 G2736 (.I(W3179), .ZN(O1557));
  INVX1 G2737 (.I(W369), .ZN(O1384));
  INVX1 G2738 (.I(W910), .ZN(O1035));
  INVX1 G2739 (.I(W378), .ZN(O1029));
  INVX1 G2740 (.I(I108), .ZN(W662));
  INVX1 G2741 (.I(W3893), .ZN(O1558));
  INVX1 G2742 (.I(W1595), .ZN(O1560));
  INVX1 G2743 (.I(W344), .ZN(W669));
  INVX1 G2744 (.I(I138), .ZN(W69));
  INVX1 G2745 (.I(I128), .ZN(W64));
  INVX1 G2746 (.I(I0), .ZN(W664));
  INVX1 G2747 (.I(W2642), .ZN(O1032));
  INVX1 G2748 (.I(W3528), .ZN(O1574));
  INVX1 G2749 (.I(I118), .ZN(W59));
  INVX1 G2750 (.I(W189), .ZN(W3404));
  INVX1 G2751 (.I(W2334), .ZN(O1019));
  INVX1 G2752 (.I(W157), .ZN(W326));
  INVX1 G2753 (.I(W2120), .ZN(O1334));
  INVX1 G2754 (.I(W675), .ZN(W684));
  INVX1 G2755 (.I(W3634), .ZN(O1381));
  INVX1 G2756 (.I(W1105), .ZN(O1016));
  INVX1 G2757 (.I(I124), .ZN(W62));
  INVX1 G2758 (.I(I106), .ZN(W53));
  INVX1 G2759 (.I(W1560), .ZN(O1014));
  INVX1 G2760 (.I(W1776), .ZN(O1013));
  INVX1 G2761 (.I(I132), .ZN(W270));
  INVX1 G2762 (.I(W474), .ZN(O1011));
  INVX1 G2763 (.I(W1835), .ZN(O1336));
  INVX1 G2764 (.I(I104), .ZN(W52));
  INVX1 G2765 (.I(W1202), .ZN(O1329));
  INVX1 G2766 (.I(W1625), .ZN(W3407));
  INVX1 G2767 (.I(W224), .ZN(O1022));
  INVX1 G2768 (.I(W651), .ZN(O1569));
  INVX1 G2769 (.I(W1694), .ZN(O1023));
  INVX1 G2770 (.I(I126), .ZN(W63));
  INVX1 G2771 (.I(W630), .ZN(O1024));
  INVX1 G2772 (.I(W2606), .ZN(O1323));
  INVX1 G2773 (.I(I134), .ZN(W674));
  INVX1 G2774 (.I(I78), .ZN(O1027));
  INVX1 G2775 (.I(W279), .ZN(O1382));
  INVX1 G2776 (.I(I130), .ZN(W65));
  INVX1 G2777 (.I(W3416), .ZN(O1565));
  INVX1 G2778 (.I(I132), .ZN(W66));
  INVX1 G2779 (.I(W335), .ZN(O1563));
  INVX1 G2780 (.I(I176), .ZN(W330));
  INVX1 G2781 (.I(I116), .ZN(O1062));
  INVX1 G2782 (.I(W534), .ZN(W626));
  INVX1 G2783 (.I(W1282), .ZN(W3466));
  INVX1 G2784 (.I(I60), .ZN(W628));
  INVX1 G2785 (.I(W3038), .ZN(O1065));
  INVX1 G2786 (.I(W606), .ZN(O1064));
  INVX1 G2787 (.I(W417), .ZN(W630));
  INVX1 G2788 (.I(W3207), .ZN(O1538));
  INVX1 G2789 (.I(I188), .ZN(W94));
  INVX1 G2790 (.I(W1379), .ZN(O1537));
  INVX1 G2791 (.I(W201), .ZN(W337));
  INVX1 G2792 (.I(I186), .ZN(W93));
  INVX1 G2793 (.I(W682), .ZN(O1541));
  INVX1 G2794 (.I(W3363), .ZN(O1061));
  INVX1 G2795 (.I(W1442), .ZN(O1060));
  INVX1 G2796 (.I(I182), .ZN(W91));
  INVX1 G2797 (.I(W2868), .ZN(O1059));
  INVX1 G2798 (.I(W66), .ZN(O1543));
  INVX1 G2799 (.I(W1), .ZN(W616));
  INVX1 G2800 (.I(I81), .ZN(W609));
  INVX1 G2801 (.I(W1462), .ZN(W3481));
  INVX1 G2802 (.I(W367), .ZN(W611));
  INVX1 G2803 (.I(I198), .ZN(W99));
  INVX1 G2804 (.I(W2684), .ZN(O1317));
  INVX1 G2805 (.I(I29), .ZN(O15));
  INVX1 G2806 (.I(W136), .ZN(W340));
  INVX1 G2807 (.I(W170), .ZN(W338));
  INVX1 G2808 (.I(W330), .ZN(O1058));
  INVX1 G2809 (.I(W2505), .ZN(O1387));
  INVX1 G2810 (.I(W472), .ZN(O1073));
  INVX1 G2811 (.I(W202), .ZN(W617));
  INVX1 G2812 (.I(W586), .ZN(W618));
  INVX1 G2813 (.I(W3162), .ZN(O1071));
  INVX1 G2814 (.I(W237), .ZN(W622));
  INVX1 G2815 (.I(W5), .ZN(W623));
  INVX1 G2816 (.I(I62), .ZN(W267));
  INVX1 G2817 (.I(W245), .ZN(W334));
  INVX1 G2818 (.I(I166), .ZN(W83));
  INVX1 G2819 (.I(I158), .ZN(W79));
  INVX1 G2820 (.I(I100), .ZN(W50));
  INVX1 G2821 (.I(I154), .ZN(W77));
  INVX1 G2822 (.I(W10), .ZN(W646));
  INVX1 G2823 (.I(I55), .ZN(W335));
  INVX1 G2824 (.I(W1488), .ZN(W3436));
  INVX1 G2825 (.I(I148), .ZN(W74));
  INVX1 G2826 (.I(I172), .ZN(W86));
  INVX1 G2827 (.I(W235), .ZN(W649));
  INVX1 G2828 (.I(I164), .ZN(W650));
  INVX1 G2829 (.I(I148), .ZN(W333));
  INVX1 G2830 (.I(W1063), .ZN(W3781));
  INVX1 G2831 (.I(I142), .ZN(W71));
  INVX1 G2832 (.I(I146), .ZN(W659));
  INVX1 G2833 (.I(I121), .ZN(W332));
  INVX1 G2834 (.I(W2301), .ZN(O1039));
  INVX1 G2835 (.I(W1028), .ZN(O1052));
  INVX1 G2836 (.I(W370), .ZN(O1544));
  INVX1 G2837 (.I(W3011), .ZN(O1545));
  INVX1 G2838 (.I(W3037), .ZN(O1055));
  INVX1 G2839 (.I(W2907), .ZN(W3452));
  INVX1 G2840 (.I(W4), .ZN(W634));
  INVX1 G2841 (.I(W1489), .ZN(O1321));
  INVX1 G2842 (.I(I176), .ZN(W88));
  INVX1 G2843 (.I(I126), .ZN(W637));
  INVX1 G2844 (.I(W417), .ZN(W660));
  INVX1 G2845 (.I(W307), .ZN(W638));
  INVX1 G2846 (.I(W1060), .ZN(O1050));
  INVX1 G2847 (.I(W2658), .ZN(O1049));
  INVX1 G2848 (.I(W3034), .ZN(O1385));
  INVX1 G2849 (.I(I92), .ZN(W641));
  INVX1 G2850 (.I(W375), .ZN(W642));
  INVX1 G2851 (.I(I117), .ZN(W643));
  INVX1 G2852 (.I(W3017), .ZN(O964));
  INVX1 G2853 (.I(I115), .ZN(W3324));
  INVX1 G2854 (.I(I49), .ZN(W311));
  INVX1 G2855 (.I(I32), .ZN(W16));
  INVX1 G2856 (.I(I198), .ZN(W759));
  INVX1 G2857 (.I(W161), .ZN(O26));
  INVX1 G2858 (.I(W1468), .ZN(W3320));
  INVX1 G2859 (.I(W2921), .ZN(O1615));
  INVX1 G2860 (.I(W3137), .ZN(O965));
  INVX1 G2861 (.I(I34), .ZN(W17));
  INVX1 G2862 (.I(W275), .ZN(W763));
  INVX1 G2863 (.I(W1049), .ZN(O962));
  INVX1 G2864 (.I(W1767), .ZN(O1616));
  INVX1 G2865 (.I(W22), .ZN(O1617));
  INVX1 G2866 (.I(W783), .ZN(W3314));
  INVX1 G2867 (.I(W1519), .ZN(O1618));
  INVX1 G2868 (.I(W1759), .ZN(O960));
  INVX1 G2869 (.I(W2563), .ZN(O1352));
  INVX1 G2870 (.I(W167), .ZN(W746));
  INVX1 G2871 (.I(I40), .ZN(W20));
  INVX1 G2872 (.I(W475), .ZN(O979));
  INVX1 G2873 (.I(W507), .ZN(W743));
  INVX1 G2874 (.I(W1154), .ZN(O978));
  INVX1 G2875 (.I(W405), .ZN(O1348));
  INVX1 G2876 (.I(W23), .ZN(W745));
  INVX1 G2877 (.I(W365), .ZN(O975));
  INVX1 G2878 (.I(I36), .ZN(W18));
  INVX1 G2879 (.I(I116), .ZN(O959));
  INVX1 G2880 (.I(W1125), .ZN(O1349));
  INVX1 G2881 (.I(W179), .ZN(O973));
  INVX1 G2882 (.I(W3128), .ZN(O972));
  INVX1 G2883 (.I(W1094), .ZN(O971));
  INVX1 G2884 (.I(W716), .ZN(O970));
  INVX1 G2885 (.I(W991), .ZN(O1612));
  INVX1 G2886 (.I(W64), .ZN(W752));
  INVX1 G2887 (.I(I112), .ZN(W753));
  INVX1 G2888 (.I(W272), .ZN(W299));
  INVX1 G2889 (.I(W1876), .ZN(O947));
  INVX1 G2890 (.I(W28), .ZN(W786));
  INVX1 G2891 (.I(W2344), .ZN(O1625));
  INVX1 G2892 (.I(W242), .ZN(W789));
  INVX1 G2893 (.I(W2496), .ZN(O1357));
  INVX1 G2894 (.I(W181), .ZN(W793));
  INVX1 G2895 (.I(W3132), .ZN(W3822));
  INVX1 G2896 (.I(I14), .ZN(W7));
  INVX1 G2897 (.I(W182), .ZN(W291));
  INVX1 G2898 (.I(W3360), .ZN(O1360));
  INVX1 G2899 (.I(W146), .ZN(W296));
  INVX1 G2900 (.I(W1794), .ZN(O1631));
  INVX1 G2901 (.I(W2919), .ZN(W3286));
  INVX1 G2902 (.I(W2010), .ZN(O1632));
  INVX1 G2903 (.I(W301), .ZN(W2033));
  INVX1 G2904 (.I(W1650), .ZN(O941));
  INVX1 G2905 (.I(W367), .ZN(W424));
  INVX1 G2906 (.I(W1872), .ZN(O952));
  INVX1 G2907 (.I(W207), .ZN(W767));
  INVX1 G2908 (.I(I16), .ZN(W308));
  INVX1 G2909 (.I(W2615), .ZN(O1354));
  INVX1 G2910 (.I(W636), .ZN(O1620));
  INVX1 G2911 (.I(W2937), .ZN(O956));
  INVX1 G2912 (.I(W458), .ZN(W770));
  INVX1 G2913 (.I(W102), .ZN(W771));
  INVX1 G2914 (.I(I24), .ZN(W12));
  INVX1 G2915 (.I(W789), .ZN(O1346));
  INVX1 G2916 (.I(W1068), .ZN(W3302));
  INVX1 G2917 (.I(W148), .ZN(W305));
  INVX1 G2918 (.I(W147), .ZN(W777));
  INVX1 G2919 (.I(W2556), .ZN(O950));
  INVX1 G2920 (.I(W2266), .ZN(O1366));
  INVX1 G2921 (.I(W644), .ZN(W783));
  INVX1 G2922 (.I(W2097), .ZN(O1623));
  INVX1 G2923 (.I(I92), .ZN(W46));
  INVX1 G2924 (.I(W205), .ZN(O23));
  INVX1 G2925 (.I(W2320), .ZN(O998));
  INVX1 G2926 (.I(I98), .ZN(W49));
  INVX1 G2927 (.I(I96), .ZN(W48));
  INVX1 G2928 (.I(W311), .ZN(W714));
  INVX1 G2929 (.I(W3870), .ZN(O1584));
  INVX1 G2930 (.I(I134), .ZN(W316));
  INVX1 G2931 (.I(W2142), .ZN(O996));
  INVX1 G2932 (.I(I0), .ZN(W0));
  INVX1 G2933 (.I(I88), .ZN(W44));
  INVX1 G2934 (.I(W194), .ZN(W282));
  INVX1 G2935 (.I(I86), .ZN(W43));
  INVX1 G2936 (.I(W813), .ZN(O1343));
  INVX1 G2937 (.I(W353), .ZN(O1590));
  INVX1 G2938 (.I(I82), .ZN(W41));
  INVX1 G2939 (.I(W439), .ZN(W719));
  INVX1 G2940 (.I(W1406), .ZN(O993));
  INVX1 G2941 (.I(W257), .ZN(W319));
  INVX1 G2942 (.I(W3389), .ZN(O1010));
  INVX1 G2943 (.I(W396), .ZN(W691));
  INVX1 G2944 (.I(W2269), .ZN(W4044));
  INVX1 G2945 (.I(W1538), .ZN(O1577));
  INVX1 G2946 (.I(W258), .ZN(W273));
  INVX1 G2947 (.I(W2820), .ZN(W3387));
  INVX1 G2948 (.I(W3599), .ZN(O1378));
  INVX1 G2949 (.I(I34), .ZN(W704));
  INVX1 G2950 (.I(W260), .ZN(W720));
  INVX1 G2951 (.I(W229), .ZN(O1004));
  INVX1 G2952 (.I(W162), .ZN(W318));
  INVX1 G2953 (.I(W1280), .ZN(W3380));
  INVX1 G2954 (.I(W2943), .ZN(W3379));
  INVX1 G2955 (.I(W3799), .ZN(O1579));
  INVX1 G2956 (.I(I194), .ZN(W707));
  INVX1 G2957 (.I(W3132), .ZN(O1580));
  INVX1 G2958 (.I(W154), .ZN(O1000));
  INVX1 G2959 (.I(I62), .ZN(W31));
  INVX1 G2960 (.I(W3038), .ZN(O986));
  INVX1 G2961 (.I(W1897), .ZN(O1372));
  INVX1 G2962 (.I(W3139), .ZN(O1599));
  INVX1 G2963 (.I(I68), .ZN(W34));
  INVX1 G2964 (.I(W399), .ZN(W735));
  INVX1 G2965 (.I(I123), .ZN(W736));
  INVX1 G2966 (.I(W669), .ZN(W737));
  INVX1 G2967 (.I(I66), .ZN(W33));
  INVX1 G2968 (.I(W175), .ZN(W732));
  INVX1 G2969 (.I(I132), .ZN(W313));
  INVX1 G2970 (.I(I58), .ZN(W29));
  INVX1 G2971 (.I(W67), .ZN(W740));
  INVX1 G2972 (.I(W3490), .ZN(O1345));
  INVX1 G2973 (.I(I52), .ZN(W26));
  INVX1 G2974 (.I(W2432), .ZN(W3343));
  INVX1 G2975 (.I(I46), .ZN(W23));
  INVX1 G2976 (.I(I164), .ZN(W285));
  INVX1 G2977 (.I(I76), .ZN(W38));
  INVX1 G2978 (.I(W977), .ZN(O1592));
  INVX1 G2979 (.I(W2537), .ZN(W3363));
  INVX1 G2980 (.I(W2376), .ZN(O1593));
  INVX1 G2981 (.I(W3035), .ZN(W3361));
  INVX1 G2982 (.I(W228), .ZN(W725));
  INVX1 G2983 (.I(W1331), .ZN(W3359));
  INVX1 G2984 (.I(W357), .ZN(W726));
  INVX1 G2985 (.I(W43), .ZN(W314));
  INVX1 G2986 (.I(W558), .ZN(O1337));
  INVX1 G2987 (.I(W3008), .ZN(O1595));
  INVX1 G2988 (.I(W1991), .ZN(O1596));
  INVX1 G2989 (.I(W3007), .ZN(O989));
  INVX1 G2990 (.I(I84), .ZN(W729));
  INVX1 G2991 (.I(I72), .ZN(W36));
  INVX1 G2992 (.I(W980), .ZN(O1598));
  INVX1 G2993 (.I(W142), .ZN(W3352));
  INVX1 G2994 (.I(W2376), .ZN(O1457));
  INVX1 G2995 (.I(W387), .ZN(O1190));
  INVX1 G2996 (.I(W84), .ZN(O1271));
  INVX1 G2997 (.I(W172), .ZN(W3622));
  INVX1 G2998 (.I(W2779), .ZN(W3621));
  INVX1 G2999 (.I(I150), .ZN(W169));
  INVX1 G3000 (.I(I182), .ZN(W168));
  INVX1 G3001 (.I(W1818), .ZN(O1189));
  INVX1 G3002 (.I(W233), .ZN(W484));
  INVX1 G3003 (.I(W1110), .ZN(O1272));
  INVX1 G3004 (.I(W131), .ZN(W480));
  INVX1 G3005 (.I(W922), .ZN(O1185));
  INVX1 G3006 (.I(W2911), .ZN(O1184));
  INVX1 G3007 (.I(W99), .ZN(W3614));
  INVX1 G3008 (.I(W2291), .ZN(O1458));
  INVX1 G3009 (.I(W1237), .ZN(O1459));
  INVX1 G3010 (.I(W3466), .ZN(O1181));
  INVX1 G3011 (.I(W358), .ZN(O11));
  INVX1 G3012 (.I(I110), .ZN(W492));
  INVX1 G3013 (.I(W169), .ZN(W475));
  INVX1 G3014 (.I(W111), .ZN(O1203));
  INVX1 G3015 (.I(W709), .ZN(O1450));
  INVX1 G3016 (.I(W3230), .ZN(O1451));
  INVX1 G3017 (.I(W174), .ZN(W239));
  INVX1 G3018 (.I(W3213), .ZN(O1200));
  INVX1 G3019 (.I(W261), .ZN(W402));
  INVX1 G3020 (.I(I82), .ZN(W473));
  INVX1 G3021 (.I(I26), .ZN(W395));
  INVX1 G3022 (.I(W332), .ZN(W493));
  INVX1 G3023 (.I(I74), .ZN(W394));
  INVX1 G3024 (.I(W2808), .ZN(W3631));
  INVX1 G3025 (.I(W302), .ZN(W393));
  INVX1 G3026 (.I(W1498), .ZN(O1197));
  INVX1 G3027 (.I(I54), .ZN(W175));
  INVX1 G3028 (.I(W2992), .ZN(O1194));
  INVX1 G3029 (.I(W2207), .ZN(O1193));
  INVX1 G3030 (.I(W2010), .ZN(O1408));
  INVX1 G3031 (.I(W1193), .ZN(W3587));
  INVX1 G3032 (.I(W23), .ZN(W247));
  INVX1 G3033 (.I(W333), .ZN(W506));
  INVX1 G3034 (.I(W93), .ZN(O1168));
  INVX1 G3035 (.I(W2657), .ZN(O1167));
  INVX1 G3036 (.I(W1911), .ZN(O1279));
  INVX1 G3037 (.I(W986), .ZN(W3590));
  INVX1 G3038 (.I(I104), .ZN(W161));
  INVX1 G3039 (.I(W622), .ZN(O1163));
  INVX1 G3040 (.I(W173), .ZN(O1469));
  INVX1 G3041 (.I(W123), .ZN(W157));
  INVX1 G3042 (.I(W914), .ZN(O1474));
  INVX1 G3043 (.I(W1777), .ZN(O1161));
  INVX1 G3044 (.I(W300), .ZN(O1280));
  INVX1 G3045 (.I(W205), .ZN(W515));
  INVX1 G3046 (.I(W119), .ZN(W249));
  INVX1 G3047 (.I(W252), .ZN(W518));
  INVX1 G3048 (.I(W1886), .ZN(O1476));
  INVX1 G3049 (.I(W282), .ZN(W495));
  INVX1 G3050 (.I(W634), .ZN(W3607));
  INVX1 G3051 (.I(W3774), .ZN(O1460));
  INVX1 G3052 (.I(W2911), .ZN(O1275));
  INVX1 G3053 (.I(W1046), .ZN(O1177));
  INVX1 G3054 (.I(I11), .ZN(W166));
  INVX1 G3055 (.I(I52), .ZN(W378));
  INVX1 G3056 (.I(I13), .ZN(O1463));
  INVX1 G3057 (.I(W1301), .ZN(O1176));
  INVX1 G3058 (.I(W3361), .ZN(O1449));
  INVX1 G3059 (.I(I8), .ZN(O1));
  INVX1 G3060 (.I(W1653), .ZN(O1174));
  INVX1 G3061 (.I(I132), .ZN(W243));
  INVX1 G3062 (.I(W3230), .ZN(O1465));
  INVX1 G3063 (.I(W37), .ZN(W499));
  INVX1 G3064 (.I(W2863), .ZN(O1467));
  INVX1 G3065 (.I(W44), .ZN(W500));
  INVX1 G3066 (.I(W3481), .ZN(O1468));
  INVX1 G3067 (.I(W1848), .ZN(O1233));
  INVX1 G3068 (.I(W288), .ZN(W434));
  INVX1 G3069 (.I(W3685), .ZN(O1427));
  INVX1 G3070 (.I(W308), .ZN(W437));
  INVX1 G3071 (.I(W1137), .ZN(O1415));
  INVX1 G3072 (.I(I80), .ZN(W211));
  INVX1 G3073 (.I(W68), .ZN(W208));
  INVX1 G3074 (.I(I5), .ZN(W438));
  INVX1 G3075 (.I(W375), .ZN(W439));
  INVX1 G3076 (.I(I3), .ZN(W216));
  INVX1 G3077 (.I(W117), .ZN(W207));
  INVX1 G3078 (.I(W931), .ZN(O1231));
  INVX1 G3079 (.I(W408), .ZN(W441));
  INVX1 G3080 (.I(W44), .ZN(W442));
  INVX1 G3081 (.I(W2238), .ZN(O1228));
  INVX1 G3082 (.I(W2950), .ZN(O1257));
  INVX1 G3083 (.I(W404), .ZN(W417));
  INVX1 G3084 (.I(W199), .ZN(O1432));
  INVX1 G3085 (.I(W558), .ZN(O1242));
  INVX1 G3086 (.I(W2913), .ZN(O1248));
  INVX1 G3087 (.I(I137), .ZN(W228));
  INVX1 G3088 (.I(I22), .ZN(W226));
  INVX1 G3089 (.I(W2126), .ZN(O1246));
  INVX1 G3090 (.I(W76), .ZN(W423));
  INVX1 G3091 (.I(W220), .ZN(W429));
  INVX1 G3092 (.I(W1600), .ZN(O1243));
  INVX1 G3093 (.I(W471), .ZN(W3685));
  INVX1 G3094 (.I(W1121), .ZN(O1433));
  INVX1 G3095 (.I(W2846), .ZN(O1241));
  INVX1 G3096 (.I(W1179), .ZN(O1251));
  INVX1 G3097 (.I(W3582), .ZN(O1252));
  INVX1 G3098 (.I(I144), .ZN(W432));
  INVX1 G3099 (.I(W32), .ZN(W222));
  INVX1 G3100 (.I(W940), .ZN(O1424));
  INVX1 G3101 (.I(W2887), .ZN(O1254));
  INVX1 G3102 (.I(W238), .ZN(W433));
  INVX1 G3103 (.I(W400), .ZN(W461));
  INVX1 G3104 (.I(W1553), .ZN(O1441));
  INVX1 G3105 (.I(I17), .ZN(W193));
  INVX1 G3106 (.I(W432), .ZN(W458));
  INVX1 G3107 (.I(W958), .ZN(W3708));
  INVX1 G3108 (.I(I58), .ZN(W191));
  INVX1 G3109 (.I(W6), .ZN(W460));
  INVX1 G3110 (.I(W1324), .ZN(O1213));
  INVX1 G3111 (.I(W3184), .ZN(O1212));
  INVX1 G3112 (.I(W1443), .ZN(W3654));
  INVX1 G3113 (.I(W2411), .ZN(O1445));
  INVX1 G3114 (.I(W2920), .ZN(O1210));
  INVX1 G3115 (.I(W1854), .ZN(O1209));
  INVX1 G3116 (.I(W607), .ZN(O1208));
  INVX1 G3117 (.I(W1528), .ZN(O1262));
  INVX1 G3118 (.I(W3663), .ZN(W3870));
  INVX1 G3119 (.I(W1031), .ZN(O1204));
  INVX1 G3120 (.I(W53), .ZN(W181));
  INVX1 G3121 (.I(W295), .ZN(W414));
  INVX1 G3122 (.I(W300), .ZN(O1227));
  INVX1 G3123 (.I(W230), .ZN(W443));
  INVX1 G3124 (.I(W44), .ZN(O3));
  INVX1 G3125 (.I(W2902), .ZN(W3702));
  INVX1 G3126 (.I(W1150), .ZN(O1434));
  INVX1 G3127 (.I(W2232), .ZN(O1412));
  INVX1 G3128 (.I(W334), .ZN(W449));
  INVX1 G3129 (.I(W1966), .ZN(W3661));
  INVX1 G3130 (.I(W1093), .ZN(O1160));
  INVX1 G3131 (.I(W1600), .ZN(O1436));
  INVX1 G3132 (.I(I86), .ZN(W454));
  INVX1 G3133 (.I(W3793), .ZN(O1437));
  INVX1 G3134 (.I(W1200), .ZN(O1219));
  INVX1 G3135 (.I(W174), .ZN(W200));
  INVX1 G3136 (.I(W3487), .ZN(O1218));
  INVX1 G3137 (.I(I64), .ZN(W413));
  INVX1 G3138 (.I(W1318), .ZN(O1217));
  INVX1 G3139 (.I(W3375), .ZN(O1106));
  INVX1 G3140 (.I(W3322), .ZN(O1516));
  INVX1 G3141 (.I(W509), .ZN(W3521));
  INVX1 G3142 (.I(W84), .ZN(W114));
  INVX1 G3143 (.I(W217), .ZN(O1518));
  INVX1 G3144 (.I(W1167), .ZN(O1108));
  INVX1 G3145 (.I(I78), .ZN(W113));
  INVX1 G3146 (.I(W4), .ZN(W112));
  INVX1 G3147 (.I(W2714), .ZN(O1303));
  INVX1 G3148 (.I(W1650), .ZN(O1110));
  INVX1 G3149 (.I(W2884), .ZN(O1105));
  INVX1 G3150 (.I(I118), .ZN(W584));
  INVX1 G3151 (.I(I181), .ZN(O1103));
  INVX1 G3152 (.I(W407), .ZN(W585));
  INVX1 G3153 (.I(W1499), .ZN(O1101));
  INVX1 G3154 (.I(W1573), .ZN(O1304));
  INVX1 G3155 (.I(W2745), .ZN(O1522));
  INVX1 G3156 (.I(W1271), .ZN(O1099));
  INVX1 G3157 (.I(W74), .ZN(W572));
  INVX1 G3158 (.I(I75), .ZN(W123));
  INVX1 G3159 (.I(W3442), .ZN(W3748));
  INVX1 G3160 (.I(W280), .ZN(W359));
  INVX1 G3161 (.I(W351), .ZN(W357));
  INVX1 G3162 (.I(W61), .ZN(W118));
  INVX1 G3163 (.I(I110), .ZN(O1119));
  INVX1 G3164 (.I(W446), .ZN(W569));
  INVX1 G3165 (.I(W3184), .ZN(O1117));
  INVX1 G3166 (.I(W554), .ZN(W3509));
  INVX1 G3167 (.I(W1847), .ZN(O1300));
  INVX1 G3168 (.I(I168), .ZN(W575));
  INVX1 G3169 (.I(W503), .ZN(W576));
  INVX1 G3170 (.I(I132), .ZN(W353));
  INVX1 G3171 (.I(W9), .ZN(W261));
  INVX1 G3172 (.I(W1536), .ZN(O1112));
  INVX1 G3173 (.I(I7), .ZN(W115));
  INVX1 G3174 (.I(W291), .ZN(W580));
  INVX1 G3175 (.I(W1790), .ZN(O1084));
  INVX1 G3176 (.I(W98), .ZN(W348));
  INVX1 G3177 (.I(W403), .ZN(W601));
  INVX1 G3178 (.I(W307), .ZN(W345));
  INVX1 G3179 (.I(W95), .ZN(W602));
  INVX1 G3180 (.I(W2477), .ZN(O1390));
  INVX1 G3181 (.I(W301), .ZN(W603));
  INVX1 G3182 (.I(W347), .ZN(W604));
  INVX1 G3183 (.I(W569), .ZN(W3490));
  INVX1 G3184 (.I(W381), .ZN(W598));
  INVX1 G3185 (.I(W1120), .ZN(O1312));
  INVX1 G3186 (.I(W2579), .ZN(O1313));
  INVX1 G3187 (.I(W3027), .ZN(O1314));
  INVX1 G3188 (.I(W418), .ZN(W608));
  INVX1 G3189 (.I(W398), .ZN(O1082));
  INVX1 G3190 (.I(I172), .ZN(W343));
  INVX1 G3191 (.I(W125), .ZN(W342));
  INVX1 G3192 (.I(W3170), .ZN(W3999));
  INVX1 G3193 (.I(W772), .ZN(O1093));
  INVX1 G3194 (.I(W726), .ZN(O1098));
  INVX1 G3195 (.I(W1160), .ZN(O1523));
  INVX1 G3196 (.I(W1095), .ZN(O1524));
  INVX1 G3197 (.I(W2372), .ZN(O1097));
  INVX1 G3198 (.I(W1553), .ZN(O1393));
  INVX1 G3199 (.I(W815), .ZN(O1525));
  INVX1 G3200 (.I(I124), .ZN(O1095));
  INVX1 G3201 (.I(W14), .ZN(O1094));
  INVX1 G3202 (.I(W470), .ZN(O1120));
  INVX1 G3203 (.I(W194), .ZN(W591));
  INVX1 G3204 (.I(W1300), .ZN(O1526));
  INVX1 G3205 (.I(I45), .ZN(O1306));
  INVX1 G3206 (.I(W129), .ZN(W594));
  INVX1 G3207 (.I(I123), .ZN(W108));
  INVX1 G3208 (.I(W59), .ZN(W3498));
  INVX1 G3209 (.I(W196), .ZN(W596));
  INVX1 G3210 (.I(W591), .ZN(W597));
  INVX1 G3211 (.I(W1542), .ZN(W3952));
  INVX1 G3212 (.I(W329), .ZN(W538));
  INVX1 G3213 (.I(W92), .ZN(W540));
  INVX1 G3214 (.I(I17), .ZN(W251));
  INVX1 G3215 (.I(W61), .ZN(W542));
  INVX1 G3216 (.I(W34), .ZN(W149));
  INVX1 G3217 (.I(W2737), .ZN(O1284));
  INVX1 G3218 (.I(W3055), .ZN(O1285));
  INVX1 G3219 (.I(W2533), .ZN(O1286));
  INVX1 G3220 (.I(W1378), .ZN(O1484));
  INVX1 G3221 (.I(W352), .ZN(W370));
  INVX1 G3222 (.I(W23), .ZN(W145));
  INVX1 G3223 (.I(I42), .ZN(W369));
  INVX1 G3224 (.I(W2337), .ZN(O1144));
  INVX1 G3225 (.I(W3661), .ZN(O1490));
  INVX1 G3226 (.I(W427), .ZN(W547));
  INVX1 G3227 (.I(W137), .ZN(W143));
  INVX1 G3228 (.I(W312), .ZN(W548));
  INVX1 G3229 (.I(W823), .ZN(O1480));
  INVX1 G3230 (.I(W443), .ZN(W519));
  INVX1 G3231 (.I(I95), .ZN(W522));
  INVX1 G3232 (.I(W566), .ZN(O1281));
  INVX1 G3233 (.I(W3525), .ZN(O1477));
  INVX1 G3234 (.I(W1536), .ZN(O1282));
  INVX1 G3235 (.I(W3521), .ZN(O1157));
  INVX1 G3236 (.I(W2939), .ZN(O1478));
  INVX1 G3237 (.I(W3264), .ZN(O1479));
  INVX1 G3238 (.I(W3492), .ZN(O1141));
  INVX1 G3239 (.I(W11), .ZN(W152));
  INVX1 G3240 (.I(W2369), .ZN(O1153));
  INVX1 G3241 (.I(W386), .ZN(W529));
  INVX1 G3242 (.I(W274), .ZN(W533));
  INVX1 G3243 (.I(W1740), .ZN(O1482));
  INVX1 G3244 (.I(W155), .ZN(W371));
  INVX1 G3245 (.I(W936), .ZN(O1149));
  INVX1 G3246 (.I(W2741), .ZN(W3731));
  INVX1 G3247 (.I(W3387), .ZN(O1507));
  INVX1 G3248 (.I(I62), .ZN(O1503));
  INVX1 G3249 (.I(I72), .ZN(W363));
  INVX1 G3250 (.I(I30), .ZN(W130));
  INVX1 G3251 (.I(I152), .ZN(W129));
  INVX1 G3252 (.I(W379), .ZN(W563));
  INVX1 G3253 (.I(W2320), .ZN(O1125));
  INVX1 G3254 (.I(W815), .ZN(O1294));
  INVX1 G3255 (.I(W2922), .ZN(O1124));
  INVX1 G3256 (.I(W142), .ZN(O1502));
  INVX1 G3257 (.I(W1394), .ZN(O1397));
  INVX1 G3258 (.I(W2035), .ZN(O1396));
  INVX1 G3259 (.I(I135), .ZN(W126));
  INVX1 G3260 (.I(W319), .ZN(W566));
  INVX1 G3261 (.I(W1952), .ZN(O1122));
  INVX1 G3262 (.I(W453), .ZN(O1297));
  INVX1 G3263 (.I(W261), .ZN(W567));
  INVX1 G3264 (.I(W3587), .ZN(O1510));
  INVX1 G3265 (.I(W160), .ZN(W556));
  INVX1 G3266 (.I(I158), .ZN(W141));
  INVX1 G3267 (.I(W1652), .ZN(O1140));
  INVX1 G3268 (.I(W1630), .ZN(O1288));
  INVX1 G3269 (.I(I132), .ZN(W137));
  INVX1 G3270 (.I(I50), .ZN(W550));
  INVX1 G3271 (.I(W501), .ZN(O1495));
  INVX1 G3272 (.I(W1505), .ZN(O1400));
  INVX1 G3273 (.I(W2891), .ZN(O1290));
  INVX1 G3274 (.I(W7), .ZN(W100));
  INVX1 G3275 (.I(W840), .ZN(O1496));
  INVX1 G3276 (.I(W492), .ZN(O1497));
  INVX1 G3277 (.I(I76), .ZN(W136));
  INVX1 G3278 (.I(W124), .ZN(W132));
  INVX1 G3279 (.I(W2438), .ZN(O1500));
  INVX1 G3280 (.I(W45), .ZN(W367));
  INVX1 G3281 (.I(I147), .ZN(W558));
  INVX1 G3282 (.I(I55), .ZN(W364));
  INVX1 G3283 (.I(W227), .ZN(W1598));
  INVX1 G3284 (.I(W1943), .ZN(O463));
  INVX1 G3285 (.I(W401), .ZN(W1585));
  INVX1 G3286 (.I(W582), .ZN(W2477));
  INVX1 G3287 (.I(W1998), .ZN(O461));
  INVX1 G3288 (.I(W1803), .ZN(W2474));
  INVX1 G3289 (.I(I153), .ZN(W2473));
  INVX1 G3290 (.I(W1688), .ZN(W2472));
  INVX1 G3291 (.I(W248), .ZN(O459));
  INVX1 G3292 (.I(W181), .ZN(W1590));
  INVX1 G3293 (.I(W1190), .ZN(W1594));
  INVX1 G3294 (.I(W742), .ZN(W1596));
  INVX1 G3295 (.I(W1390), .ZN(O151));
  INVX1 G3296 (.I(W1729), .ZN(W2480));
  INVX1 G3297 (.I(W1744), .ZN(O454));
  INVX1 G3298 (.I(W1303), .ZN(O452));
  INVX1 G3299 (.I(W1965), .ZN(O451));
  INVX1 G3300 (.I(W2348), .ZN(W2455));
  INVX1 G3301 (.I(W2003), .ZN(O450));
  INVX1 G3302 (.I(W587), .ZN(W2453));
  INVX1 G3303 (.I(W1032), .ZN(W2452));
  INVX1 G3304 (.I(W668), .ZN(W2448));
  INVX1 G3305 (.I(W1158), .ZN(W1604));
  INVX1 G3306 (.I(W468), .ZN(W1606));
  INVX1 G3307 (.I(W682), .ZN(W1609));
  INVX1 G3308 (.I(W409), .ZN(O155));
  INVX1 G3309 (.I(W1851), .ZN(O472));
  INVX1 G3310 (.I(W1381), .ZN(W1534));
  INVX1 G3311 (.I(W1217), .ZN(O481));
  INVX1 G3312 (.I(W61), .ZN(W1536));
  INVX1 G3313 (.I(W1150), .ZN(W2520));
  INVX1 G3314 (.I(W147), .ZN(W1537));
  INVX1 G3315 (.I(W849), .ZN(W1540));
  INVX1 G3316 (.I(W1473), .ZN(O478));
  INVX1 G3317 (.I(W737), .ZN(W1545));
  INVX1 G3318 (.I(W1341), .ZN(W1546));
  INVX1 G3319 (.I(W1472), .ZN(W2508));
  INVX1 G3320 (.I(W624), .ZN(W1548));
  INVX1 G3321 (.I(W1495), .ZN(O137));
  INVX1 G3322 (.I(W1504), .ZN(W1613));
  INVX1 G3323 (.I(W479), .ZN(W2501));
  INVX1 G3324 (.I(W1246), .ZN(W1555));
  INVX1 G3325 (.I(W951), .ZN(W2498));
  INVX1 G3326 (.I(W287), .ZN(W1563));
  INVX1 G3327 (.I(W1128), .ZN(W1564));
  INVX1 G3328 (.I(W378), .ZN(O145));
  INVX1 G3329 (.I(W1170), .ZN(W1569));
  INVX1 G3330 (.I(W1389), .ZN(W1575));
  INVX1 G3331 (.I(W396), .ZN(W1581));
  INVX1 G3332 (.I(W104), .ZN(O464));
  INVX1 G3333 (.I(W140), .ZN(W1582));
  INVX1 G3334 (.I(W2103), .ZN(W2481));
  INVX1 G3335 (.I(W46), .ZN(O415));
  INVX1 G3336 (.I(W303), .ZN(W1669));
  INVX1 G3337 (.I(W665), .ZN(O423));
  INVX1 G3338 (.I(I54), .ZN(W1672));
  INVX1 G3339 (.I(W2301), .ZN(O422));
  INVX1 G3340 (.I(W2268), .ZN(W2388));
  INVX1 G3341 (.I(W1584), .ZN(O178));
  INVX1 G3342 (.I(W949), .ZN(O419));
  INVX1 G3343 (.I(W811), .ZN(O179));
  INVX1 G3344 (.I(W1687), .ZN(O418));
  INVX1 G3345 (.I(W781), .ZN(O417));
  INVX1 G3346 (.I(W917), .ZN(O180));
  INVX1 G3347 (.I(W2226), .ZN(O416));
  INVX1 G3348 (.I(W439), .ZN(W1665));
  INVX1 G3349 (.I(W257), .ZN(W2373));
  INVX1 G3350 (.I(I137), .ZN(W2372));
  INVX1 G3351 (.I(W104), .ZN(O414));
  INVX1 G3352 (.I(I2), .ZN(W2370));
  INVX1 G3353 (.I(W331), .ZN(W1685));
  INVX1 G3354 (.I(W2324), .ZN(W2368));
  INVX1 G3355 (.I(W1235), .ZN(W1686));
  INVX1 G3356 (.I(W348), .ZN(W1687));
  INVX1 G3357 (.I(W1142), .ZN(W1688));
  INVX1 G3358 (.I(W611), .ZN(O412));
  INVX1 G3359 (.I(W1373), .ZN(O409));
  INVX1 G3360 (.I(W1601), .ZN(W1692));
  INVX1 G3361 (.I(W387), .ZN(O439));
  INVX1 G3362 (.I(W194), .ZN(W1619));
  INVX1 G3363 (.I(W1108), .ZN(O157));
  INVX1 G3364 (.I(W1455), .ZN(W1622));
  INVX1 G3365 (.I(W1522), .ZN(W2432));
  INVX1 G3366 (.I(W311), .ZN(O445));
  INVX1 G3367 (.I(I26), .ZN(O444));
  INVX1 G3368 (.I(W1452), .ZN(W2429));
  INVX1 G3369 (.I(W598), .ZN(O443));
  INVX1 G3370 (.I(W429), .ZN(O158));
  INVX1 G3371 (.I(I4), .ZN(O441));
  INVX1 G3372 (.I(W518), .ZN(W1628));
  INVX1 G3373 (.I(W1618), .ZN(W1629));
  INVX1 G3374 (.I(W1324), .ZN(W1532));
  INVX1 G3375 (.I(W2360), .ZN(W2420));
  INVX1 G3376 (.I(W304), .ZN(O161));
  INVX1 G3377 (.I(W221), .ZN(W1634));
  INVX1 G3378 (.I(W190), .ZN(W1635));
  INVX1 G3379 (.I(W589), .ZN(O162));
  INVX1 G3380 (.I(W1001), .ZN(O168));
  INVX1 G3381 (.I(W1301), .ZN(O170));
  INVX1 G3382 (.I(W505), .ZN(O430));
  INVX1 G3383 (.I(W842), .ZN(W2404));
  INVX1 G3384 (.I(W326), .ZN(W2401));
  INVX1 G3385 (.I(W845), .ZN(O172));
  INVX1 G3386 (.I(W1111), .ZN(W2608));
  INVX1 G3387 (.I(W139), .ZN(W1449));
  INVX1 G3388 (.I(W1159), .ZN(W1450));
  INVX1 G3389 (.I(W1264), .ZN(W2625));
  INVX1 G3390 (.I(W892), .ZN(W1451));
  INVX1 G3391 (.I(W932), .ZN(W1452));
  INVX1 G3392 (.I(W412), .ZN(W1453));
  INVX1 G3393 (.I(W2295), .ZN(O532));
  INVX1 G3394 (.I(W594), .ZN(O528));
  INVX1 G3395 (.I(W1570), .ZN(O527));
  INVX1 G3396 (.I(W2354), .ZN(O526));
  INVX1 G3397 (.I(W408), .ZN(O525));
  INVX1 G3398 (.I(W907), .ZN(O524));
  INVX1 G3399 (.I(W2412), .ZN(W2628));
  INVX1 G3400 (.I(W481), .ZN(W1462));
  INVX1 G3401 (.I(W179), .ZN(W2605));
  INVX1 G3402 (.I(W1323), .ZN(W1465));
  INVX1 G3403 (.I(W1375), .ZN(W2603));
  INVX1 G3404 (.I(W1174), .ZN(W1466));
  INVX1 G3405 (.I(W1394), .ZN(W1467));
  INVX1 G3406 (.I(W2212), .ZN(W2600));
  INVX1 G3407 (.I(W1186), .ZN(W1469));
  INVX1 G3408 (.I(W2559), .ZN(O520));
  INVX1 G3409 (.I(W251), .ZN(O519));
  INVX1 G3410 (.I(W1067), .ZN(W1471));
  INVX1 G3411 (.I(W221), .ZN(W2593));
  INVX1 G3412 (.I(W1113), .ZN(W1420));
  INVX1 G3413 (.I(W588), .ZN(W1405));
  INVX1 G3414 (.I(W633), .ZN(W1407));
  INVX1 G3415 (.I(W1075), .ZN(W1409));
  INVX1 G3416 (.I(W550), .ZN(W1412));
  INVX1 G3417 (.I(W300), .ZN(W2659));
  INVX1 G3418 (.I(W1503), .ZN(W2658));
  INVX1 G3419 (.I(W408), .ZN(W2657));
  INVX1 G3420 (.I(W911), .ZN(W2656));
  INVX1 G3421 (.I(W274), .ZN(W2655));
  INVX1 G3422 (.I(W759), .ZN(O549));
  INVX1 G3423 (.I(W261), .ZN(W2650));
  INVX1 G3424 (.I(W2601), .ZN(O548));
  INVX1 G3425 (.I(W1560), .ZN(O518));
  INVX1 G3426 (.I(W154), .ZN(W1421));
  INVX1 G3427 (.I(W1034), .ZN(O543));
  INVX1 G3428 (.I(W670), .ZN(O119));
  INVX1 G3429 (.I(I126), .ZN(O541));
  INVX1 G3430 (.I(I191), .ZN(W1427));
  INVX1 G3431 (.I(W2242), .ZN(O540));
  INVX1 G3432 (.I(W2166), .ZN(O539));
  INVX1 G3433 (.I(W1233), .ZN(O122));
  INVX1 G3434 (.I(W327), .ZN(O123));
  INVX1 G3435 (.I(W1870), .ZN(W2632));
  INVX1 G3436 (.I(W750), .ZN(W1443));
  INVX1 G3437 (.I(W1452), .ZN(O491));
  INVX1 G3438 (.I(W525), .ZN(W1499));
  INVX1 G3439 (.I(W361), .ZN(W1503));
  INVX1 G3440 (.I(W1204), .ZN(W1505));
  INVX1 G3441 (.I(W1806), .ZN(O498));
  INVX1 G3442 (.I(W1956), .ZN(W2556));
  INVX1 G3443 (.I(W1078), .ZN(O495));
  INVX1 G3444 (.I(W1073), .ZN(W1512));
  INVX1 G3445 (.I(W725), .ZN(W2548));
  INVX1 G3446 (.I(W1389), .ZN(W2547));
  INVX1 G3447 (.I(W1685), .ZN(O492));
  INVX1 G3448 (.I(W870), .ZN(W2545));
  INVX1 G3449 (.I(I28), .ZN(W1516));
  INVX1 G3450 (.I(W1654), .ZN(W2562));
  INVX1 G3451 (.I(I71), .ZN(W1517));
  INVX1 G3452 (.I(W1055), .ZN(O490));
  INVX1 G3453 (.I(W2129), .ZN(O489));
  INVX1 G3454 (.I(W2287), .ZN(W2538));
  INVX1 G3455 (.I(W268), .ZN(W1522));
  INVX1 G3456 (.I(W1820), .ZN(W2533));
  INVX1 G3457 (.I(W1755), .ZN(O486));
  INVX1 G3458 (.I(W168), .ZN(W1527));
  INVX1 G3459 (.I(W2516), .ZN(O485));
  INVX1 G3460 (.I(I17), .ZN(O484));
  INVX1 G3461 (.I(I122), .ZN(W2527));
  INVX1 G3462 (.I(W735), .ZN(W1530));
  INVX1 G3463 (.I(W213), .ZN(O510));
  INVX1 G3464 (.I(W340), .ZN(W1472));
  INVX1 G3465 (.I(W1802), .ZN(W2589));
  INVX1 G3466 (.I(W909), .ZN(W1475));
  INVX1 G3467 (.I(W783), .ZN(O515));
  INVX1 G3468 (.I(I30), .ZN(W1476));
  INVX1 G3469 (.I(W1275), .ZN(O127));
  INVX1 G3470 (.I(W1004), .ZN(W1478));
  INVX1 G3471 (.I(W865), .ZN(W1480));
  INVX1 G3472 (.I(W1218), .ZN(O511));
  INVX1 G3473 (.I(W719), .ZN(W1481));
  INVX1 G3474 (.I(W1737), .ZN(W2580));
  INVX1 G3475 (.I(W477), .ZN(W2579));
  INVX1 G3476 (.I(W1465), .ZN(W1695));
  INVX1 G3477 (.I(W985), .ZN(W1484));
  INVX1 G3478 (.I(W498), .ZN(O129));
  INVX1 G3479 (.I(W1644), .ZN(W2573));
  INVX1 G3480 (.I(W1387), .ZN(O507));
  INVX1 G3481 (.I(W2096), .ZN(O506));
  INVX1 G3482 (.I(I126), .ZN(O131));
  INVX1 G3483 (.I(W2157), .ZN(O504));
  INVX1 G3484 (.I(W41), .ZN(O503));
  INVX1 G3485 (.I(W1293), .ZN(W1497));
  INVX1 G3486 (.I(W319), .ZN(O500));
  INVX1 G3487 (.I(W586), .ZN(W2563));
  INVX1 G3488 (.I(W1074), .ZN(O250));
  INVX1 G3489 (.I(W1145), .ZN(W1912));
  INVX1 G3490 (.I(W284), .ZN(W2152));
  INVX1 G3491 (.I(W1569), .ZN(W2149));
  INVX1 G3492 (.I(W60), .ZN(W1917));
  INVX1 G3493 (.I(I39), .ZN(W1919));
  INVX1 G3494 (.I(W269), .ZN(W1920));
  INVX1 G3495 (.I(W530), .ZN(W2145));
  INVX1 G3496 (.I(W1419), .ZN(W2144));
  INVX1 G3497 (.I(W71), .ZN(W2142));
  INVX1 G3498 (.I(W926), .ZN(W1923));
  INVX1 G3499 (.I(W930), .ZN(O319));
  INVX1 G3500 (.I(W271), .ZN(W2139));
  INVX1 G3501 (.I(W1450), .ZN(W1911));
  INVX1 G3502 (.I(W1555), .ZN(W1926));
  INVX1 G3503 (.I(W1147), .ZN(W1927));
  INVX1 G3504 (.I(W706), .ZN(W1933));
  INVX1 G3505 (.I(W1205), .ZN(W1935));
  INVX1 G3506 (.I(W936), .ZN(O254));
  INVX1 G3507 (.I(I3), .ZN(W1942));
  INVX1 G3508 (.I(W1288), .ZN(W1944));
  INVX1 G3509 (.I(W89), .ZN(W1948));
  INVX1 G3510 (.I(W1315), .ZN(W2116));
  INVX1 G3511 (.I(W913), .ZN(O308));
  INVX1 G3512 (.I(W779), .ZN(W1957));
  INVX1 G3513 (.I(W1337), .ZN(W1958));
  INVX1 G3514 (.I(W1409), .ZN(W2175));
  INVX1 G3515 (.I(W1007), .ZN(O235));
  INVX1 G3516 (.I(W1159), .ZN(W2192));
  INVX1 G3517 (.I(W90), .ZN(W2189));
  INVX1 G3518 (.I(W957), .ZN(O237));
  INVX1 G3519 (.I(W206), .ZN(W1876));
  INVX1 G3520 (.I(W972), .ZN(W2183));
  INVX1 G3521 (.I(W473), .ZN(W2182));
  INVX1 G3522 (.I(W1325), .ZN(O331));
  INVX1 G3523 (.I(W1289), .ZN(W2179));
  INVX1 G3524 (.I(W183), .ZN(W2178));
  INVX1 G3525 (.I(W328), .ZN(W1885));
  INVX1 G3526 (.I(W1600), .ZN(W1887));
  INVX1 G3527 (.I(W175), .ZN(W2112));
  INVX1 G3528 (.I(W920), .ZN(W1892));
  INVX1 G3529 (.I(W1272), .ZN(W2170));
  INVX1 G3530 (.I(W371), .ZN(W1895));
  INVX1 G3531 (.I(W67), .ZN(W1896));
  INVX1 G3532 (.I(W1631), .ZN(W1897));
  INVX1 G3533 (.I(W858), .ZN(O242));
  INVX1 G3534 (.I(W1886), .ZN(W1899));
  INVX1 G3535 (.I(W1067), .ZN(O323));
  INVX1 G3536 (.I(W740), .ZN(W1903));
  INVX1 G3537 (.I(I51), .ZN(W1906));
  INVX1 G3538 (.I(W451), .ZN(W2156));
  INVX1 G3539 (.I(W517), .ZN(W2155));
  INVX1 G3540 (.I(W1821), .ZN(W2055));
  INVX1 G3541 (.I(W1548), .ZN(O268));
  INVX1 G3542 (.I(W664), .ZN(W2078));
  INVX1 G3543 (.I(W1937), .ZN(O297));
  INVX1 G3544 (.I(W1542), .ZN(O270));
  INVX1 G3545 (.I(W941), .ZN(W1996));
  INVX1 G3546 (.I(W723), .ZN(W2067));
  INVX1 G3547 (.I(W1862), .ZN(W2001));
  INVX1 G3548 (.I(W775), .ZN(W2002));
  INVX1 G3549 (.I(I71), .ZN(O293));
  INVX1 G3550 (.I(I20), .ZN(W2003));
  INVX1 G3551 (.I(W846), .ZN(W2060));
  INVX1 G3552 (.I(W1244), .ZN(W2010));
  INVX1 G3553 (.I(W1064), .ZN(W2080));
  INVX1 G3554 (.I(W388), .ZN(O288));
  INVX1 G3555 (.I(W262), .ZN(W2013));
  INVX1 G3556 (.I(W852), .ZN(W2016));
  INVX1 G3557 (.I(W677), .ZN(W2022));
  INVX1 G3558 (.I(W79), .ZN(O283));
  INVX1 G3559 (.I(W1318), .ZN(W2026));
  INVX1 G3560 (.I(W715), .ZN(O282));
  INVX1 G3561 (.I(W1725), .ZN(W2041));
  INVX1 G3562 (.I(W1330), .ZN(W2029));
  INVX1 G3563 (.I(W340), .ZN(O280));
  INVX1 G3564 (.I(W1864), .ZN(O278));
  INVX1 G3565 (.I(W1996), .ZN(W2037));
  INVX1 G3566 (.I(W387), .ZN(W2095));
  INVX1 G3567 (.I(W251), .ZN(W1960));
  INVX1 G3568 (.I(W1887), .ZN(W1961));
  INVX1 G3569 (.I(W1830), .ZN(O304));
  INVX1 G3570 (.I(W504), .ZN(W2107));
  INVX1 G3571 (.I(W354), .ZN(O262));
  INVX1 G3572 (.I(W1445), .ZN(W1965));
  INVX1 G3573 (.I(W171), .ZN(W2103));
  INVX1 G3574 (.I(W286), .ZN(W2102));
  INVX1 G3575 (.I(W827), .ZN(W1967));
  INVX1 G3576 (.I(W1774), .ZN(O263));
  INVX1 G3577 (.I(W1902), .ZN(W2097));
  INVX1 G3578 (.I(I75), .ZN(W2096));
  INVX1 G3579 (.I(W204), .ZN(O234));
  INVX1 G3580 (.I(W1349), .ZN(O265));
  INVX1 G3581 (.I(W91), .ZN(W1973));
  INVX1 G3582 (.I(W251), .ZN(W1976));
  INVX1 G3583 (.I(W989), .ZN(O301));
  INVX1 G3584 (.I(W1638), .ZN(W1978));
  INVX1 G3585 (.I(I42), .ZN(W1979));
  INVX1 G3586 (.I(W821), .ZN(W2086));
  INVX1 G3587 (.I(W1780), .ZN(O267));
  INVX1 G3588 (.I(W1787), .ZN(W2084));
  INVX1 G3589 (.I(I19), .ZN(W1982));
  INVX1 G3590 (.I(W557), .ZN(W1984));
  INVX1 G3591 (.I(W1288), .ZN(W2293));
  INVX1 G3592 (.I(W343), .ZN(W2311));
  INVX1 G3593 (.I(W774), .ZN(W2310));
  INVX1 G3594 (.I(W1006), .ZN(W1755));
  INVX1 G3595 (.I(W131), .ZN(W2306));
  INVX1 G3596 (.I(W1830), .ZN(W2305));
  INVX1 G3597 (.I(W1360), .ZN(W1761));
  INVX1 G3598 (.I(W1311), .ZN(W2301));
  INVX1 G3599 (.I(W53), .ZN(O386));
  INVX1 G3600 (.I(W823), .ZN(O202));
  INVX1 G3601 (.I(W1167), .ZN(O384));
  INVX1 G3602 (.I(W1411), .ZN(W2295));
  INVX1 G3603 (.I(W85), .ZN(W2294));
  INVX1 G3604 (.I(W2222), .ZN(O392));
  INVX1 G3605 (.I(W2101), .ZN(W2292));
  INVX1 G3606 (.I(I82), .ZN(W2291));
  INVX1 G3607 (.I(W910), .ZN(W1766));
  INVX1 G3608 (.I(W1490), .ZN(W1770));
  INVX1 G3609 (.I(W1269), .ZN(W1772));
  INVX1 G3610 (.I(W269), .ZN(O379));
  INVX1 G3611 (.I(W1822), .ZN(O378));
  INVX1 G3612 (.I(W1598), .ZN(W1774));
  INVX1 G3613 (.I(W691), .ZN(W1775));
  INVX1 G3614 (.I(W1722), .ZN(W1776));
  INVX1 G3615 (.I(W164), .ZN(W2278));
  INVX1 G3616 (.I(W844), .ZN(W1779));
  INVX1 G3617 (.I(W727), .ZN(W1723));
  INVX1 G3618 (.I(W1383), .ZN(W1697));
  INVX1 G3619 (.I(I28), .ZN(W2351));
  INVX1 G3620 (.I(W337), .ZN(W2350));
  INVX1 G3621 (.I(W1238), .ZN(O403));
  INVX1 G3622 (.I(W1576), .ZN(W2347));
  INVX1 G3623 (.I(W1335), .ZN(W1712));
  INVX1 G3624 (.I(W1624), .ZN(W1715));
  INVX1 G3625 (.I(W1278), .ZN(O400));
  INVX1 G3626 (.I(I49), .ZN(W2341));
  INVX1 G3627 (.I(W500), .ZN(W1716));
  INVX1 G3628 (.I(I115), .ZN(W1719));
  INVX1 G3629 (.I(W5), .ZN(O193));
  INVX1 G3630 (.I(W251), .ZN(W1784));
  INVX1 G3631 (.I(W821), .ZN(W2335));
  INVX1 G3632 (.I(W292), .ZN(W2334));
  INVX1 G3633 (.I(W1601), .ZN(O194));
  INVX1 G3634 (.I(W379), .ZN(O398));
  INVX1 G3635 (.I(W425), .ZN(W1726));
  INVX1 G3636 (.I(W515), .ZN(W2324));
  INVX1 G3637 (.I(W760), .ZN(W1738));
  INVX1 G3638 (.I(W1564), .ZN(O393));
  INVX1 G3639 (.I(I137), .ZN(W1746));
  INVX1 G3640 (.I(W476), .ZN(W2316));
  INVX1 G3641 (.I(W2156), .ZN(W2315));
  INVX1 G3642 (.I(W1772), .ZN(O222));
  INVX1 G3643 (.I(W138), .ZN(W1820));
  INVX1 G3644 (.I(W2069), .ZN(O358));
  INVX1 G3645 (.I(W148), .ZN(W1823));
  INVX1 G3646 (.I(W980), .ZN(W2231));
  INVX1 G3647 (.I(W389), .ZN(W1825));
  INVX1 G3648 (.I(W1407), .ZN(O220));
  INVX1 G3649 (.I(W74), .ZN(W1829));
  INVX1 G3650 (.I(W1739), .ZN(W1832));
  INVX1 G3651 (.I(W667), .ZN(O221));
  INVX1 G3652 (.I(W859), .ZN(W1834));
  INVX1 G3653 (.I(W283), .ZN(W2222));
  INVX1 G3654 (.I(W732), .ZN(W1835));
  INVX1 G3655 (.I(W1396), .ZN(O360));
  INVX1 G3656 (.I(I81), .ZN(W1839));
  INVX1 G3657 (.I(W534), .ZN(O223));
  INVX1 G3658 (.I(W710), .ZN(W1842));
  INVX1 G3659 (.I(W551), .ZN(O347));
  INVX1 G3660 (.I(W475), .ZN(W1847));
  INVX1 G3661 (.I(W1062), .ZN(O228));
  INVX1 G3662 (.I(W1364), .ZN(O343));
  INVX1 G3663 (.I(W1268), .ZN(W2207));
  INVX1 G3664 (.I(I40), .ZN(W2203));
  INVX1 G3665 (.I(W567), .ZN(O230));
  INVX1 G3666 (.I(W614), .ZN(O340));
  INVX1 G3667 (.I(W574), .ZN(W1862));
  INVX1 G3668 (.I(W25), .ZN(W2255));
  INVX1 G3669 (.I(W337), .ZN(O372));
  INVX1 G3670 (.I(W1684), .ZN(O371));
  INVX1 G3671 (.I(W1349), .ZN(W1787));
  INVX1 G3672 (.I(W304), .ZN(O370));
  INVX1 G3673 (.I(W960), .ZN(O209));
  INVX1 G3674 (.I(W922), .ZN(W2266));
  INVX1 G3675 (.I(W1416), .ZN(W1795));
  INVX1 G3676 (.I(W265), .ZN(O367));
  INVX1 G3677 (.I(W1373), .ZN(W2263));
  INVX1 G3678 (.I(W1907), .ZN(W2262));
  INVX1 G3679 (.I(W46), .ZN(W1800));
  INVX1 G3680 (.I(W471), .ZN(O211));
  INVX1 G3681 (.I(W843), .ZN(O555));
  INVX1 G3682 (.I(W184), .ZN(W2254));
  INVX1 G3683 (.I(W563), .ZN(W2253));
  INVX1 G3684 (.I(W2210), .ZN(W2252));
  INVX1 G3685 (.I(W346), .ZN(W1805));
  INVX1 G3686 (.I(W526), .ZN(O212));
  INVX1 G3687 (.I(W1780), .ZN(W2248));
  INVX1 G3688 (.I(I111), .ZN(W1812));
  INVX1 G3689 (.I(W640), .ZN(O362));
  INVX1 G3690 (.I(W1110), .ZN(O361));
  INVX1 G3691 (.I(W982), .ZN(W1814));
  INVX1 G3692 (.I(W1564), .ZN(W1819));
  INVX1 G3693 (.I(W1974), .ZN(O788));
  INVX1 G3694 (.I(W105), .ZN(O50));
  INVX1 G3695 (.I(W2426), .ZN(O800));
  INVX1 G3696 (.I(W2065), .ZN(O799));
  INVX1 G3697 (.I(W954), .ZN(W3089));
  INVX1 G3698 (.I(W2597), .ZN(W3084));
  INVX1 G3699 (.I(W398), .ZN(W1002));
  INVX1 G3700 (.I(W825), .ZN(W1004));
  INVX1 G3701 (.I(W97), .ZN(W1006));
  INVX1 G3702 (.I(W2380), .ZN(O791));
  INVX1 G3703 (.I(W864), .ZN(O790));
  INVX1 G3704 (.I(W710), .ZN(W1007));
  INVX1 G3705 (.I(W958), .ZN(O789));
  INVX1 G3706 (.I(W488), .ZN(W989));
  INVX1 G3707 (.I(W2295), .ZN(W3074));
  INVX1 G3708 (.I(W2241), .ZN(O787));
  INVX1 G3709 (.I(I132), .ZN(O52));
  INVX1 G3710 (.I(W1752), .ZN(O784));
  INVX1 G3711 (.I(W773), .ZN(O783));
  INVX1 G3712 (.I(W853), .ZN(W1012));
  INVX1 G3713 (.I(W2129), .ZN(O781));
  INVX1 G3714 (.I(W969), .ZN(W1017));
  INVX1 G3715 (.I(W923), .ZN(W1018));
  INVX1 G3716 (.I(W472), .ZN(W1019));
  INVX1 G3717 (.I(W1), .ZN(W1023));
  INVX1 G3718 (.I(W955), .ZN(W1025));
  INVX1 G3719 (.I(W298), .ZN(W973));
  INVX1 G3720 (.I(I186), .ZN(W957));
  INVX1 G3721 (.I(W87), .ZN(W3129));
  INVX1 G3722 (.I(I166), .ZN(W3128));
  INVX1 G3723 (.I(W1702), .ZN(O822));
  INVX1 G3724 (.I(W2719), .ZN(O821));
  INVX1 G3725 (.I(W2659), .ZN(W3124));
  INVX1 G3726 (.I(W1930), .ZN(O819));
  INVX1 G3727 (.I(W1239), .ZN(W3120));
  INVX1 G3728 (.I(W699), .ZN(W966));
  INVX1 G3729 (.I(W939), .ZN(O817));
  INVX1 G3730 (.I(W868), .ZN(W968));
  INVX1 G3731 (.I(W476), .ZN(W969));
  INVX1 G3732 (.I(W802), .ZN(O775));
  INVX1 G3733 (.I(W2352), .ZN(W3114));
  INVX1 G3734 (.I(I24), .ZN(O48));
  INVX1 G3735 (.I(W748), .ZN(W976));
  INVX1 G3736 (.I(I142), .ZN(W979));
  INVX1 G3737 (.I(W1839), .ZN(O809));
  INVX1 G3738 (.I(W2092), .ZN(W3105));
  INVX1 G3739 (.I(W32), .ZN(W984));
  INVX1 G3740 (.I(W2551), .ZN(O808));
  INVX1 G3741 (.I(W2627), .ZN(O807));
  INVX1 G3742 (.I(W2142), .ZN(O806));
  INVX1 G3743 (.I(W1228), .ZN(W3099));
  INVX1 G3744 (.I(I174), .ZN(W988));
  INVX1 G3745 (.I(W2409), .ZN(O748));
  INVX1 G3746 (.I(W2717), .ZN(W3019));
  INVX1 G3747 (.I(W2077), .ZN(O756));
  INVX1 G3748 (.I(W2051), .ZN(W3017));
  INVX1 G3749 (.I(W300), .ZN(W1061));
  INVX1 G3750 (.I(W110), .ZN(W1063));
  INVX1 G3751 (.I(W1564), .ZN(W3013));
  INVX1 G3752 (.I(W1361), .ZN(O753));
  INVX1 G3753 (.I(W1475), .ZN(W3011));
  INVX1 G3754 (.I(W2198), .ZN(O752));
  INVX1 G3755 (.I(I45), .ZN(W1067));
  INVX1 G3756 (.I(W599), .ZN(W1070));
  INVX1 G3757 (.I(I136), .ZN(W1071));
  INVX1 G3758 (.I(W1384), .ZN(W3020));
  INVX1 G3759 (.I(W722), .ZN(O747));
  INVX1 G3760 (.I(W2460), .ZN(O746));
  INVX1 G3761 (.I(W989), .ZN(O745));
  INVX1 G3762 (.I(W377), .ZN(W1075));
  INVX1 G3763 (.I(W752), .ZN(W2997));
  INVX1 G3764 (.I(W2018), .ZN(W2996));
  INVX1 G3765 (.I(W1084), .ZN(O741));
  INVX1 G3766 (.I(W1870), .ZN(O740));
  INVX1 G3767 (.I(W632), .ZN(O738));
  INVX1 G3768 (.I(W749), .ZN(W1083));
  INVX1 G3769 (.I(W743), .ZN(O737));
  INVX1 G3770 (.I(W579), .ZN(W1085));
  INVX1 G3771 (.I(W2934), .ZN(O768));
  INVX1 G3772 (.I(W2516), .ZN(W3056));
  INVX1 G3773 (.I(W523), .ZN(W3055));
  INVX1 G3774 (.I(W1012), .ZN(W1029));
  INVX1 G3775 (.I(W2081), .ZN(W3049));
  INVX1 G3776 (.I(W786), .ZN(W1031));
  INVX1 G3777 (.I(W808), .ZN(W1036));
  INVX1 G3778 (.I(W699), .ZN(W1037));
  INVX1 G3779 (.I(I146), .ZN(O56));
  INVX1 G3780 (.I(W35), .ZN(W1040));
  INVX1 G3781 (.I(W464), .ZN(W1041));
  INVX1 G3782 (.I(W332), .ZN(W3042));
  INVX1 G3783 (.I(W1910), .ZN(O769));
  INVX1 G3784 (.I(W568), .ZN(O47));
  INVX1 G3785 (.I(W1239), .ZN(W3038));
  INVX1 G3786 (.I(W289), .ZN(W1045));
  INVX1 G3787 (.I(W1511), .ZN(O767));
  INVX1 G3788 (.I(W458), .ZN(W1046));
  INVX1 G3789 (.I(W685), .ZN(W1047));
  INVX1 G3790 (.I(W544), .ZN(W1049));
  INVX1 G3791 (.I(W631), .ZN(O764));
  INVX1 G3792 (.I(W524), .ZN(O763));
  INVX1 G3793 (.I(W287), .ZN(W1051));
  INVX1 G3794 (.I(I114), .ZN(W1053));
  INVX1 G3795 (.I(W236), .ZN(O59));
  INVX1 G3796 (.I(W44), .ZN(W867));
  INVX1 G3797 (.I(W57), .ZN(W849));
  INVX1 G3798 (.I(W854), .ZN(W3243));
  INVX1 G3799 (.I(W2171), .ZN(W3242));
  INVX1 G3800 (.I(W805), .ZN(O35));
  INVX1 G3801 (.I(W987), .ZN(W3239));
  INVX1 G3802 (.I(W602), .ZN(W853));
  INVX1 G3803 (.I(W245), .ZN(W857));
  INVX1 G3804 (.I(W29), .ZN(W858));
  INVX1 G3805 (.I(W1136), .ZN(O901));
  INVX1 G3806 (.I(W8), .ZN(W859));
  INVX1 G3807 (.I(W2449), .ZN(O899));
  INVX1 G3808 (.I(W647), .ZN(W865));
  INVX1 G3809 (.I(W1684), .ZN(O910));
  INVX1 G3810 (.I(W927), .ZN(O895));
  INVX1 G3811 (.I(W670), .ZN(W869));
  INVX1 G3812 (.I(W2733), .ZN(O893));
  INVX1 G3813 (.I(W3162), .ZN(O892));
  INVX1 G3814 (.I(W269), .ZN(O36));
  INVX1 G3815 (.I(W692), .ZN(O891));
  INVX1 G3816 (.I(I85), .ZN(W875));
  INVX1 G3817 (.I(W276), .ZN(W877));
  INVX1 G3818 (.I(I137), .ZN(W881));
  INVX1 G3819 (.I(W3188), .ZN(W3214));
  INVX1 G3820 (.I(W751), .ZN(W884));
  INVX1 G3821 (.I(W329), .ZN(O884));
  INVX1 G3822 (.I(W501), .ZN(W821));
  INVX1 G3823 (.I(W675), .ZN(W802));
  INVX1 G3824 (.I(I88), .ZN(W803));
  INVX1 G3825 (.I(W2828), .ZN(W3278));
  INVX1 G3826 (.I(W812), .ZN(O933));
  INVX1 G3827 (.I(W241), .ZN(W812));
  INVX1 G3828 (.I(W2066), .ZN(O931));
  INVX1 G3829 (.I(I21), .ZN(W813));
  INVX1 G3830 (.I(W2658), .ZN(O930));
  INVX1 G3831 (.I(I48), .ZN(W814));
  INVX1 G3832 (.I(W505), .ZN(W816));
  INVX1 G3833 (.I(W538), .ZN(O926));
  INVX1 G3834 (.I(W621), .ZN(O32));
  INVX1 G3835 (.I(W2411), .ZN(O883));
  INVX1 G3836 (.I(W282), .ZN(W3263));
  INVX1 G3837 (.I(W366), .ZN(O33));
  INVX1 G3838 (.I(I66), .ZN(W832));
  INVX1 G3839 (.I(I108), .ZN(W833));
  INVX1 G3840 (.I(W1362), .ZN(O918));
  INVX1 G3841 (.I(W1246), .ZN(W3254));
  INVX1 G3842 (.I(W156), .ZN(W836));
  INVX1 G3843 (.I(W677), .ZN(W837));
  INVX1 G3844 (.I(W673), .ZN(W838));
  INVX1 G3845 (.I(W460), .ZN(W844));
  INVX1 G3846 (.I(W123), .ZN(W3249));
  INVX1 G3847 (.I(W55), .ZN(O44));
  INVX1 G3848 (.I(W1383), .ZN(W3168));
  INVX1 G3849 (.I(W847), .ZN(W924));
  INVX1 G3850 (.I(W208), .ZN(O852));
  INVX1 G3851 (.I(W1185), .ZN(W3165));
  INVX1 G3852 (.I(W699), .ZN(W926));
  INVX1 G3853 (.I(W2014), .ZN(O850));
  INVX1 G3854 (.I(W432), .ZN(W927));
  INVX1 G3855 (.I(I62), .ZN(W3161));
  INVX1 G3856 (.I(W861), .ZN(O847));
  INVX1 G3857 (.I(W1467), .ZN(O844));
  INVX1 G3858 (.I(W908), .ZN(O842));
  INVX1 G3859 (.I(W516), .ZN(W935));
  INVX1 G3860 (.I(W467), .ZN(W3169));
  INVX1 G3861 (.I(W505), .ZN(W943));
  INVX1 G3862 (.I(W465), .ZN(W944));
  INVX1 G3863 (.I(W903), .ZN(O45));
  INVX1 G3864 (.I(W1762), .ZN(O833));
  INVX1 G3865 (.I(W587), .ZN(O832));
  INVX1 G3866 (.I(I84), .ZN(W948));
  INVX1 G3867 (.I(W414), .ZN(W950));
  INVX1 G3868 (.I(W408), .ZN(W951));
  INVX1 G3869 (.I(W1988), .ZN(W3137));
  INVX1 G3870 (.I(W1098), .ZN(O829));
  INVX1 G3871 (.I(W891), .ZN(W952));
  INVX1 G3872 (.I(W931), .ZN(W955));
  INVX1 G3873 (.I(W861), .ZN(O41));
  INVX1 G3874 (.I(W2041), .ZN(O881));
  INVX1 G3875 (.I(W376), .ZN(W3207));
  INVX1 G3876 (.I(W1751), .ZN(O880));
  INVX1 G3877 (.I(W787), .ZN(O879));
  INVX1 G3878 (.I(W558), .ZN(O878));
  INVX1 G3879 (.I(W21), .ZN(W886));
  INVX1 G3880 (.I(W1756), .ZN(W3200));
  INVX1 G3881 (.I(W2918), .ZN(W3198));
  INVX1 G3882 (.I(W1553), .ZN(O873));
  INVX1 G3883 (.I(W84), .ZN(W895));
  INVX1 G3884 (.I(W1973), .ZN(O868));
  INVX1 G3885 (.I(W474), .ZN(W903));
  INVX1 G3886 (.I(W2336), .ZN(W2984));
  INVX1 G3887 (.I(W344), .ZN(W905));
  INVX1 G3888 (.I(W1869), .ZN(W3184));
  INVX1 G3889 (.I(W879), .ZN(W909));
  INVX1 G3890 (.I(W168), .ZN(O863));
  INVX1 G3891 (.I(I197), .ZN(W910));
  INVX1 G3892 (.I(W100), .ZN(W913));
  INVX1 G3893 (.I(W841), .ZN(W914));
  INVX1 G3894 (.I(W412), .ZN(W915));
  INVX1 G3895 (.I(I152), .ZN(W917));
  INVX1 G3896 (.I(W393), .ZN(W923));
  INVX1 G3897 (.I(W944), .ZN(W3170));
  INVX1 G3898 (.I(W324), .ZN(W1308));
  INVX1 G3899 (.I(W812), .ZN(W1289));
  INVX1 G3900 (.I(W601), .ZN(O95));
  INVX1 G3901 (.I(W1063), .ZN(W1292));
  INVX1 G3902 (.I(W1575), .ZN(O622));
  INVX1 G3903 (.I(W75), .ZN(W1293));
  INVX1 G3904 (.I(I27), .ZN(W1298));
  INVX1 G3905 (.I(W1288), .ZN(W1299));
  INVX1 G3906 (.I(W2519), .ZN(W2774));
  INVX1 G3907 (.I(W929), .ZN(O97));
  INVX1 G3908 (.I(W2094), .ZN(O616));
  INVX1 G3909 (.I(W771), .ZN(W1304));
  INVX1 G3910 (.I(W62), .ZN(W1305));
  INVX1 G3911 (.I(W18), .ZN(W1288));
  INVX1 G3912 (.I(W1134), .ZN(O98));
  INVX1 G3913 (.I(W706), .ZN(O99));
  INVX1 G3914 (.I(W2203), .ZN(W2764));
  INVX1 G3915 (.I(W299), .ZN(W2763));
  INVX1 G3916 (.I(W2), .ZN(O612));
  INVX1 G3917 (.I(W1165), .ZN(O100));
  INVX1 G3918 (.I(W1089), .ZN(W1314));
  INVX1 G3919 (.I(W2472), .ZN(O608));
  INVX1 G3920 (.I(W34), .ZN(W2756));
  INVX1 G3921 (.I(W668), .ZN(W2755));
  INVX1 G3922 (.I(W648), .ZN(W1318));
  INVX1 G3923 (.I(W1145), .ZN(W1322));
  INVX1 G3924 (.I(I66), .ZN(W1269));
  INVX1 G3925 (.I(I126), .ZN(O87));
  INVX1 G3926 (.I(W263), .ZN(W1248));
  INVX1 G3927 (.I(W2441), .ZN(W2821));
  INVX1 G3928 (.I(W53), .ZN(W1250));
  INVX1 G3929 (.I(W677), .ZN(O89));
  INVX1 G3930 (.I(W2764), .ZN(O650));
  INVX1 G3931 (.I(W1131), .ZN(O648));
  INVX1 G3932 (.I(W2563), .ZN(W2813));
  INVX1 G3933 (.I(W245), .ZN(W1262));
  INVX1 G3934 (.I(W723), .ZN(W1263));
  INVX1 G3935 (.I(W610), .ZN(O642));
  INVX1 G3936 (.I(I66), .ZN(W1267));
  INVX1 G3937 (.I(W794), .ZN(W1323));
  INVX1 G3938 (.I(W540), .ZN(W1270));
  INVX1 G3939 (.I(W1024), .ZN(W1279));
  INVX1 G3940 (.I(W662), .ZN(O635));
  INVX1 G3941 (.I(W2754), .ZN(O633));
  INVX1 G3942 (.I(W2357), .ZN(O632));
  INVX1 G3943 (.I(W2009), .ZN(O631));
  INVX1 G3944 (.I(W752), .ZN(W1282));
  INVX1 G3945 (.I(W960), .ZN(O93));
  INVX1 G3946 (.I(W972), .ZN(W1285));
  INVX1 G3947 (.I(W1036), .ZN(W1286));
  INVX1 G3948 (.I(W2781), .ZN(W2787));
  INVX1 G3949 (.I(W584), .ZN(W2691));
  INVX1 G3950 (.I(W393), .ZN(O584));
  INVX1 G3951 (.I(W557), .ZN(W1363));
  INVX1 G3952 (.I(I171), .ZN(O109));
  INVX1 G3953 (.I(W658), .ZN(O579));
  INVX1 G3954 (.I(W871), .ZN(W1377));
  INVX1 G3955 (.I(I18), .ZN(W1379));
  INVX1 G3956 (.I(W870), .ZN(W1380));
  INVX1 G3957 (.I(I140), .ZN(O577));
  INVX1 G3958 (.I(W1180), .ZN(O576));
  INVX1 G3959 (.I(W804), .ZN(W2697));
  INVX1 G3960 (.I(W1457), .ZN(O575));
  INVX1 G3961 (.I(W2148), .ZN(O571));
  INVX1 G3962 (.I(W833), .ZN(W1362));
  INVX1 G3963 (.I(W854), .ZN(W1385));
  INVX1 G3964 (.I(W79), .ZN(W1389));
  INVX1 G3965 (.I(I120), .ZN(O565));
  INVX1 G3966 (.I(W269), .ZN(W2678));
  INVX1 G3967 (.I(W985), .ZN(W2677));
  INVX1 G3968 (.I(W40), .ZN(W1398));
  INVX1 G3969 (.I(I90), .ZN(O561));
  INVX1 G3970 (.I(W1127), .ZN(W2673));
  INVX1 G3971 (.I(W1296), .ZN(O114));
  INVX1 G3972 (.I(W2615), .ZN(O559));
  INVX1 G3973 (.I(W729), .ZN(O557));
  INVX1 G3974 (.I(W477), .ZN(W1402));
  INVX1 G3975 (.I(W2623), .ZN(O595));
  INVX1 G3976 (.I(W380), .ZN(W1324));
  INVX1 G3977 (.I(W294), .ZN(W2747));
  INVX1 G3978 (.I(W1013), .ZN(W1325));
  INVX1 G3979 (.I(W525), .ZN(O104));
  INVX1 G3980 (.I(W229), .ZN(W2744));
  INVX1 G3981 (.I(W1424), .ZN(O601));
  INVX1 G3982 (.I(W584), .ZN(W1329));
  INVX1 G3983 (.I(W982), .ZN(O600));
  INVX1 G3984 (.I(W75), .ZN(W1331));
  INVX1 G3985 (.I(W510), .ZN(W1334));
  INVX1 G3986 (.I(W1029), .ZN(W1337));
  INVX1 G3987 (.I(W852), .ZN(O596));
  INVX1 G3988 (.I(W69), .ZN(O651));
  INVX1 G3989 (.I(W1121), .ZN(W2730));
  INVX1 G3990 (.I(W529), .ZN(O591));
  INVX1 G3991 (.I(W750), .ZN(W1347));
  INVX1 G3992 (.I(W49), .ZN(W1348));
  INVX1 G3993 (.I(W595), .ZN(W1350));
  INVX1 G3994 (.I(W330), .ZN(W1352));
  INVX1 G3995 (.I(I166), .ZN(O588));
  INVX1 G3996 (.I(W2368), .ZN(W2717));
  INVX1 G3997 (.I(W1716), .ZN(O587));
  INVX1 G3998 (.I(W797), .ZN(W1361));
  INVX1 G3999 (.I(W1452), .ZN(W2713));
  INVX1 G4000 (.I(W2154), .ZN(W2927));
  INVX1 G4001 (.I(W218), .ZN(W1116));
  INVX1 G4002 (.I(W0), .ZN(W1117));
  INVX1 G4003 (.I(W463), .ZN(W1118));
  INVX1 G4004 (.I(I26), .ZN(W1119));
  INVX1 G4005 (.I(W849), .ZN(W1121));
  INVX1 G4006 (.I(W683), .ZN(W1124));
  INVX1 G4007 (.I(I66), .ZN(W1127));
  INVX1 G4008 (.I(W1582), .ZN(W2935));
  INVX1 G4009 (.I(W2819), .ZN(W2933));
  INVX1 G4010 (.I(I102), .ZN(W1131));
  INVX1 G4011 (.I(W188), .ZN(W1133));
  INVX1 G4012 (.I(W1076), .ZN(O708));
  INVX1 G4013 (.I(I110), .ZN(W1115));
  INVX1 G4014 (.I(W374), .ZN(W1136));
  INVX1 G4015 (.I(W1706), .ZN(O706));
  INVX1 G4016 (.I(W706), .ZN(W2924));
  INVX1 G4017 (.I(W1564), .ZN(O705));
  INVX1 G4018 (.I(I13), .ZN(W1138));
  INVX1 G4019 (.I(W1130), .ZN(O66));
  INVX1 G4020 (.I(W53), .ZN(W2920));
  INVX1 G4021 (.I(W1616), .ZN(W2913));
  INVX1 G4022 (.I(W1634), .ZN(W2911));
  INVX1 G4023 (.I(W1061), .ZN(O69));
  INVX1 G4024 (.I(W2291), .ZN(O699));
  INVX1 G4025 (.I(W424), .ZN(W1157));
  INVX1 G4026 (.I(W1697), .ZN(W2964));
  INVX1 G4027 (.I(W1326), .ZN(O735));
  INVX1 G4028 (.I(W4), .ZN(O734));
  INVX1 G4029 (.I(W1875), .ZN(O733));
  INVX1 G4030 (.I(I7), .ZN(W2979));
  INVX1 G4031 (.I(W448), .ZN(O732));
  INVX1 G4032 (.I(W1370), .ZN(W2974));
  INVX1 G4033 (.I(W2315), .ZN(O729));
  INVX1 G4034 (.I(W470), .ZN(O728));
  INVX1 G4035 (.I(W1788), .ZN(O727));
  INVX1 G4036 (.I(W968), .ZN(W1092));
  INVX1 G4037 (.I(I76), .ZN(O725));
  INVX1 G4038 (.I(I36), .ZN(W1094));
  INVX1 G4039 (.I(W674), .ZN(W1161));
  INVX1 G4040 (.I(W151), .ZN(W2963));
  INVX1 G4041 (.I(W69), .ZN(W1098));
  INVX1 G4042 (.I(W57), .ZN(W1099));
  INVX1 G4043 (.I(I56), .ZN(W1100));
  INVX1 G4044 (.I(W180), .ZN(W1105));
  INVX1 G4045 (.I(W438), .ZN(W1108));
  INVX1 G4046 (.I(W2900), .ZN(W2952));
  INVX1 G4047 (.I(W2620), .ZN(O717));
  INVX1 G4048 (.I(I34), .ZN(W2950));
  INVX1 G4049 (.I(I138), .ZN(O715));
  INVX1 G4050 (.I(W2826), .ZN(W2947));
  INVX1 G4051 (.I(W2765), .ZN(O660));
  INVX1 G4052 (.I(W2736), .ZN(W2857));
  INVX1 G4053 (.I(W475), .ZN(W1212));
  INVX1 G4054 (.I(W946), .ZN(W1218));
  INVX1 G4055 (.I(W1838), .ZN(O667));
  INVX1 G4056 (.I(W600), .ZN(W1219));
  INVX1 G4057 (.I(W2388), .ZN(W2850));
  INVX1 G4058 (.I(W105), .ZN(O81));
  INVX1 G4059 (.I(W1109), .ZN(W1222));
  INVX1 G4060 (.I(W1880), .ZN(O664));
  INVX1 G4061 (.I(W1048), .ZN(W1225));
  INVX1 G4062 (.I(W1909), .ZN(O662));
  INVX1 G4063 (.I(W1846), .ZN(O661));
  INVX1 G4064 (.I(W833), .ZN(W1210));
  INVX1 G4065 (.I(W1007), .ZN(O659));
  INVX1 G4066 (.I(W239), .ZN(W1227));
  INVX1 G4067 (.I(W901), .ZN(O657));
  INVX1 G4068 (.I(W97), .ZN(W1228));
  INVX1 G4069 (.I(W434), .ZN(W1234));
  INVX1 G4070 (.I(W2551), .ZN(O653));
  INVX1 G4071 (.I(W1618), .ZN(W2832));
  INVX1 G4072 (.I(W481), .ZN(W2830));
  INVX1 G4073 (.I(W266), .ZN(W1240));
  INVX1 G4074 (.I(W1167), .ZN(O85));
  INVX1 G4075 (.I(W2628), .ZN(W2826));
  INVX1 G4076 (.I(W1046), .ZN(O86));
  INVX1 G4077 (.I(W269), .ZN(W1195));
  INVX1 G4078 (.I(W658), .ZN(W1162));
  INVX1 G4079 (.I(I12), .ZN(W1170));
  INVX1 G4080 (.I(W1051), .ZN(W1172));
  INVX1 G4081 (.I(W683), .ZN(W1176));
  INVX1 G4082 (.I(I144), .ZN(W1177));
  INVX1 G4083 (.I(W2344), .ZN(O691));
  INVX1 G4084 (.I(W84), .ZN(W1183));
  INVX1 G4085 (.I(W472), .ZN(W1185));
  INVX1 G4086 (.I(I60), .ZN(O687));
  INVX1 G4087 (.I(W1050), .ZN(W1192));
  INVX1 G4088 (.I(I138), .ZN(O685));
  INVX1 G4089 (.I(W887), .ZN(W2881));
  INVX1 G4090 (.I(W425), .ZN(W801));
  INVX1 G4091 (.I(W1372), .ZN(O682));
  INVX1 G4092 (.I(W2588), .ZN(O681));
  INVX1 G4093 (.I(I29), .ZN(O680));
  INVX1 G4094 (.I(W716), .ZN(O77));
  INVX1 G4095 (.I(W322), .ZN(W2873));
  INVX1 G4096 (.I(W2527), .ZN(O677));
  INVX1 G4097 (.I(W179), .ZN(O676));
  INVX1 G4098 (.I(W1024), .ZN(W1201));
  INVX1 G4099 (.I(W371), .ZN(W1202));
  INVX1 G4100 (.I(W2562), .ZN(W2861));
  INVX1 G4101 (.I(W302), .ZN(W2860));
endmodule
