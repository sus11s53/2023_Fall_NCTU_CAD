module hidden_6 (I0, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I16, I17, I18, I19, I20, I21, I22, I23, I24, I26, I27, I28, I29, I30, I31, I32, I34, I36, I38, I39, I40, I42, I43, I44, I45, I46, I48, I49, I50, I51, I52, I54, I55, I56, I57, I58, I60, I61, I62, I64, I65, I66, I68, I70, I71, I72, I74, I75, I76, I78, I79, I80, I81, I82, I84, I85, I86, I88, I90, I91, I92, I94, I95, I96, I98, I100, I102, I103, I104, I106, I108, I109, I110, I111, I112, I113, I114, I115, I116, I117, I118, I120, I121, I122, I123, I124, I126, I128, I130, I132, I134, I135, I136, I137, I138, I140, I142, I144, I145, I146, I147, I148, I150, I151, I152, I153, I154, I156, I157, I158, I160, I161, I162, I163, I164, I165, I166, I168, I169, I170, I171, I172, I174, I175, I176, I178, I179, I180, I181, I182, I184, I185, I186, I188, I190, I191, I192, I193, I194, I195, I196, I197, I198, I200, I202, I203, I204, I206, I207, I208, I209, I210, I212, I213, I214, I215, I216, I217, I218, I219, I220, I221, I222, I223, I224, I225, I226, I227, I228, I229, I230, I231, I232, I233, I234, I235, I236, I237, I238, I239, I240, I241, I242, I243, I244, I245, I246, I247, I248, I249, I250, I252, I253, I254, I255, I256, I257, I258, I259, I260, I261, I262, I263, I264, I266, I267, I268, I269, I270, I271, I272, I274, I276, I277, I278, I280, I282, I283, I284, I285, I286, I288, I289, I290, I291, I292, I294, I296, I297, I298, I299, I300, I301, I302, I303, I304, I305, I306, I308, I309, I310, I312, I313, I314, I315, I316, I317, I318, I319, I320, I322, I323, I324, I326, I328, I329, I330, I331, I332, I334, I335, I336, I337, I338, I339, I340, I342, I344, I346, I347, I348, I349, I350, I351, I352, I353, I354, I355, I356, I357, I358, I360, I361, I362, I364, I365, I366, I368, I370, I371, I372, I374, I375, I376, I378, I380, I382, I384, I385, I386, I387, I388, I389, I390, I391, I392, I393, I394, I396, I398, I400, I401, I402, I404, I405, I406, I407, I408, I409, I410, I412, I413, I414, I415, I416, I417, I418, I420, I421, I422, I423, I424, I426, I428, I429, I430, I431, I432, I433, I434, I435, I436, I437, I438, I439, I440, I441, I442, I443, I444, I445, I446, I447, I448, I450, I451, I452, I454, I455, I456, I457, I458, I459, I460, I462, I463, I464, I466, I467, I468, I469, I470, I471, I472, I474, I475, I476, I477, I478, I479, I480, I481, I482, I483, I484, I485, I486, I488, I489, I490, I491, I492, I493, I494, I495, I496, I498, I499, I500, I501, I502, I503, I504, I505, I506, I507, I508, I509, I510, I511, I512, I514, I516, I517, I518, I519, I520, I521, I522, I524, I525, I526, I527, I528, I530, I531, I532, I533, I534, I535, I536, I537, I538, I539, I540, I541, I542, I543, I544, I546, I547, I548, I549, I550, I551, I552, I554, I555, I556, I557, I558, I559, I560, I562, I563, I564, I565, I566, I567, I568, I570, I572, I574, I575, I576, I578, I579, I580, I581, I582, I583, I584, I586, I587, I588, I590, I592, I594, I595, I596, I597, I598, I600, I601, I602, I603, I604, I605, I606, I607, I608, I609, I610, I612, I613, I614, I615, I616, I618, I619, I620, I621, I622, I623, I624, I625, I626, I628, I629, I630, I631, I632, I633, I634, I635, I636, I637, I638, I639, I640, I641, I642, I643, I644, I646, I647, I648, I649, I650, I652, I654, I655, I656, I657, I658, I659, I660, I661, I662, I664, I665, I666, I668, I669, I670, I671, I672, I673, I674, I675, I676, I677, I678, I679, I680, I681, I682, I683, I684, I685, I686, I687, I688, I690, I691, I692, I693, I694, I695, I696, I697, I698, I700, I701, I702, I704, I705, I706, I707, I708, I710, I711, I712, I713, I714, I715, I716, I718, I719, I720, I721, I722, I723, I724, I725, I726, I727, I728, I729, I730, I731, I732, I734, I735, I736, I737, I738, I740, I741, I742, I743, I744, I745, I746, I747, I748, I750, I752, I753, I754, I755, I756, I758, I759, I760, I762, I764, I765, I766, I767, I768, I770, I771, I772, I773, I774, I776, I777, I778, I779, I780, I781, I782, I784, I785, I786, I787, I788, I790, I791, I792, I793, I794, I796, I797, I798, I799, I800, I802, I804, I806, I808, I809, I810, I811, I812, I813, I814, I815, I816, I817, I818, I819, I820, I821, I822, I824, I825, I826, I827, I828, I829, I830, I831, I832, I833, I834, I836, I838, I839, I840, I842, I843, I844, I846, I848, I849, I850, I852, I853, I854, I856, I857, I858, I859, I860, I861, I862, I863, I864, I866, I868, I870, I871, I872, I873, I874, I875, I876, I877, I878, I879, I880, I881, I882, I884, I885, I886, I887, I888, I889, I890, I892, I893, I894, I895, I896, I898, I900, I901, I902, I903, I904, I905, I906, I907, I908, I909, I910, I911, I912, I913, I914, I915, I916, I917, I918, I919, I920, I921, I922, I923, I924, I925, I926, I927, I928, I929, I930, I932, I933, I934, I936, I937, I938, I939, I940, I941, I942, I943, I944, I945, I946, I947, I948, I950, I952, I953, I954, I956, I957, I958, I960, I962, I963, I964, I965, I966, I967, I968, I969, I970, I972, I973, I974, I975, I976, I977, I978, I980, I981, I982, I983, I984, I986, I987, I988, I989, I990, I991, I992, I993, I994, I995, I996, I998, I999, I1000, I1001, I1002, I1003, I1004, I1005, I1006, I1008, I1010, I1011, I1012, I1013, I1014, I1015, I1016, I1018, I1019, I1020, I1021, I1022, I1024, I1025, I1026, I1027, I1028, I1029, I1030, I1031, I1032, I1033, I1034, I1036, I1038, I1040, I1041, I1042, I1043, I1044, I1045, I1046, I1047, I1048, I1049, I1050, I1051, I1052, I1053, I1054, I1055, I1056, I1058, I1059, I1060, I1062, I1064, I1065, I1066, I1067, I1068, I1069, I1070, I1072, I1073, I1074, I1075, I1076, I1078, I1079, I1080, I1082, I1084, I1086, I1087, I1088, I1089, I1090, I1091, I1092, I1094, I1095, I1096, I1098, I1100, I1102, I1103, I1104, I1105, I1106, I1107, I1108, I1110, I1111, I1112, I1113, I1114, I1115, I1116, I1117, I1118, I1119, I1120, I1121, I1122, I1123, I1124, I1126, I1127, I1128, I1129, I1130, I1131, I1132, I1133, I1134, I1135, I1136, I1138, I1139, I1140, I1141, I1142, I1143, I1144, I1145, I1146, I1147, I1148, I1149, I1150, I1151, I1152, I1153, I1154, I1156, I1157, I1158, I1159, I1160, I1161, I1162, I1163, I1164, I1165, I1166, I1167, I1168, I1170, I1171, I1172, I1173, I1174, I1175, I1176, I1177, I1178, I1179, I1180, I1181, I1182, I1184, I1186, I1187, I1188, I1189, I1190, I1192, I1193, I1194, I1195, I1196, I1197, I1198, I1199, I1200, I1201, I1202, I1204, I1206, I1208, I1209, I1210, I1211, I1212, I1213, I1214, I1215, I1216, I1217, I1218, I1219, I1220, I1221, I1222, I1224, I1225, I1226, I1228, I1229, I1230, I1231, I1232, I1233, I1234, I1235, I1236, I1238, I1239, I1240, I1242, I1243, I1244, I1245, I1246, I1247, I1248, I1250, I1251, I1252, I1253, I1254, I1255, I1256, I1258, I1259, I1260, I1261, I1262, I1263, I1264, I1265, I1266, I1267, I1268, I1270, I1271, I1272, I1273, I1274, I1276, I1277, I1278, I1280, I1281, I1282, I1283, I1284, I1286, I1287, I1288, I1289, I1290, I1292, I1293, I1294, I1296, I1298, I1299, I1300, I1301, I1302, I1303, I1304, I1305, I1306, I1307, I1308, I1310, I1312, I1314, I1316, I1317, I1318, I1319, I1320, I1321, I1322, I1323, I1324, I1325, I1326, I1328, I1329, I1330, I1331, I1332, I1333, I1334, I1336, I1337, I1338, I1339, I1340, I1341, I1342, I1343, I1344, I1345, I1346, I1347, I1348, I1350, I1352, I1353, I1354, I1355, I1356, I1357, I1358, I1360, I1361, I1362, I1364, I1365, I1366, I1367, I1368, I1370, I1372, I1373, I1374, I1375, I1376, I1377, I1378, I1380, I1381, I1382, I1384, I1385, I1386, I1388, I1389, I1390, I1391, I1392, I1393, I1394, I1395, I1396, I1398, I1399, I1400, I1401, I1402, I1403, I1404, I1406, I1407, I1408, I1409, I1410, I1411, I1412, I1414, I1415, I1416, I1418, I1419, I1420, I1421, I1422, I1423, I1424, I1425, I1426, I1427, I1428, I1429, I1430, I1431, I1432, I1434, I1435, I1436, I1437, I1438, I1439, I1440, I1441, I1442, I1444, I1445, I1446, I1447, I1448, I1449, I1450, I1452, I1453, I1454, I1455, I1456, I1457, I1458, I1459, I1460, I1461, I1462, I1463, I1464, I1465, I1466, I1467, I1468, I1470, I1471, I1472, I1473, I1474, I1475, I1476, I1477, I1478, I1480, I1482, I1483, I1484, I1486, I1488, I1489, I1490, I1491, I1492, I1493, I1494, I1495, I1496, I1497, I1498, I1500, I1501, I1502, I1503, I1504, I1505, I1506, I1507, I1508, I1509, I1510, I1512, I1513, I1514, I1516, I1518, I1519, I1520, I1522, I1523, I1524, I1526, I1528, I1529, I1530, I1531, I1532, I1533, I1534, I1535, I1536, I1538, I1540, I1541, I1542, I1544, I1545, I1546, I1547, I1548, I1550, I1552, I1553, I1554, I1556, I1557, I1558, I1560, I1561, I1562, I1563, I1564, I1565, I1566, I1568, I1569, I1570, I1571, I1572, I1573, I1574, I1575, I1576, I1577, I1578, I1579, I1580, I1582, I1584, I1585, I1586, I1588, I1589, I1590, I1591, I1592, I1593, I1594, I1596, I1597, I1598, I1599, I1600, I1602, I1603, I1604, I1606, I1608, I1609, I1610, I1611, I1612, I1614, I1616, I1617, I1618, I1619, I1620, I1621, I1622, I1624, I1626, I1628, I1629, I1630, I1632, I1633, I1634, I1636, I1637, I1638, I1639, I1640, I1642, I1644, I1646, I1647, I1648, I1649, I1650, I1651, I1652, I1653, I1654, I1656, I1657, I1658, I1659, I1660, I1662, I1663, I1664, I1665, I1666, I1667, I1668, I1669, I1670, I1671, I1672, I1674, I1675, I1676, I1677, I1678, I1679, I1680, I1681, I1682, I1684, I1685, I1686, I1687, I1688, I1689, I1690, I1692, I1694, I1695, I1696, I1697, I1698, I1700, I1701, I1702, I1703, I1704, I1706, I1707, I1708, I1709, I1710, I1711, I1712, I1714, I1715, I1716, I1717, I1718, I1719, I1720, I1722, I1724, I1725, I1726, I1727, I1728, I1729, I1730, I1731, I1732, I1733, I1734, I1736, I1737, I1738, I1739, I1740, I1742, I1743, I1744, I1746, I1747, I1748, I1749, I1750, I1751, I1752, I1753, I1754, I1755, I1756, I1758, I1759, I1760, I1761, I1762, I1763, I1764, I1766, I1768, I1769, I1770, I1772, I1773, I1774, I1775, I1776, I1777, I1778, I1779, I1780, I1782, I1783, I1784, I1786, I1788, I1790, I1792, I1793, I1794, I1795, I1796, I1798, I1799, I1800, I1801, I1802, I1803, I1804, I1806, I1807, I1808, I1809, I1810, I1811, I1812, I1813, I1814, I1815, I1816, I1818, I1819, I1820, I1822, I1824, I1825, I1826, I1828, I1830, I1831, I1832, I1834, I1835, I1836, I1837, I1838, I1839, I1840, I1841, I1842, I1843, I1844, I1846, I1847, I1848, I1850, I1851, I1852, I1853, I1854, I1856, I1858, I1859, I1860, I1861, I1862, I1863, I1864, I1865, I1866, I1868, I1870, I1872, I1873, I1874, I1875, I1876, I1877, I1878, I1880, I1881, I1882, I1883, I1884, I1886, I1887, I1888, I1889, I1890, I1892, I1893, I1894, I1895, I1896, I1898, I1900, I1901, I1902, I1903, I1904, I1906, I1907, I1908, I1909, I1910, I1911, I1912, I1913, I1914, I1915, I1916, I1917, I1918, I1919, I1920, I1921, I1922, I1923, I1924, I1925, I1926, I1927, I1928, I1930, I1931, I1932, I1933, I1934, I1935, I1936, I1937, I1938, I1939, I1940, I1941, I1942, I1943, I1944, I1945, I1946, I1948, I1949, I1950, I1952, I1953, I1954, I1955, I1956, I1957, I1958, I1959, I1960, I1962, I1963, I1964, I1965, I1966, I1968, I1969, I1970, I1972, I1974, I1975, I1976, I1977, I1978, I1979, I1980, I1981, I1982, I1983, I1984, I1985, I1986, I1987, I1988, I1990, I1991, I1992, I1993, I1994, I1996, I1997, I1998, O0, O1, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15, O16, O17, O18, O19, O20, O21, O22, O23, O24, O25, O26, O27, O28, O29, O30, O31, O32, O33, O34, O35, O36, O37, O38, O39, O40, O41, O42, O43, O44, O45, O46, O47, O48, O49, O50, O51, O52, O53, O54, O55, O56, O57, O58, O59, O60, O61, O62, O63, O64, O65, O66, O67, O68, O69, O70, O71, O72, O73, O74, O75, O76, O77, O78, O79, O80, O81, O82, O83, O84, O85, O86, O87, O88, O89, O90, O91, O92, O93, O94, O95, O96, O97, O98, O99, O100, O101, O102, O103, O104, O105, O106, O107, O108, O109, O110, O111, O112, O113, O114, O115, O116, O117, O118, O119, O120, O121, O122, O123, O124, O125, O126, O127, O128, O129, O130, O131, O132, O133, O134, O135, O136, O137, O138, O139, O140, O141, O142, O143, O144, O145, O146, O147, O148, O149, O150, O151, O152, O153, O154, O155, O156, O157, O158, O159, O160, O161, O162, O163, O164, O165, O166, O167, O168, O169, O170, O171, O172, O173, O174, O175, O176, O177, O178, O179, O180, O181, O182, O183, O184, O185, O186, O187, O188, O189, O190, O191, O192, O193, O194, O195, O196, O197, O198, O199, O200, O201, O202, O203, O204, O205, O206, O207, O208, O209, O210, O211, O212, O213, O214, O215, O216, O217, O218, O219, O220, O221, O222, O223, O224, O225, O226, O227, O228, O229, O230, O231, O232, O233, O234, O235, O236, O237, O238, O239, O240, O241, O242, O243, O244, O245, O246, O247, O248, O249, O250, O251, O252, O253, O254, O255, O256, O257, O258, O259, O260, O261, O262, O263, O264, O265, O266, O267, O268, O269, O270, O271, O272, O273, O274, O275, O276, O277, O278, O279, O280, O281, O282, O283, O284, O285, O286, O287, O288, O289, O290, O291, O292, O293, O294, O295, O296, O297, O298, O299, O300, O301, O302, O303, O304, O305, O306, O307, O308, O309, O310, O311, O312, O313, O314, O315, O316, O317, O318, O319, O320, O321, O322, O323, O324, O325, O326, O327, O328, O329, O330, O331, O332, O333, O334, O335, O336, O337, O338, O339, O340, O341, O342, O343, O344, O345, O346, O347, O348, O349, O350, O351, O352, O353, O354, O355, O356, O357, O358, O359, O360, O361, O362, O363, O364, O365, O366, O367, O368, O369, O370, O371, O372, O373, O374, O375, O376, O377, O378, O379, O380, O381, O382, O383, O384, O385, O386, O387, O388, O389, O390, O391, O392, O393, O394, O395, O396, O397, O398, O399, O400, O401, O402, O403, O404, O405, O406, O407, O408, O409, O410, O411, O412, O413, O414, O415, O416, O417, O418, O419, O420, O421, O422, O423, O424, O425, O426, O427, O428, O429, O430, O431, O432, O433, O434, O435, O436, O437, O438, O439, O440, O441, O442, O443, O444, O445, O446, O447, O448, O449, O450, O451, O452, O453, O454, O455, O456, O457, O458, O459, O460, O461, O462, O463, O464, O465, O466, O467, O468, O469, O470, O471, O472, O473, O474, O475, O476, O477, O478, O479, O480, O481, O482, O483, O484, O485, O486, O487, O488, O489, O490, O491, O492, O493, O494, O495, O496, O497, O498, O499, O500, O501, O502, O503, O504, O505, O506, O507, O508, O509, O510, O511, O512, O513, O514, O515, O516, O517, O518, O519, O520, O521, O522, O523, O524, O525, O526, O527, O528, O529, O530, O531, O532, O533, O534, O535, O536, O537, O538, O539, O540, O541, O542, O543, O544, O545, O546, O547, O548, O549, O550, O551, O552, O553, O554, O555, O556, O557, O558, O559, O560, O561, O562, O563, O564, O565, O566, O567, O568, O569, O570, O571, O572, O573, O574, O575, O576, O577, O578, O579, O580, O581, O582, O583, O584, O585, O586, O587, O588, O589, O590, O591, O592, O593, O594, O595, O596, O597, O598, O599, O600, O601, O602, O603, O604, O605, O606, O607, O608, O609, O610, O611, O612, O613, O614, O615, O616, O617, O618, O619, O620, O621, O622, O623, O624, O625, O626, O627, O628, O629, O630, O631, O632, O633, O634, O635, O636, O637, O638, O639, O640, O641, O642, O643, O644, O645, O646, O647, O648, O649, O650, O651, O652, O653, O654, O655, O656, O657, O658, O659, O660, O661, O662, O663, O664, O665, O666, O667, O668, O669, O670, O671, O672, O673, O674, O675, O676, O677, O678, O679, O680, O681, O682, O683, O684, O685, O686, O687, O688, O689, O690, O691, O692, O693, O694, O695, O696, O697, O698, O699, O700, O701, O702, O703, O704, O705, O706, O707, O708, O709, O710, O711, O712, O713, O714, O715, O716, O717, O718, O719, O720, O721, O722, O723, O724, O725, O726, O727, O728, O729, O730, O731, O732, O733, O734, O735, O736, O737, O738, O739, O740, O741, O742, O743, O744, O745, O746, O747, O748, O749, O750, O751, O752, O753, O754, O755, O756, O757, O758, O759, O760, O761, O762, O763, O764, O765, O766, O767, O768, O769, O770, O771, O772, O773, O774, O775, O776, O777, O778, O779, O780, O781, O782, O783, O784, O785, O786, O787, O788, O789, O790, O791, O792, O793, O794, O795, O796, O797, O798, O799, O800, O801, O802, O803, O804, O805, O806, O807, O808, O809, O810, O811, O812, O813, O814, O815, O816, O817, O818, O819, O820, O821, O822, O823, O824, O825, O826, O827, O828, O829, O830, O831, O832, O833, O834, O835, O836, O837, O838, O839, O840, O841, O842, O843, O844, O845, O846, O847, O848, O849, O850, O851, O852, O853, O854, O855, O856, O857, O858, O859, O860, O861, O862, O863, O864, O865, O866, O867, O868, O869, O870, O871, O872, O873, O874, O875, O876, O877, O878, O879, O880, O881, O882, O883, O884, O885, O886, O887, O888, O889, O890, O891, O892, O893, O894, O895, O896, O897, O898, O899, O900, O901, O902, O903, O904, O905, O906, O907, O908, O909, O910, O911, O912, O913, O914, O915, O916, O917, O918, O919, O920, O921, O922, O923, O924, O925, O926, O927, O928, O929, O930, O931, O932, O933, O934, O935, O936, O937, O938, O939, O940, O941, O942, O943, O944, O945, O946, O947, O948, O949, O950, O951, O952, O953, O954, O955, O956, O957, O958, O959, O960, O961, O962, O963, O964, O965, O966, O967, O968, O969, O970, O971, O972, O973, O974, O975, O976, O977, O978, O979, O980, O981, O982, O983, O984, O985, O986, O987, O988, O989, O990, O991, O992, O993, O994, O995, O996, O997, O998, O999, O1000, O1001, O1002, O1003, O1004, O1005, O1006, O1007, O1008, O1009, O1010, O1011, O1012, O1013, O1014, O1015, O1016, O1017, O1018, O1019, O1020, O1021, O1022, O1023, O1024, O1025, O1026, O1027, O1028, O1029, O1030, O1031, O1032, O1033, O1034, O1035, O1036, O1037, O1038, O1039, O1040, O1041, O1042, O1043, O1044, O1045, O1046, O1047, O1048, O1049, O1050, O1051, O1052, O1053, O1054, O1055, O1056, O1057, O1058, O1059, O1060, O1061, O1062, O1063, O1064, O1065, O1066, O1067, O1068, O1069, O1070, O1071, O1072, O1073, O1074, O1075, O1076, O1077, O1078, O1079, O1080, O1081, O1082, O1083, O1084, O1085, O1086, O1087, O1088, O1089, O1090, O1091, O1092, O1093, O1094, O1095, O1096, O1097, O1098, O1099, O1100, O1101, O1102, O1103, O1104, O1105, O1106, O1107, O1108, O1109, O1110, O1111, O1112, O1113, O1114, O1115, O1116, O1117, O1118, O1119, O1120, O1121, O1122, O1123, O1124, O1125, O1126, O1127, O1128, O1129, O1130, O1131, O1132, O1133, O1134, O1135, O1136, O1137, O1138, O1139, O1140, O1141, O1142, O1143, O1144, O1145, O1146, O1147, O1148, O1149, O1150, O1151, O1152, O1153, O1154, O1155, O1156, O1157, O1158, O1159, O1160, O1161, O1162, O1163, O1164, O1165, O1166, O1167, O1168, O1169, O1170, O1171, O1172, O1173, O1174, O1175, O1176, O1177, O1178, O1179, O1180, O1181, O1182, O1183, O1184, O1185, O1186, O1187, O1188, O1189, O1190, O1191, O1192, O1193, O1194, O1195, O1196, O1197, O1198, O1199, O1200, O1201, O1202, O1203, O1204, O1205, O1206, O1207, O1208, O1209, O1210, O1211, O1212, O1213, O1214, O1215, O1216, O1217, O1218, O1219, O1220, O1221, O1222, O1223, O1224, O1225, O1226, O1227, O1228, O1229, O1230, O1231, O1232, O1233, O1234, O1235, O1236, O1237, O1238, O1239, O1240, O1241, O1242, O1243, O1244, O1245, O1246, O1247, O1248, O1249, O1250, O1251, O1252, O1253, O1254, O1255, O1256, O1257, O1258, O1259, O1260, O1261, O1262, O1263, O1264, O1265, O1266, O1267, O1268, O1269, O1270, O1271, O1272, O1273, O1274, O1275, O1276, O1277, O1278, O1279, O1280, O1281, O1282, O1283, O1284, O1285, O1286, O1287, O1288, O1289, O1290, O1291, O1292, O1293, O1294, O1295, O1296, O1297, O1298, O1299, O1300, O1301, O1302, O1303, O1304, O1305, O1306, O1307, O1308, O1309, O1310, O1311, O1312, O1313, O1314, O1315, O1316, O1317, O1318, O1319, O1320, O1321, O1322, O1323, O1324, O1325, O1326, O1327, O1328, O1329, O1330, O1331, O1332, O1333, O1334, O1335, O1336, O1337, O1338, O1339, O1340, O1341, O1342, O1343, O1344, O1345, O1346, O1347, O1348, O1349, O1350, O1351, O1352, O1353, O1354, O1355, O1356, O1357, O1358, O1359, O1360, O1361, O1362, O1363, O1364, O1365, O1366, O1367, O1368, O1369, O1370, O1371, O1372, O1373, O1374, O1375, O1376, O1377, O1378, O1379, O1380, O1381, O1382, O1383, O1384, O1385, O1386, O1387, O1388, O1389, O1390, O1391, O1392, O1393, O1394, O1395, O1396, O1397, O1398, O1399, O1400, O1401, O1402, O1403, O1404, O1405, O1406, O1407, O1408, O1409, O1410, O1411, O1412, O1413, O1414, O1415, O1416, O1417, O1418, O1419, O1420, O1421, O1422, O1423, O1424, O1425, O1426, O1427, O1428, O1429, O1430, O1431, O1432, O1433, O1434, O1435, O1436, O1437, O1438, O1439, O1440, O1441, O1442, O1443, O1444, O1445, O1446, O1447, O1448, O1449, O1450, O1451, O1452, O1453, O1454, O1455, O1456, O1457, O1458, O1459, O1460, O1461, O1462, O1463, O1464, O1465, O1466, O1467, O1468, O1469, O1470, O1471, O1472, O1473, O1474, O1475, O1476, O1477, O1478, O1479, O1480, O1481, O1482, O1483, O1484, O1485, O1486, O1487, O1488, O1489, O1490, O1491, O1492, O1493, O1494, O1495, O1496, O1497, O1498, O1499, O1500, O1501, O1502, O1503, O1504, O1505, O1506, O1507, O1508, O1509, O1510, O1511, O1512, O1513, O1514, O1515, O1516, O1517, O1518, O1519, O1520, O1521, O1522, O1523, O1524, O1525, O1526, O1527, O1528, O1529, O1530, O1531, O1532, O1533, O1534, O1535, O1536, O1537, O1538, O1539, O1540, O1541, O1542, O1543, O1544, O1545, O1546, O1547, O1548, O1549, O1550, O1551, O1552, O1553, O1554, O1555, O1556, O1557, O1558, O1559, O1560, O1561, O1562, O1563, O1564, O1565, O1566, O1567, O1568, O1569, O1570, O1571, O1572, O1573, O1574, O1575, O1576, O1577, O1578, O1579, O1580, O1581, O1582, O1583, O1584, O1585, O1586, O1587, O1588, O1589, O1590, O1591, O1592, O1593, O1594, O1595, O1596, O1597, O1598, O1599, O1600, O1601, O1602, O1603, O1604, O1605, O1606, O1607, O1608, O1609, O1610, O1611, O1612, O1613, O1614, O1615, O1616, O1617, O1618, O1619, O1620, O1621, O1622, O1623, O1624, O1625, O1626, O1627, O1628, O1629, O1630, O1631, O1632, O1633, O1634, O1635, O1636, O1637, O1638, O1639, O1640, O1641, O1642, O1643, O1644, O1645, O1646, O1647, O1648, O1649, O1650, O1651, O1652, O1653, O1654, O1655, O1656, O1657, O1658, O1659, O1660, O1661, O1662, O1663, O1664, O1665, O1666, O1667, O1668, O1669, O1670, O1671, O1672, O1673, O1674, O1675, O1676, O1677, O1678, O1679, O1680, O1681, O1682, O1683, O1684, O1685, O1686, O1687, O1688, O1689, O1690, O1691, O1692, O1693, O1694, O1695, O1696, O1697, O1698, O1699, O1700, O1701, O1702, O1703, O1704, O1705, O1706, O1707, O1708, O1709, O1710, O1711, O1712, O1713, O1714, O1715, O1716, O1717, O1718, O1719, O1720, O1721, O1722, O1723, O1724, O1725, O1726, O1727, O1728, O1729, O1730, O1731, O1732, O1733, O1734, O1735, O1736, O1737, O1738, O1739, O1740, O1741, O1742, O1743, O1744, O1745, O1746, O1747, O1748, O1749, O1750, O1751, O1752, O1753, O1754, O1755, O1756, O1757, O1758, O1759, O1760, O1761, O1762, O1763, O1764, O1765, O1766, O1767, O1768, O1769, O1770, O1771, O1772, O1773, O1774, O1775, O1776, O1777, O1778, O1779, O1780, O1781, O1782, O1783, O1784, O1785, O1786, O1787, O1788, O1789, O1790, O1791, O1792, O1793, O1794, O1795, O1796, O1797, O1798, O1799, O1800, O1801, O1802, O1803, O1804, O1805, O1806, O1807, O1808, O1809, O1810, O1811, O1812, O1813, O1814, O1815, O1816, O1817, O1818, O1819, O1820, O1821, O1822, O1823, O1824, O1825, O1826, O1827, O1828, O1829, O1830, O1831, O1832, O1833, O1834, O1835, O1836, O1837, O1838, O1839, O1840, O1841, O1842, O1843, O1844, O1845, O1846, O1847, O1848, O1849, O1850, O1851, O1852, O1853, O1854, O1855, O1856, O1857, O1858, O1859, O1860, O1861, O1862, O1863, O1864, O1865, O1866, O1867, O1868, O1869, O1870, O1871, O1872, O1873, O1874, O1875, O1876, O1877, O1878, O1879, O1880, O1881, O1882, O1883, O1884, O1885, O1886, O1887, O1888, O1889, O1890, O1891, O1892, O1893, O1894, O1895, O1896, O1897, O1898, O1899, O1900, O1901, O1902, O1903, O1904, O1905, O1906, O1907, O1908, O1909, O1910, O1911, O1912, O1913, O1914, O1915, O1916, O1917, O1918, O1919, O1920, O1921, O1922, O1923, O1924, O1925, O1926, O1927, O1928, O1929, O1930, O1931, O1932, O1933, O1934, O1935, O1936, O1937, O1938, O1939, O1940, O1941, O1942, O1943, O1944, O1945, O1946, O1947, O1948, O1949, O1950, O1951, O1952, O1953, O1954, O1955, O1956, O1957, O1958, O1959, O1960, O1961, O1962, O1963, O1964, O1965, O1966, O1967, O1968, O1969, O1970, O1971, O1972, O1973, O1974, O1975, O1976, O1977, O1978, O1979, O1980, O1981, O1982, O1983, O1984, O1985, O1986, O1987, O1988, O1989, O1990, O1991, O1992, O1993, O1994, O1995, O1996, O1997, O1998, O1999, O2000, O2001, O2002, O2003, O2004, O2005, O2006, O2007, O2008, O2009, O2010, O2011, O2012, O2013, O2014, O2015, O2016, O2017, O2018, O2019, O2020, O2021, O2022, O2023, O2024, O2025, O2026, O2027, O2028, O2029, O2030, O2031, O2032, O2033, O2034, O2035, O2036, O2037, O2038, O2039, O2040, O2041, O2042, O2043, O2044, O2045, O2046, O2047, O2048, O2049, O2050, O2051, O2052, O2053, O2054, O2055, O2056, O2057, O2058, O2059, O2060, O2061, O2062, O2063, O2064, O2065, O2066, O2067, O2068, O2069, O2070, O2071, O2072, O2073, O2074, O2075, O2076, O2077, O2078, O2079, O2080, O2081, O2082, O2083, O2084, O2085, O2086, O2087, O2088, O2089, O2090, O2091, O2092, O2093, O2094, O2095, O2096, O2097, O2098, O2099, O2100, O2101, O2102, O2103, O2104, O2105, O2106, O2107, O2108, O2109, O2110, O2111, O2112, O2113, O2114, O2115, O2116, O2117, O2118, O2119, O2120, O2121, O2122, O2123, O2124, O2125, O2126, O2127, O2128, O2129, O2130, O2131, O2132, O2133, O2134, O2135, O2136, O2137, O2138, O2139, O2140, O2141, O2142, O2143, O2144, O2145, O2146, O2147, O2148, O2149, O2150, O2151, O2152, O2153, O2154, O2155, O2156, O2157, O2158, O2159, O2160, O2161, O2162, O2163, O2164, O2165, O2166, O2167, O2168, O2169, O2170, O2171, O2172, O2173, O2174, O2175, O2176, O2177, O2178, O2179, O2180, O2181, O2182, O2183, O2184, O2185, O2186, O2187, O2188, O2189, O2190, O2191, O2192, O2193, O2194, O2195, O2196, O2197, O2198, O2199, O2200, O2201, O2202, O2203, O2204, O2205, O2206, O2207, O2208, O2209, O2210, O2211, O2212, O2213, O2214, O2215, O2216, O2217, O2218, O2219, O2220, O2221, O2222, O2223, O2224, O2225, O2226, O2227, O2228, O2229, O2230, O2231, O2232, O2233, O2234, O2235, O2236, O2237, O2238, O2239, O2240, O2241, O2242, O2243, O2244, O2245, O2246, O2247, O2248, O2249, O2250, O2251, O2252, O2253, O2254, O2255, O2256, O2257, O2258, O2259, O2260, O2261, O2262, O2263, O2264, O2265, O2266, O2267, O2268, O2269, O2270, O2271, O2272, O2273, O2274, O2275, O2276, O2277, O2278, O2279, O2280, O2281, O2282, O2283, O2284, O2285, O2286, O2287, O2288, O2289, O2290, O2291, O2292, O2293, O2294, O2295, O2296, O2297, O2298, O2299, O2300, O2301, O2302, O2303, O2304, O2305, O2306, O2307, O2308, O2309, O2310, O2311, O2312, O2313, O2314, O2315, O2316, O2317, O2318, O2319, O2320, O2321, O2322, O2323, O2324, O2325, O2326, O2327, O2328, O2329, O2330, O2331, O2332, O2333, O2334, O2335, O2336, O2337, O2338, O2339, O2340, O2341, O2342, O2343, O2344, O2345, O2346, O2347, O2348, O2349, O2350, O2351, O2352, O2353, O2354, O2355, O2356, O2357, O2358, O2359, O2360, O2361, O2362, O2363, O2364, O2365, O2366, O2367, O2368, O2369, O2370, O2371, O2372, O2373, O2374, O2375, O2376, O2377, O2378, O2379, O2380, O2381, O2382, O2383, O2384, O2385, O2386, O2387, O2388, O2389, O2390, O2391, O2392, O2393, O2394, O2395, O2396, O2397, O2398, O2399, O2400, O2401, O2402, O2403, O2404, O2405, O2406, O2407, O2408, O2409, O2410, O2411, O2412, O2413, O2414, O2415, O2416, O2417, O2418, O2419, O2420, O2421, O2422, O2423, O2424, O2425, O2426, O2427, O2428, O2429, O2430, O2431, O2432, O2433, O2434, O2435, O2436, O2437, O2438, O2439, O2440, O2441, O2442, O2443, O2444, O2445, O2446, O2447, O2448, O2449, O2450, O2451, O2452, O2453, O2454, O2455, O2456, O2457, O2458, O2459, O2460, O2461, O2462, O2463, O2464, O2465, O2466, O2467, O2468, O2469, O2470, O2471, O2472, O2473, O2474, O2475, O2476, O2477, O2478, O2479, O2480, O2481, O2482, O2483, O2484, O2485, O2486, O2487, O2488, O2489, O2490, O2491, O2492, O2493, O2494, O2495, O2496, O2497, O2498, O2499, O2500, O2501, O2502, O2503, O2504, O2505, O2506, O2507, O2508, O2509, O2510, O2511, O2512, O2513, O2514, O2515, O2516, O2517, O2518, O2519, O2520, O2521, O2522, O2523, O2524, O2525, O2526, O2527, O2528, O2529, O2530, O2531, O2532, O2533, O2534, O2535, O2536, O2537, O2538, O2539, O2540, O2541, O2542, O2543, O2544, O2545, O2546, O2547, O2548, O2549, O2550, O2551, O2552, O2553, O2554, O2555, O2556, O2557, O2558, O2559, O2560, O2561, O2562, O2563, O2564, O2565, O2566, O2567, O2568, O2569, O2570, O2571, O2572, O2573, O2574, O2575, O2576, O2577, O2578, O2579, O2580, O2581, O2582, O2583, O2584, O2585, O2586, O2587, O2588, O2589, O2590, O2591, O2592, O2593, O2594, O2595, O2596, O2597, O2598, O2599, O2600, O2601, O2602, O2603, O2604, O2605, O2606, O2607, O2608, O2609, O2610, O2611, O2612, O2613, O2614, O2615, O2616, O2617, O2618, O2619, O2620, O2621, O2622, O2623, O2624, O2625, O2626, O2627, O2628, O2629, O2630, O2631, O2632, O2633, O2634, O2635, O2636, O2637, O2638, O2639, O2640, O2641, O2642, O2643, O2644, O2645, O2646, O2647, O2648, O2649, O2650, O2651, O2652, O2653, O2654, O2655, O2656, O2657, O2658, O2659, O2660, O2661, O2662, O2663, O2664, O2665, O2666, O2667, O2668, O2669, O2670, O2671, O2672, O2673, O2674, O2675, O2676, O2677, O2678, O2679, O2680, O2681, O2682, O2683, O2684, O2685, O2686, O2687, O2688, O2689, O2690, O2691, O2692, O2693, O2694, O2695, O2696, O2697, O2698, O2699, O2700, O2701, O2702, O2703, O2704, O2705, O2706, O2707, O2708, O2709, O2710, O2711, O2712, O2713, O2714, O2715, O2716, O2717, O2718, O2719, O2720, O2721, O2722, O2723, O2724, O2725, O2726, O2727, O2728, O2729, O2730, O2731, O2732, O2733, O2734, O2735, O2736, O2737, O2738, O2739, O2740, O2741, O2742, O2743, O2744, O2745, O2746, O2747, O2748, O2749, O2750, O2751, O2752, O2753, O2754, O2755, O2756, O2757, O2758, O2759, O2760, O2761, O2762, O2763, O2764, O2765, O2766, O2767, O2768, O2769, O2770, O2771, O2772, O2773, O2774, O2775, O2776, O2777, O2778, O2779, O2780, O2781, O2782, O2783, O2784, O2785, O2786, O2787, O2788, O2789, O2790, O2791, O2792, O2793, O2794, O2795, O2796, O2797, O2798, O2799, O2800, O2801, O2802, O2803, O2804, O2805, O2806, O2807, O2808, O2809, O2810, O2811, O2812, O2813, O2814, O2815, O2816, O2817, O2818, O2819, O2820, O2821, O2822, O2823, O2824, O2825, O2826, O2827, O2828, O2829, O2830, O2831, O2832, O2833, O2834, O2835, O2836, O2837, O2838, O2839, O2840, O2841, O2842, O2843, O2844, O2845, O2846, O2847, O2848, O2849, O2850, O2851, O2852, O2853, O2854, O2855, O2856, O2857, O2858, O2859, O2860, O2861, O2862, O2863, O2864, O2865, O2866, O2867, O2868, O2869, O2870, O2871, O2872, O2873, O2874, O2875, O2876, O2877, O2878, O2879, O2880, O2881, O2882, O2883, O2884, O2885, O2886, O2887, O2888, O2889, O2890, O2891, O2892, O2893, O2894, O2895, O2896, O2897, O2898, O2899, O2900, O2901, O2902, O2903, O2904, O2905, O2906, O2907, O2908, O2909, O2910, O2911, O2912, O2913, O2914, O2915, O2916, O2917, O2918, O2919, O2920, O2921, O2922, O2923, O2924, O2925, O2926, O2927, O2928, O2929, O2930, O2931, O2932, O2933, O2934, O2935, O2936, O2937, O2938, O2939, O2940, O2941, O2942, O2943, O2944, O2945, O2946, O2947, O2948, O2949, O2950, O2951, O2952, O2953, O2954, O2955, O2956, O2957, O2958, O2959, O2960, O2961, O2962, O2963, O2964, O2965, O2966, O2967, O2968, O2969, O2970, O2971, O2972, O2973, O2974, O2975, O2976, O2977, O2978, O2979, O2980, O2981, O2982, O2983, O2984, O2985, O2986, O2987, O2988, O2989, O2990, O2991, O2992, O2993, O2994, O2995, O2996, O2997, O2998, O2999, O3000, O3001, O3002, O3003, O3004, O3005, O3006, O3007, O3008, O3009, O3010, O3011, O3012, O3013, O3014, O3015, O3016, O3017, O3018, O3019, O3020, O3021, O3022, O3023, O3024, O3025, O3026, O3027, O3028, O3029, O3030, O3031, O3032, O3033, O3034, O3035, O3036, O3037, O3038, O3039, O3040, O3041, O3042, O3043, O3044, O3045, O3046, O3047, O3048, O3049, O3050, O3051, O3052, O3053, O3054, O3055, O3056, O3057, O3058, O3059, O3060, O3061, O3062, O3063, O3064, O3065, O3066, O3067, O3068, O3069, O3070, O3071, O3072, O3073, O3074, O3075, O3076, O3077, O3078, O3079, O3080, O3081, O3082, O3083, O3084, O3085, O3086, O3087, O3088, O3089, O3090, O3091, O3092, O3093, O3094, O3095, O3096, O3097, O3098, O3099, O3100, O3101, O3102, O3103, O3104, O3105, O3106, O3107, O3108, O3109, O3110, O3111, O3112, O3113, O3114, O3115, O3116, O3117, O3118, O3119, O3120, O3121, O3122, O3123, O3124, O3125, O3126, O3127, O3128, O3129, O3130, O3131, O3132, O3133, O3134, O3135, O3136, O3137, O3138, O3139, O3140, O3141, O3142, O3143, O3144, O3145, O3146, O3147, O3148, O3149, O3150, O3151, O3152, O3153, O3154, O3155, O3156, O3157, O3158, O3159, O3160, O3161, O3162, O3163, O3164, O3165, O3166, O3167, O3168, O3169, O3170, O3171, O3172, O3173, O3174, O3175, O3176, O3177, O3178, O3179, O3180, O3181, O3182, O3183, O3184, O3185, O3186, O3187, O3188, O3189, O3190, O3191, O3192, O3193, O3194, O3195, O3196, O3197, O3198, O3199, O3200, O3201, O3202, O3203, O3204, O3205, O3206, O3207, O3208, O3209, O3210, O3211, O3212, O3213, O3214, O3215, O3216, O3217, O3218, O3219, O3220, O3221, O3222, O3223, O3224, O3225, O3226, O3227, O3228, O3229, O3230, O3231, O3232, O3233, O3234, O3235, O3236, O3237, O3238, O3239, O3240, O3241, O3242, O3243, O3244, O3245, O3246, O3247, O3248, O3249, O3250, O3251, O3252, O3253, O3254, O3255, O3256, O3257, O3258, O3259, O3260, O3261, O3262, O3263, O3264, O3265, O3266, O3267, O3268, O3269, O3270, O3271, O3272, O3273, O3274, O3275, O3276, O3277, O3278, O3279, O3280, O3281, O3282, O3283, O3284, O3285, O3286, O3287, O3288, O3289, O3290, O3291, O3292, O3293, O3294, O3295, O3296, O3297, O3298, O3299, O3300, O3301, O3302, O3303, O3304, O3305, O3306, O3307, O3308, O3309, O3310, O3311, O3312, O3313, O3314, O3315, O3316, O3317, O3318, O3319, O3320, O3321, O3322, O3323, O3324, O3325, O3326, O3327, O3328, O3329, O3330, O3331, O3332, O3333, O3334, O3335, O3336, O3337, O3338, O3339, O3340, O3341, O3342, O3343, O3344, O3345, O3346, O3347, O3348, O3349, O3350, O3351, O3352, O3353, O3354, O3355, O3356, O3357, O3358, O3359, O3360, O3361, O3362, O3363, O3364, O3365, O3366, O3367, O3368, O3369, O3370, O3371, O3372, O3373, O3374, O3375, O3376, O3377, O3378, O3379, O3380, O3381, O3382, O3383, O3384, O3385, O3386, O3387, O3388, O3389, O3390, O3391, O3392, O3393, O3394, O3395, O3396, O3397, O3398, O3399, O3400, O3401, O3402, O3403, O3404, O3405, O3406, O3407, O3408, O3409, O3410, O3411, O3412, O3413, O3414, O3415, O3416, O3417, O3418, O3419, O3420, O3421, O3422, O3423, O3424, O3425, O3426, O3427, O3428, O3429, O3430, O3431, O3432, O3433, O3434, O3435, O3436, O3437, O3438, O3439, O3440, O3441, O3442, O3443, O3444, O3445, O3446, O3447, O3448, O3449, O3450, O3451, O3452, O3453, O3454, O3455, O3456, O3457, O3458, O3459, O3460, O3461, O3462, O3463, O3464, O3465, O3466, O3467, O3468, O3469, O3470, O3471, O3472, O3473, O3474, O3475, O3476, O3477, O3478, O3479, O3480, O3481, O3482, O3483, O3484, O3485, O3486, O3487, O3488, O3489, O3490, O3491, O3492, O3493, O3494, O3495, O3496, O3497, O3498, O3499, O3500, O3501, O3502, O3503, O3504, O3505, O3506, O3507, O3508, O3509, O3510, O3511, O3512, O3513, O3514, O3515, O3516, O3517, O3518, O3519, O3520, O3521, O3522, O3523, O3524, O3525, O3526, O3527, O3528, O3529, O3530, O3531, O3532, O3533, O3534, O3535, O3536, O3537, O3538, O3539, O3540, O3541, O3542, O3543, O3544, O3545, O3546, O3547, O3548, O3549, O3550, O3551, O3552, O3553, O3554, O3555, O3556, O3557, O3558, O3559, O3560, O3561, O3562, O3563, O3564, O3565, O3566, O3567, O3568, O3569, O3570, O3571, O3572, O3573, O3574, O3575, O3576, O3577, O3578, O3579, O3580, O3581, O3582, O3583, O3584, O3585, O3586, O3587, O3588, O3589, O3590, O3591, O3592, O3593, O3594, O3595, O3596, O3597, O3598, O3599, O3600, O3601, O3602, O3603, O3604, O3605, O3606, O3607, O3608, O3609, O3610, O3611, O3612, O3613, O3614, O3615, O3616, O3617, O3618, O3619, O3620, O3621, O3622, O3623, O3624, O3625, O3626, O3627, O3628, O3629, O3630, O3631, O3632, O3633, O3634, O3635, O3636, O3637, O3638, O3639, O3640, O3641, O3642, O3643, O3644, O3645, O3646, O3647, O3648, O3649, O3650, O3651, O3652, O3653, O3654, O3655, O3656, O3657, O3658, O3659, O3660, O3661, O3662, O3663, O3664, O3665, O3666, O3667, O3668, O3669, O3670, O3671, O3672, O3673, O3674, O3675, O3676, O3677, O3678, O3679, O3680, O3681, O3682, O3683, O3684, O3685, O3686, O3687, O3688, O3689, O3690, O3691, O3692, O3693, O3694, O3695, O3696, O3697, O3698, O3699, O3700, O3701, O3702, O3703, O3704, O3705, O3706, O3707, O3708, O3709, O3710, O3711, O3712, O3713, O3714, O3715, O3716, O3717, O3718, O3719, O3720, O3721, O3722, O3723, O3724, O3725, O3726, O3727, O3728, O3729, O3730, O3731, O3732, O3733, O3734, O3735, O3736, O3737, O3738, O3739, O3740, O3741, O3742, O3743, O3744, O3745, O3746, O3747, O3748, O3749, O3750, O3751, O3752, O3753, O3754, O3755, O3756, O3757, O3758, O3759, O3760, O3761, O3762, O3763, O3764, O3765, O3766, O3767, O3768, O3769, O3770, O3771, O3772, O3773, O3774, O3775, O3776, O3777, O3778, O3779, O3780, O3781, O3782, O3783, O3784, O3785, O3786, O3787, O3788, O3789, O3790, O3791, O3792, O3793, O3794, O3795, O3796, O3797, O3798, O3799, O3800, O3801, O3802, O3803, O3804, O3805, O3806, O3807, O3808, O3809, O3810, O3811, O3812, O3813, O3814, O3815, O3816, O3817, O3818, O3819, O3820, O3821, O3822, O3823, O3824, O3825, O3826, O3827, O3828, O3829, O3830, O3831, O3832, O3833, O3834, O3835, O3836, O3837, O3838, O3839, O3840, O3841, O3842, O3843, O3844, O3845, O3846, O3847, O3848, O3849, O3850, O3851, O3852, O3853, O3854, O3855, O3856, O3857, O3858, O3859, O3860, O3861, O3862, O3863, O3864, O3865, O3866, O3867, O3868, O3869, O3870, O3871, O3872, O3873, O3874, O3875, O3876, O3877, O3878, O3879, O3880, O3881, O3882, O3883, O3884, O3885, O3886, O3887, O3888, O3889, O3890, O3891, O3892, O3893, O3894, O3895, O3896, O3897, O3898, O3899, O3900, O3901, O3902, O3903, O3904, O3905, O3906, O3907, O3908, O3909, O3910, O3911, O3912, O3913, O3914, O3915, O3916, O3917, O3918, O3919, O3920, O3921, O3922, O3923, O3924, O3925, O3926, O3927, O3928, O3929, O3930, O3931, O3932, O3933, O3934, O3935, O3936, O3937, O3938, O3939, O3940, O3941, O3942, O3943, O3944, O3945, O3946, O3947, O3948, O3949, O3950, O3951, O3952, O3953, O3954, O3955, O3956, O3957, O3958, O3959, O3960, O3961, O3962, O3963, O3964, O3965, O3966, O3967, O3968, O3969, O3970, O3971, O3972, O3973, O3974, O3975, O3976, O3977, O3978, O3979, O3980, O3981, O3982, O3983, O3984, O3985, O3986, O3987, O3988, O3989, O3990, O3991, O3992, O3993, O3994, O3995, O3996, O3997, O3998, O3999, O4000, O4001, O4002, O4003, O4004, O4005, O4006, O4007, O4008, O4009, O4010, O4011, O4012, O4013, O4014, O4015, O4016, O4017, O4018, O4019, O4020, O4021, O4022, O4023, O4024, O4025, O4026, O4027, O4028, O4029, O4030, O4031, O4032, O4033, O4034, O4035, O4036, O4037, O4038, O4039, O4040, O4041, O4042, O4043, O4044, O4045, O4046, O4047, O4048, O4049, O4050, O4051, O4052, O4053, O4054, O4055, O4056, O4057, O4058, O4059, O4060, O4061, O4062, O4063, O4064, O4065, O4066, O4067, O4068, O4069, O4070, O4071, O4072, O4073, O4074, O4075, O4076, O4077, O4078, O4079, O4080, O4081, O4082, O4083, O4084, O4085, O4086, O4087, O4088, O4089, O4090, O4091, O4092, O4093, O4094, O4095, O4096, O4097, O4098, O4099, O4100, O4101, O4102, O4103, O4104, O4105, O4106, O4107, O4108, O4109, O4110, O4111, O4112, O4113, O4114, O4115, O4116, O4117, O4118, O4119, O4120, O4121, O4122, O4123, O4124, O4125, O4126, O4127, O4128, O4129, O4130, O4131, O4132, O4133, O4134, O4135, O4136, O4137, O4138, O4139, O4140, O4141, O4142, O4143, O4144, O4145, O4146, O4147, O4148, O4149, O4150, O4151, O4152, O4153, O4154, O4155, O4156, O4157, O4158, O4159, O4160, O4161, O4162, O4163, O4164, O4165, O4166, O4167, O4168, O4169, O4170, O4171, O4172, O4173, O4174, O4175, O4176, O4177, O4178, O4179, O4180, O4181, O4182, O4183, O4184, O4185, O4186, O4187, O4188, O4189, O4190, O4191, O4192, O4193, O4194, O4195, O4196, O4197, O4198, O4199, O4200, O4201, O4202, O4203, O4204, O4205, O4206, O4207, O4208, O4209, O4210, O4211, O4212, O4213, O4214, O4215, O4216, O4217, O4218, O4219, O4220, O4221, O4222, O4223, O4224, O4225, O4226, O4227, O4228, O4229, O4230, O4231, O4232, O4233, O4234, O4235, O4236, O4237, O4238, O4239, O4240, O4241, O4242, O4243, O4244, O4245, O4246, O4247, O4248, O4249, O4250, O4251, O4252, O4253, O4254, O4255, O4256, O4257, O4258, O4259, O4260, O4261, O4262, O4263, O4264, O4265, O4266, O4267, O4268, O4269, O4270, O4271, O4272, O4273, O4274, O4275, O4276, O4277, O4278, O4279, O4280, O4281, O4282, O4283, O4284, O4285, O4286, O4287, O4288, O4289, O4290, O4291, O4292, O4293, O4294, O4295, O4296, O4297, O4298, O4299, O4300, O4301, O4302, O4303, O4304, O4305, O4306, O4307, O4308, O4309, O4310, O4311, O4312, O4313, O4314, O4315, O4316, O4317, O4318, O4319, O4320, O4321, O4322, O4323, O4324, O4325, O4326, O4327, O4328, O4329, O4330, O4331, O4332, O4333, O4334, O4335, O4336, O4337, O4338, O4339, O4340, O4341, O4342, O4343, O4344, O4345, O4346, O4347, O4348, O4349, O4350, O4351, O4352, O4353, O4354, O4355, O4356, O4357, O4358, O4359, O4360, O4361, O4362, O4363, O4364, O4365, O4366, O4367, O4368, O4369, O4370, O4371, O4372, O4373, O4374, O4375, O4376, O4377, O4378, O4379, O4380, O4381, O4382, O4383, O4384, O4385, O4386, O4387, O4388, O4389, O4390, O4391, O4392, O4393, O4394, O4395, O4396, O4397, O4398, O4399, O4400, O4401, O4402, O4403, O4404, O4405, O4406, O4407, O4408, O4409, O4410, O4411, O4412, O4413, O4414, O4415, O4416, O4417, O4418, O4419, O4420, O4421, O4422, O4423, O4424, O4425, O4426, O4427, O4428, O4429, O4430, O4431, O4432, O4433, O4434, O4435, O4436, O4437, O4438, O4439, O4440, O4441, O4442, O4443, O4444, O4445, O4446, O4447, O4448, O4449, O4450, O4451, O4452, O4453, O4454, O4455, O4456, O4457, O4458, O4459, O4460, O4461, O4462, O4463, O4464, O4465, O4466, O4467, O4468, O4469, O4470, O4471, O4472, O4473, O4474, O4475, O4476, O4477, O4478, O4479, O4480, O4481, O4482, O4483, O4484, O4485, O4486, O4487, O4488, O4489, O4490, O4491, O4492, O4493, O4494, O4495, O4496, O4497, O4498, O4499, O4500, O4501, O4502, O4503, O4504, O4505, O4506, O4507, O4508, O4509, O4510, O4511, O4512, O4513, O4514, O4515, O4516, O4517, O4518, O4519, O4520, O4521, O4522, O4523, O4524, O4525, O4526, O4527, O4528, O4529, O4530, O4531, O4532, O4533, O4534, O4535, O4536, O4537, O4538, O4539, O4540, O4541, O4542, O4543, O4544, O4545, O4546, O4547, O4548, O4549, O4550, O4551, O4552, O4553, O4554, O4555, O4556, O4557, O4558, O4559, O4560, O4561, O4562, O4563, O4564, O4565, O4566, O4567, O4568, O4569, O4570, O4571, O4572, O4573, O4574, O4575, O4576, O4577, O4578, O4579, O4580, O4581, O4582, O4583, O4584, O4585, O4586, O4587, O4588, O4589, O4590, O4591, O4592, O4593, O4594, O4595, O4596, O4597, O4598, O4599, O4600, O4601, O4602, O4603, O4604, O4605, O4606, O4607, O4608, O4609, O4610, O4611, O4612, O4613, O4614, O4615, O4616, O4617, O4618, O4619, O4620, O4621, O4622, O4623, O4624, O4625, O4626, O4627, O4628, O4629, O4630, O4631, O4632, O4633, O4634, O4635, O4636, O4637, O4638, O4639, O4640, O4641, O4642, O4643, O4644, O4645, O4646, O4647, O4648, O4649, O4650, O4651, O4652, O4653, O4654, O4655, O4656, O4657, O4658, O4659, O4660, O4661, O4662, O4663, O4664, O4665, O4666, O4667, O4668, O4669, O4670, O4671, O4672, O4673, O4674, O4675, O4676, O4677, O4678, O4679, O4680, O4681, O4682, O4683, O4684, O4685, O4686, O4687, O4688, O4689, O4690, O4691, O4692, O4693, O4694, O4695, O4696, O4697, O4698, O4699, O4700, O4701, O4702, O4703, O4704, O4705, O4706, O4707, O4708, O4709, O4710, O4711, O4712, O4713, O4714, O4715, O4716, O4717, O4718, O4719, O4720, O4721, O4722, O4723, O4724, O4725, O4726, O4727, O4728, O4729, O4730, O4731, O4732, O4733, O4734, O4735, O4736, O4737, O4738, O4739, O4740, O4741, O4742, O4743, O4744, O4745, O4746, O4747, O4748, O4749, O4750, O4751, O4752, O4753, O4754, O4755, O4756, O4757, O4758, O4759, O4760, O4761, O4762, O4763, O4764, O4765, O4766, O4767, O4768, O4769, O4770, O4771, O4772, O4773, O4774, O4775, O4776, O4777, O4778, O4779, O4780, O4781, O4782, O4783, O4784, O4785, O4786, O4787, O4788, O4789, O4790, O4791, O4792, O4793, O4794, O4795, O4796, O4797, O4798, O4799, O4800, O4801, O4802, O4803, O4804, O4805, O4806, O4807, O4808, O4809, O4810, O4811, O4812, O4813, O4814, O4815, O4816, O4817, O4818, O4819, O4820, O4821, O4822, O4823, O4824, O4825, O4826, O4827, O4828, O4829, O4830, O4831, O4832, O4833, O4834, O4835, O4836, O4837, O4838, O4839, O4840, O4841, O4842, O4843, O4844, O4845, O4846, O4847, O4848, O4849, O4850, O4851, O4852, O4853, O4854, O4855, O4856, O4857, O4858, O4859, O4860, O4861, O4862, O4863, O4864, O4865, O4866, O4867, O4868, O4869, O4870, O4871, O4872, O4873, O4874, O4875, O4876, O4877, O4878, O4879, O4880, O4881, O4882, O4883, O4884, O4885, O4886, O4887, O4888, O4889, O4890, O4891, O4892, O4893, O4894, O4895, O4896, O4897, O4898, O4899, O4900, O4901, O4902, O4903, O4904, O4905, O4906, O4907, O4908, O4909, O4910, O4911, O4912, O4913, O4914, O4915, O4916, O4917, O4918, O4919, O4920, O4921, O4922, O4923, O4924, O4925, O4926, O4927, O4928, O4929, O4930, O4931, O4932, O4933, O4934, O4935, O4936, O4937, O4938, O4939, O4940, O4941, O4942, O4943, O4944, O4945, O4946, O4947, O4948, O4949, O4950, O4951, O4952, O4953, O4954, O4955, O4956, O4957, O4958, O4959, O4960, O4961, O4962, O4963, O4964, O4965, O4966, O4967, O4968, O4969, O4970, O4971, O4972, O4973, O4974, O4975, O4976, O4977, O4978, O4979, O4980, O4981, O4982, O4983, O4984, O4985, O4986, O4987, O4988, O4989, O4990, O4991, O4992, O4993, O4994, O4995, O4996, O4997, O4998, O4999, O5000, O5001, O5002, O5003, O5004, O5005, O5006, O5007, O5008, O5009, O5010, O5011, O5012, O5013, O5014, O5015, O5016, O5017, O5018, O5019, O5020, O5021, O5022, O5023, O5024, O5025, O5026, O5027, O5028, O5029, O5030, O5031, O5032, O5033, O5034, O5035, O5036, O5037, O5038, O5039, O5040, O5041, O5042, O5043, O5044, O5045, O5046, O5047, O5048, O5049, O5050, O5051, O5052, O5053, O5054, O5055, O5056, O5057, O5058, O5059, O5060, O5061, O5062, O5063, O5064, O5065, O5066, O5067, O5068, O5069, O5070, O5071, O5072, O5073, O5074, O5075, O5076, O5077, O5078, O5079, O5080, O5081, O5082, O5083, O5084, O5085, O5086, O5087, O5088, O5089, O5090, O5091, O5092, O5093, O5094, O5095, O5096, O5097, O5098, O5099, O5100, O5101, O5102, O5103, O5104, O5105, O5106, O5107, O5108, O5109, O5110, O5111, O5112, O5113, O5114, O5115, O5116, O5117, O5118, O5119, O5120, O5121, O5122, O5123, O5124, O5125, O5126, O5127, O5128, O5129, O5130, O5131, O5132, O5133, O5134, O5135, O5136, O5137, O5138, O5139, O5140, O5141, O5142, O5143, O5144, O5145, O5146, O5147, O5148, O5149, O5150, O5151, O5152, O5153, O5154, O5155, O5156, O5157, O5158, O5159, O5160, O5161, O5162, O5163, O5164, O5165, O5166, O5167, O5168, O5169, O5170, O5171, O5172, O5173, O5174, O5175, O5176, O5177, O5178, O5179, O5180, O5181, O5182, O5183, O5184, O5185, O5186, O5187, O5188, O5189, O5190, O5191, O5192, O5193, O5194, O5195, O5196, O5197, O5198, O5199, O5200, O5201, O5202, O5203, O5204, O5205, O5206, O5207, O5208, O5209, O5210, O5211, O5212, O5213, O5214, O5215, O5216, O5217, O5218, O5219, O5220, O5221, O5222, O5223, O5224, O5225, O5226, O5227, O5228, O5229, O5230, O5231, O5232, O5233, O5234, O5235, O5236, O5237, O5238, O5239, O5240, O5241, O5242, O5243, O5244, O5245, O5246, O5247, O5248, O5249, O5250, O5251, O5252, O5253, O5254, O5255, O5256, O5257, O5258, O5259, O5260, O5261, O5262, O5263, O5264, O5265, O5266, O5267, O5268, O5269, O5270, O5271, O5272, O5273, O5274, O5275, O5276, O5277, O5278, O5279, O5280, O5281, O5282, O5283, O5284, O5285, O5286, O5287, O5288, O5289, O5290, O5291, O5292, O5293, O5294, O5295, O5296, O5297, O5298, O5299, O5300, O5301, O5302, O5303, O5304, O5305, O5306, O5307, O5308, O5309, O5310, O5311, O5312, O5313, O5314, O5315, O5316, O5317, O5318, O5319, O5320, O5321, O5322, O5323, O5324, O5325, O5326, O5327, O5328, O5329, O5330, O5331, O5332, O5333, O5334, O5335, O5336, O5337, O5338, O5339, O5340, O5341, O5342, O5343, O5344, O5345, O5346, O5347, O5348, O5349, O5350, O5351, O5352, O5353, O5354, O5355, O5356, O5357, O5358, O5359, O5360, O5361, O5362, O5363, O5364, O5365, O5366, O5367, O5368, O5369, O5370, O5371, O5372, O5373, O5374, O5375, O5376, O5377, O5378, O5379, O5380, O5381, O5382, O5383, O5384, O5385, O5386, O5387, O5388, O5389, O5390, O5391, O5392, O5393, O5394, O5395, O5396, O5397, O5398, O5399, O5400, O5401, O5402, O5403, O5404, O5405, O5406, O5407, O5408, O5409, O5410, O5411, O5412, O5413, O5414, O5415, O5416, O5417, O5418, O5419, O5420, O5421, O5422, O5423, O5424, O5425, O5426, O5427, O5428, O5429, O5430, O5431, O5432, O5433, O5434, O5435, O5436, O5437, O5438, O5439, O5440, O5441, O5442, O5443, O5444, O5445, O5446, O5447, O5448, O5449, O5450, O5451, O5452, O5453, O5454, O5455, O5456, O5457, O5458, O5459, O5460, O5461, O5462, O5463, O5464, O5465, O5466, O5467, O5468, O5469, O5470, O5471, O5472, O5473, O5474, O5475, O5476, O5477, O5478, O5479, O5480, O5481, O5482, O5483, O5484, O5485, O5486, O5487, O5488, O5489, O5490, O5491, O5492, O5493, O5494, O5495, O5496, O5497, O5498, O5499, O5500, O5501, O5502, O5503, O5504, O5505, O5506, O5507, O5508, O5509, O5510, O5511, O5512, O5513, O5514, O5515, O5516, O5517, O5518, O5519, O5520, O5521, O5522, O5523, O5524, O5525, O5526, O5527, O5528, O5529, O5530, O5531, O5532, O5533, O5534, O5535, O5536, O5537, O5538, O5539, O5540, O5541, O5542, O5543, O5544, O5545, O5546, O5547, O5548, O5549, O5550, O5551, O5552, O5553, O5554, O5555, O5556, O5557, O5558, O5559, O5560, O5561, O5562, O5563, O5564, O5565, O5566, O5567, O5568, O5569, O5570, O5571, O5572, O5573, O5574, O5575, O5576, O5577, O5578, O5579, O5580, O5581, O5582, O5583, O5584, O5585, O5586, O5587, O5588, O5589, O5590, O5591, O5592, O5593, O5594, O5595, O5596, O5597, O5598, O5599, O5600, O5601, O5602, O5603, O5604, O5605, O5606, O5607, O5608, O5609, O5610, O5611, O5612, O5613, O5614, O5615, O5616, O5617, O5618, O5619, O5620, O5621, O5622, O5623, O5624, O5625, O5626, O5627, O5628, O5629, O5630, O5631, O5632, O5633, O5634, O5635, O5636, O5637, O5638, O5639, O5640, O5641, O5642, O5643, O5644, O5645, O5646, O5647, O5648, O5649, O5650, O5651, O5652, O5653, O5654, O5655, O5656, O5657, O5658, O5659, O5660, O5661, O5662, O5663, O5664, O5665, O5666, O5667, O5668, O5669, O5670, O5671, O5672, O5673, O5674, O5675, O5676, O5677, O5678, O5679, O5680, O5681, O5682, O5683, O5684, O5685, O5686, O5687, O5688, O5689, O5690, O5691, O5692, O5693, O5694, O5695, O5696, O5697, O5698, O5699, O5700, O5701, O5702, O5703, O5704, O5705, O5706, O5707, O5708, O5709, O5710, O5711, O5712, O5713, O5714, O5715, O5716, O5717, O5718, O5719, O5720, O5721, O5722, O5723, O5724, O5725, O5726, O5727, O5728, O5729, O5730, O5731, O5732, O5733, O5734, O5735, O5736, O5737, O5738, O5739, O5740, O5741, O5742, O5743, O5744, O5745, O5746, O5747, O5748, O5749, O5750, O5751, O5752, O5753, O5754, O5755, O5756, O5757, O5758, O5759, O5760, O5761, O5762, O5763, O5764, O5765, O5766, O5767, O5768, O5769, O5770, O5771, O5772, O5773, O5774, O5775, O5776, O5777, O5778, O5779, O5780, O5781, O5782, O5783, O5784, O5785, O5786, O5787, O5788, O5789, O5790, O5791, O5792, O5793, O5794, O5795, O5796, O5797, O5798, O5799, O5800, O5801, O5802, O5803, O5804, O5805, O5806, O5807, O5808, O5809, O5810, O5811, O5812, O5813, O5814, O5815, O5816, O5817, O5818, O5819, O5820, O5821, O5822, O5823, O5824, O5825, O5826, O5827, O5828, O5829, O5830, O5831, O5832, O5833, O5834, O5835, O5836, O5837, O5838, O5839, O5840, O5841, O5842, O5843, O5844, O5845, O5846, O5847, O5848, O5849, O5850, O5851, O5852, O5853, O5854, O5855, O5856, O5857, O5858, O5859, O5860, O5861, O5862, O5863, O5864, O5865, O5866, O5867, O5868, O5869, O5870, O5871, O5872, O5873, O5874, O5875, O5876, O5877, O5878, O5879, O5880, O5881, O5882, O5883, O5884, O5885, O5886, O5887, O5888, O5889, O5890, O5891, O5892, O5893, O5894, O5895, O5896, O5897, O5898, O5899, O5900, O5901, O5902, O5903, O5904, O5905, O5906, O5907, O5908, O5909, O5910, O5911, O5912, O5913, O5914, O5915, O5916, O5917, O5918, O5919, O5920, O5921, O5922, O5923, O5924, O5925, O5926, O5927, O5928, O5929, O5930, O5931, O5932, O5933, O5934, O5935, O5936, O5937, O5938, O5939, O5940, O5941, O5942, O5943, O5944, O5945, O5946, O5947, O5948, O5949, O5950, O5951, O5952, O5953, O5954, O5955, O5956, O5957, O5958, O5959, O5960, O5961, O5962, O5963, O5964, O5965, O5966, O5967, O5968, O5969, O5970, O5971, O5972, O5973, O5974, O5975, O5976, O5977, O5978, O5979, O5980, O5981, O5982, O5983, O5984, O5985, O5986, O5987, O5988, O5989, O5990, O5991, O5992, O5993, O5994, O5995, O5996, O5997, O5998, O5999, O6000, O6001, O6002, O6003, O6004, O6005, O6006, O6007, O6008, O6009, O6010, O6011, O6012, O6013, O6014, O6015, O6016, O6017, O6018, O6019, O6020, O6021, O6022, O6023, O6024, O6025, O6026, O6027, O6028, O6029, O6030, O6031, O6032, O6033, O6034, O6035, O6036, O6037, O6038, O6039, O6040, O6041, O6042, O6043, O6044, O6045, O6046, O6047, O6048, O6049, O6050, O6051, O6052, O6053, O6054, O6055, O6056, O6057, O6058, O6059, O6060, O6061, O6062, O6063, O6064, O6065, O6066, O6067, O6068, O6069, O6070, O6071, O6072, O6073, O6074, O6075, O6076, O6077, O6078, O6079, O6080, O6081, O6082, O6083, O6084, O6085, O6086, O6087, O6088, O6089, O6090, O6091, O6092, O6093, O6094, O6095, O6096, O6097, O6098, O6099, O6100, O6101, O6102, O6103, O6104, O6105, O6106, O6107, O6108, O6109, O6110, O6111, O6112, O6113, O6114, O6115, O6116, O6117, O6118, O6119, O6120, O6121, O6122, O6123, O6124, O6125, O6126, O6127, O6128, O6129, O6130, O6131, O6132, O6133, O6134, O6135, O6136, O6137, O6138, O6139, O6140, O6141, O6142, O6143, O6144, O6145, O6146, O6147, O6148, O6149, O6150, O6151, O6152, O6153, O6154, O6155, O6156, O6157, O6158, O6159, O6160, O6161, O6162, O6163, O6164, O6165, O6166, O6167, O6168, O6169, O6170, O6171, O6172, O6173, O6174, O6175, O6176, O6177, O6178, O6179, O6180, O6181, O6182, O6183, O6184, O6185, O6186, O6187, O6188, O6189, O6190, O6191, O6192, O6193, O6194, O6195, O6196, O6197, O6198, O6199, O6200, O6201, O6202, O6203, O6204, O6205, O6206, O6207, O6208, O6209, O6210, O6211, O6212, O6213, O6214, O6215, O6216, O6217, O6218, O6219, O6220, O6221, O6222, O6223, O6224, O6225, O6226, O6227, O6228, O6229, O6230, O6231, O6232, O6233, O6234, O6235, O6236, O6237, O6238, O6239, O6240, O6241, O6242, O6243, O6244, O6245, O6246, O6247, O6248, O6249, O6250, O6251, O6252, O6253, O6254, O6255, O6256, O6257, O6258, O6259, O6260, O6261, O6262, O6263, O6264, O6265, O6266, O6267, O6268, O6269, O6270, O6271, O6272, O6273, O6274, O6275, O6276, O6277, O6278, O6279, O6280, O6281, O6282, O6283, O6284, O6285, O6286, O6287, O6288, O6289, O6290, O6291, O6292, O6293, O6294, O6295, O6296, O6297, O6298, O6299, O6300, O6301, O6302, O6303, O6304, O6305, O6306, O6307, O6308, O6309, O6310, O6311, O6312, O6313, O6314, O6315, O6316, O6317, O6318, O6319, O6320, O6321, O6322, O6323, O6324, O6325, O6326, O6327, O6328, O6329, O6330, O6331, O6332, O6333, O6334, O6335, O6336, O6337, O6338, O6339, O6340, O6341, O6342, O6343, O6344, O6345, O6346, O6347, O6348, O6349, O6350, O6351, O6352, O6353, O6354, O6355, O6356, O6357, O6358, O6359, O6360, O6361, O6362, O6363, O6364, O6365, O6366, O6367, O6368, O6369, O6370, O6371, O6372, O6373, O6374, O6375, O6376, O6377, O6378, O6379, O6380, O6381, O6382, O6383, O6384, O6385, O6386, O6387, O6388, O6389, O6390, O6391, O6392, O6393, O6394, O6395, O6396, O6397, O6398, O6399, O6400, O6401, O6402, O6403, O6404, O6405, O6406, O6407, O6408, O6409, O6410, O6411, O6412, O6413, O6414, O6415, O6416, O6417, O6418, O6419, O6420, O6421, O6422, O6423, O6424, O6425, O6426, O6427, O6428, O6429, O6430, O6431, O6432, O6433, O6434, O6435, O6436, O6437, O6438, O6439, O6440, O6441, O6442, O6443, O6444, O6445, O6446, O6447, O6448, O6449, O6450, O6451, O6452, O6453, O6454, O6455, O6456, O6457, O6458, O6459, O6460, O6461, O6462, O6463, O6464, O6465, O6466, O6467, O6468, O6469, O6470, O6471, O6472, O6473, O6474, O6475, O6476, O6477, O6478, O6479, O6480, O6481, O6482, O6483, O6484, O6485, O6486, O6487, O6488, O6489, O6490, O6491, O6492, O6493, O6494, O6495, O6496, O6497, O6498, O6499, O6500, O6501, O6502, O6503, O6504, O6505, O6506, O6507, O6508, O6509, O6510, O6511, O6512, O6513, O6514, O6515, O6516, O6517, O6518, O6519, O6520, O6521, O6522, O6523, O6524, O6525, O6526, O6527, O6528, O6529, O6530, O6531, O6532, O6533, O6534, O6535, O6536, O6537, O6538, O6539, O6540, O6541, O6542, O6543, O6544, O6545, O6546, O6547, O6548, O6549, O6550, O6551, O6552, O6553, O6554, O6555, O6556, O6557, O6558, O6559, O6560, O6561, O6562, O6563, O6564, O6565, O6566, O6567, O6568, O6569, O6570, O6571, O6572, O6573, O6574, O6575, O6576, O6577, O6578, O6579, O6580, O6581, O6582, O6583, O6584, O6585, O6586, O6587, O6588, O6589, O6590, O6591, O6592, O6593, O6594, O6595, O6596, O6597, O6598, O6599, O6600, O6601, O6602, O6603, O6604, O6605, O6606, O6607, O6608, O6609, O6610, O6611, O6612, O6613, O6614, O6615, O6616, O6617, O6618, O6619, O6620, O6621, O6622, O6623, O6624, O6625, O6626, O6627, O6628, O6629, O6630, O6631, O6632, O6633, O6634, O6635, O6636, O6637, O6638, O6639, O6640, O6641, O6642, O6643, O6644, O6645, O6646, O6647, O6648, O6649, O6650, O6651, O6652, O6653, O6654, O6655, O6656, O6657, O6658, O6659, O6660, O6661, O6662, O6663, O6664, O6665, O6666, O6667, O6668, O6669, O6670, O6671, O6672, O6673, O6674, O6675, O6676, O6677, O6678, O6679, O6680, O6681, O6682, O6683, O6684, O6685, O6686, O6687, O6688, O6689, O6690, O6691, O6692, O6693, O6694, O6695, O6696, O6697, O6698, O6699, O6700, O6701, O6702, O6703, O6704, O6705, O6706, O6707, O6708, O6709, O6710, O6711, O6712, O6713, O6714, O6715, O6716, O6717, O6718, O6719, O6720, O6721, O6722, O6723, O6724, O6725, O6726, O6727, O6728, O6729, O6730, O6731, O6732, O6733, O6734, O6735, O6736, O6737, O6738, O6739, O6740, O6741, O6742, O6743, O6744, O6745, O6746, O6747, O6748, O6749, O6750, O6751, O6752, O6753, O6754, O6755, O6756, O6757, O6758, O6759, O6760, O6761, O6762, O6763, O6764, O6765, O6766, O6767, O6768, O6769, O6770, O6771, O6772, O6773, O6774, O6775, O6776, O6777, O6778, O6779, O6780, O6781, O6782, O6783, O6784, O6785, O6786, O6787, O6788, O6789, O6790, O6791, O6792, O6793, O6794, O6795, O6796, O6797, O6798, O6799, O6800, O6801, O6802, O6803, O6804, O6805, O6806, O6807, O6808, O6809, O6810, O6811, O6812, O6813, O6814, O6815, O6816, O6817, O6818, O6819, O6820, O6821, O6822, O6823, O6824, O6825, O6826, O6827, O6828, O6829, O6830, O6831, O6832, O6833, O6834, O6835, O6836, O6837, O6838, O6839, O6840, O6841, O6842, O6843, O6844, O6845, O6846, O6847, O6848, O6849, O6850, O6851, O6852, O6853, O6854, O6855, O6856, O6857, O6858, O6859, O6860, O6861, O6862, O6863, O6864, O6865, O6866, O6867, O6868, O6869, O6870, O6871, O6872, O6873, O6874, O6875, O6876, O6877, O6878, O6879, O6880, O6881, O6882, O6883, O6884, O6885, O6886, O6887, O6888, O6889, O6890, O6891, O6892, O6893, O6894, O6895, O6896, O6897, O6898, O6899, O6900, O6901, O6902, O6903, O6904, O6905, O6906, O6907, O6908, O6909, O6910, O6911, O6912, O6913, O6914, O6915, O6916, O6917, O6918, O6919, O6920, O6921, O6922, O6923, O6924, O6925, O6926, O6927, O6928, O6929, O6930, O6931, O6932, O6933, O6934, O6935, O6936, O6937, O6938, O6939, O6940, O6941, O6942, O6943, O6944, O6945, O6946, O6947, O6948, O6949, O6950, O6951, O6952, O6953, O6954, O6955, O6956, O6957, O6958, O6959, O6960, O6961, O6962, O6963, O6964, O6965, O6966, O6967, O6968, O6969, O6970, O6971, O6972, O6973, O6974, O6975, O6976, O6977, O6978, O6979, O6980, O6981, O6982, O6983, O6984, O6985, O6986, O6987, O6988, O6989, O6990, O6991, O6992, O6993, O6994, O6995, O6996, O6997, O6998, O6999, O7000, O7001, O7002, O7003, O7004, O7005, O7006, O7007, O7008, O7009, O7010, O7011, O7012, O7013, O7014, O7015, O7016, O7017, O7018, O7019, O7020, O7021, O7022, O7023, O7024, O7025, O7026, O7027, O7028, O7029, O7030, O7031, O7032, O7033, O7034, O7035, O7036, O7037, O7038, O7039, O7040, O7041, O7042, O7043, O7044, O7045, O7046, O7047, O7048, O7049, O7050, O7051, O7052, O7053, O7054, O7055, O7056, O7057, O7058, O7059, O7060, O7061, O7062, O7063, O7064, O7065, O7066, O7067, O7068, O7069, O7070, O7071, O7072, O7073, O7074, O7075, O7076, O7077, O7078, O7079, O7080, O7081, O7082, O7083, O7084, O7085, O7086, O7087, O7088, O7089, O7090, O7091, O7092, O7093, O7094, O7095, O7096, O7097, O7098, O7099, O7100, O7101, O7102, O7103, O7104, O7105, O7106, O7107, O7108, O7109, O7110, O7111, O7112, O7113, O7114, O7115, O7116, O7117, O7118, O7119, O7120, O7121, O7122, O7123, O7124, O7125, O7126, O7127, O7128, O7129, O7130, O7131, O7132, O7133, O7134, O7135, O7136, O7137, O7138, O7139, O7140, O7141, O7142, O7143, O7144, O7145, O7146, O7147, O7148, O7149, O7150, O7151, O7152, O7153, O7154, O7155, O7156, O7157, O7158, O7159, O7160, O7161, O7162, O7163, O7164, O7165, O7166, O7167, O7168, O7169, O7170, O7171, O7172, O7173, O7174, O7175, O7176, O7177, O7178, O7179, O7180, O7181, O7182, O7183, O7184, O7185, O7186, O7187, O7188, O7189, O7190, O7191, O7192, O7193, O7194, O7195, O7196, O7197, O7198, O7199, O7200, O7201, O7202, O7203, O7204, O7205, O7206, O7207, O7208, O7209, O7210, O7211, O7212, O7213, O7214, O7215, O7216, O7217, O7218, O7219, O7220, O7221, O7222, O7223, O7224, O7225, O7226, O7227, O7228, O7229, O7230, O7231, O7232, O7233, O7234, O7235, O7236, O7237, O7238, O7239, O7240, O7241, O7242, O7243, O7244, O7245, O7246, O7247, O7248, O7249, O7250, O7251, O7252, O7253, O7254, O7255, O7256, O7257, O7258, O7259, O7260, O7261, O7262, O7263, O7264, O7265, O7266, O7267, O7268, O7269, O7270, O7271, O7272, O7273, O7274, O7275, O7276, O7277, O7278, O7279, O7280, O7281, O7282, O7283, O7284, O7285, O7286, O7287, O7288, O7289, O7290, O7291, O7292, O7293, O7294, O7295, O7296, O7297, O7298, O7299, O7300, O7301, O7302, O7303, O7304, O7305, O7306, O7307, O7308, O7309, O7310, O7311, O7312, O7313, O7314, O7315, O7316, O7317, O7318, O7319, O7320, O7321, O7322, O7323, O7324, O7325, O7326, O7327, O7328, O7329, O7330, O7331, O7332, O7333, O7334, O7335, O7336, O7337, O7338, O7339, O7340, O7341, O7342, O7343, O7344, O7345, O7346, O7347, O7348, O7349, O7350, O7351, O7352, O7353, O7354, O7355, O7356, O7357, O7358, O7359, O7360, O7361, O7362, O7363, O7364, O7365, O7366, O7367, O7368, O7369, O7370, O7371, O7372, O7373, O7374, O7375, O7376, O7377, O7378, O7379, O7380, O7381, O7382, O7383, O7384, O7385, O7386, O7387, O7388, O7389, O7390, O7391, O7392, O7393, O7394, O7395, O7396, O7397, O7398, O7399, O7400, O7401, O7402, O7403, O7404, O7405, O7406, O7407, O7408, O7409, O7410, O7411, O7412, O7413, O7414, O7415, O7416, O7417, O7418, O7419, O7420, O7421, O7422, O7423, O7424, O7425, O7426, O7427, O7428, O7429, O7430, O7431, O7432, O7433, O7434, O7435, O7436, O7437, O7438, O7439, O7440, O7441, O7442, O7443, O7444, O7445, O7446, O7447, O7448, O7449, O7450, O7451, O7452, O7453, O7454, O7455, O7456, O7457, O7458, O7459, O7460, O7461, O7462, O7463, O7464, O7465, O7466, O7467, O7468, O7469, O7470, O7471, O7472, O7473, O7474, O7475, O7476, O7477, O7478, O7479, O7480, O7481, O7482, O7483, O7484, O7485, O7486, O7487, O7488, O7489, O7490, O7491, O7492, O7493, O7494, O7495, O7496, O7497, O7498, O7499, O7500, O7501, O7502, O7503, O7504, O7505, O7506, O7507, O7508, O7509, O7510, O7511, O7512, O7513, O7514, O7515, O7516, O7517, O7518, O7519, O7520, O7521, O7522, O7523, O7524, O7525, O7526, O7527, O7528, O7529, O7530, O7531, O7532, O7533, O7534, O7535, O7536, O7537, O7538, O7539, O7540, O7541, O7542, O7543, O7544, O7545, O7546, O7547, O7548, O7549, O7550, O7551, O7552, O7553, O7554, O7555, O7556, O7557, O7558, O7559, O7560, O7561, O7562, O7563, O7564, O7565, O7566, O7567, O7568, O7569, O7570, O7571, O7572, O7573, O7574, O7575, O7576, O7577, O7578, O7579, O7580, O7581, O7582, O7583, O7584, O7585, O7586, O7587, O7588, O7589, O7590, O7591, O7592, O7593, O7594, O7595, O7596, O7597, O7598, O7599, O7600, O7601, O7602, O7603, O7604, O7605, O7606, O7607, O7608, O7609, O7610, O7611, O7612, O7613, O7614, O7615, O7616, O7617, O7618, O7619, O7620, O7621, O7622, O7623, O7624, O7625, O7626, O7627, O7628, O7629, O7630, O7631, O7632, O7633, O7634, O7635, O7636, O7637, O7638, O7639, O7640, O7641, O7642, O7643, O7644, O7645, O7646, O7647, O7648, O7649, O7650, O7651, O7652, O7653, O7654, O7655, O7656, O7657, O7658, O7659, O7660, O7661, O7662, O7663, O7664, O7665, O7666, O7667, O7668, O7669, O7670, O7671, O7672, O7673, O7674, O7675, O7676, O7677, O7678, O7679, O7680, O7681, O7682, O7683, O7684, O7685, O7686, O7687, O7688, O7689, O7690, O7691, O7692, O7693, O7694, O7695, O7696, O7697, O7698, O7699, O7700, O7701, O7702, O7703, O7704, O7705, O7706, O7707, O7708, O7709, O7710, O7711, O7712, O7713, O7714, O7715, O7716, O7717, O7718, O7719, O7720, O7721, O7722, O7723, O7724, O7725, O7726, O7727, O7728, O7729, O7730, O7731, O7732, O7733, O7734, O7735, O7736, O7737, O7738, O7739, O7740, O7741, O7742, O7743, O7744, O7745, O7746, O7747, O7748, O7749, O7750, O7751, O7752, O7753, O7754, O7755, O7756, O7757, O7758, O7759, O7760, O7761, O7762, O7763, O7764, O7765, O7766, O7767, O7768, O7769, O7770, O7771, O7772, O7773, O7774, O7775, O7776, O7777, O7778, O7779, O7780, O7781, O7782, O7783, O7784, O7785, O7786, O7787, O7788, O7789, O7790, O7791, O7792, O7793, O7794, O7795, O7796, O7797, O7798, O7799, O7800, O7801, O7802, O7803, O7804, O7805, O7806, O7807, O7808, O7809, O7810, O7811, O7812, O7813, O7814, O7815, O7816, O7817, O7818, O7819, O7820, O7821, O7822, O7823, O7824, O7825, O7826, O7827, O7828, O7829, O7830, O7831, O7832, O7833, O7834, O7835, O7836, O7837, O7838, O7839, O7840, O7841, O7842, O7843, O7844, O7845, O7846, O7847, O7848, O7849, O7850, O7851, O7852, O7853, O7854, O7855, O7856, O7857, O7858, O7859, O7860, O7861, O7862, O7863, O7864, O7865, O7866, O7867, O7868, O7869, O7870, O7871, O7872, O7873, O7874, O7875, O7876, O7877, O7878, O7879, O7880, O7881, O7882, O7883, O7884, O7885, O7886, O7887, O7888, O7889, O7890, O7891, O7892, O7893, O7894, O7895, O7896, O7897, O7898, O7899, O7900, O7901, O7902, O7903, O7904, O7905, O7906, O7907, O7908, O7909, O7910, O7911, O7912, O7913, O7914, O7915, O7916, O7917, O7918, O7919, O7920, O7921, O7922, O7923, O7924, O7925, O7926, O7927, O7928, O7929, O7930, O7931, O7932, O7933, O7934, O7935, O7936, O7937, O7938, O7939, O7940, O7941, O7942, O7943, O7944, O7945, O7946, O7947, O7948, O7949, O7950, O7951, O7952, O7953, O7954, O7955, O7956, O7957, O7958, O7959, O7960, O7961, O7962, O7963, O7964, O7965, O7966, O7967, O7968, O7969, O7970, O7971, O7972, O7973, O7974, O7975, O7976, O7977, O7978, O7979, O7980, O7981, O7982, O7983, O7984, O7985, O7986, O7987, O7988, O7989, O7990, O7991, O7992, O7993, O7994, O7995, O7996, O7997, O7998, O7999, O8000, O8001, O8002, O8003, O8004, O8005, O8006, O8007, O8008, O8009, O8010, O8011, O8012, O8013, O8014, O8015, O8016, O8017, O8018, O8019, O8020, O8021, O8022, O8023, O8024, O8025, O8026, O8027, O8028, O8029, O8030, O8031, O8032, O8033, O8034, O8035, O8036, O8037, O8038, O8039, O8040, O8041, O8042, O8043, O8044, O8045, O8046, O8047, O8048, O8049, O8050, O8051, O8052, O8053, O8054, O8055, O8056, O8057, O8058, O8059, O8060, O8061, O8062, O8063, O8064, O8065, O8066, O8067, O8068, O8069, O8070, O8071, O8072, O8073, O8074, O8075, O8076, O8077, O8078, O8079, O8080, O8081, O8082, O8083, O8084, O8085, O8086, O8087, O8088, O8089, O8090, O8091, O8092, O8093, O8094, O8095, O8096, O8097, O8098, O8099, O8100, O8101, O8102, O8103, O8104, O8105, O8106, O8107, O8108, O8109, O8110, O8111, O8112, O8113, O8114, O8115, O8116, O8117, O8118, O8119, O8120, O8121, O8122, O8123, O8124, O8125, O8126, O8127, O8128, O8129, O8130, O8131, O8132, O8133, O8134, O8135, O8136, O8137, O8138, O8139, O8140, O8141, O8142, O8143, O8144, O8145, O8146, O8147, O8148, O8149, O8150, O8151, O8152, O8153, O8154, O8155, O8156, O8157, O8158, O8159, O8160, O8161, O8162, O8163, O8164, O8165, O8166, O8167, O8168, O8169, O8170, O8171, O8172, O8173, O8174, O8175, O8176, O8177, O8178, O8179, O8180, O8181, O8182, O8183, O8184, O8185, O8186, O8187, O8188, O8189, O8190, O8191, O8192, O8193, O8194, O8195, O8196, O8197, O8198, O8199, O8200, O8201, O8202, O8203, O8204, O8205, O8206, O8207, O8208, O8209, O8210, O8211, O8212, O8213, O8214, O8215, O8216, O8217, O8218, O8219, O8220, O8221, O8222, O8223, O8224, O8225, O8226, O8227, O8228, O8229, O8230, O8231, O8232, O8233, O8234, O8235, O8236, O8237, O8238, O8239, O8240, O8241, O8242, O8243, O8244, O8245, O8246, O8247, O8248, O8249, O8250, O8251, O8252, O8253, O8254, O8255, O8256, O8257, O8258, O8259, O8260, O8261, O8262, O8263, O8264, O8265, O8266, O8267, O8268, O8269, O8270, O8271, O8272, O8273, O8274, O8275, O8276, O8277, O8278, O8279, O8280, O8281, O8282, O8283, O8284, O8285, O8286, O8287, O8288, O8289, O8290, O8291, O8292, O8293, O8294, O8295, O8296, O8297, O8298, O8299, O8300, O8301, O8302, O8303, O8304, O8305, O8306, O8307, O8308, O8309, O8310, O8311, O8312, O8313, O8314, O8315, O8316, O8317, O8318, O8319, O8320, O8321, O8322, O8323, O8324, O8325, O8326, O8327, O8328, O8329, O8330, O8331, O8332, O8333, O8334, O8335, O8336, O8337, O8338, O8339, O8340, O8341, O8342, O8343, O8344, O8345, O8346, O8347, O8348, O8349, O8350, O8351, O8352, O8353, O8354, O8355, O8356, O8357, O8358, O8359, O8360, O8361, O8362, O8363, O8364, O8365, O8366, O8367, O8368, O8369, O8370, O8371, O8372, O8373, O8374, O8375, O8376, O8377, O8378, O8379, O8380, O8381, O8382, O8383, O8384, O8385, O8386, O8387, O8388, O8389, O8390, O8391, O8392, O8393, O8394, O8395, O8396, O8397, O8398, O8399, O8400, O8401, O8402, O8403, O8404, O8405, O8406, O8407, O8408, O8409, O8410, O8411, O8412, O8413, O8414, O8415, O8416, O8417, O8418, O8419, O8420, O8421, O8422, O8423, O8424, O8425, O8426, O8427, O8428, O8429, O8430, O8431, O8432, O8433, O8434, O8435, O8436, O8437, O8438, O8439, O8440, O8441, O8442, O8443, O8444, O8445, O8446, O8447, O8448, O8449, O8450, O8451, O8452, O8453, O8454, O8455, O8456, O8457, O8458, O8459, O8460, O8461, O8462, O8463, O8464, O8465, O8466, O8467, O8468, O8469, O8470, O8471, O8472, O8473, O8474, O8475, O8476, O8477, O8478, O8479, O8480, O8481, O8482, O8483, O8484, O8485, O8486, O8487, O8488, O8489, O8490, O8491, O8492, O8493, O8494, O8495, O8496, O8497, O8498, O8499, O8500, O8501, O8502, O8503, O8504, O8505, O8506, O8507, O8508, O8509, O8510, O8511, O8512, O8513, O8514, O8515, O8516, O8517, O8518, O8519, O8520, O8521, O8522, O8523, O8524, O8525, O8526, O8527, O8528, O8529, O8530, O8531, O8532, O8533, O8534, O8535, O8536, O8537, O8538, O8539, O8540, O8541, O8542, O8543, O8544, O8545, O8546, O8547, O8548, O8549, O8550, O8551, O8552, O8553, O8554, O8555, O8556, O8557, O8558, O8559, O8560, O8561, O8562, O8563, O8564, O8565, O8566, O8567, O8568, O8569, O8570, O8571, O8572, O8573, O8574, O8575, O8576, O8577, O8578, O8579, O8580, O8581, O8582, O8583, O8584, O8585, O8586, O8587, O8588, O8589, O8590, O8591, O8592, O8593, O8594, O8595, O8596, O8597, O8598, O8599, O8600, O8601, O8602, O8603, O8604, O8605, O8606, O8607, O8608, O8609, O8610, O8611, O8612, O8613, O8614, O8615, O8616, O8617, O8618, O8619, O8620, O8621, O8622, O8623, O8624, O8625, O8626, O8627, O8628, O8629, O8630, O8631, O8632, O8633, O8634, O8635, O8636, O8637, O8638, O8639, O8640, O8641, O8642, O8643, O8644, O8645, O8646, O8647, O8648, O8649, O8650, O8651, O8652, O8653, O8654, O8655, O8656, O8657, O8658, O8659, O8660, O8661, O8662, O8663, O8664, O8665, O8666, O8667, O8668, O8669, O8670, O8671, O8672, O8673, O8674, O8675, O8676, O8677, O8678, O8679, O8680, O8681, O8682, O8683, O8684, O8685, O8686, O8687, O8688, O8689, O8690, O8691, O8692, O8693, O8694, O8695, O8696, O8697, O8698, O8699, O8700, O8701, O8702, O8703, O8704, O8705, O8706, O8707, O8708, O8709, O8710, O8711, O8712, O8713, O8714, O8715, O8716, O8717, O8718, O8719, O8720, O8721, O8722, O8723, O8724, O8725, O8726, O8727, O8728, O8729, O8730, O8731, O8732, O8733, O8734, O8735, O8736, O8737, O8738, O8739, O8740, O8741, O8742, O8743, O8744, O8745, O8746, O8747, O8748, O8749, O8750, O8751, O8752, O8753, O8754, O8755, O8756, O8757, O8758, O8759, O8760, O8761, O8762, O8763, O8764, O8765, O8766, O8767, O8768, O8769, O8770, O8771, O8772, O8773, O8774, O8775, O8776, O8777, O8778, O8779, O8780, O8781, O8782, O8783, O8784, O8785, O8786, O8787, O8788, O8789, O8790, O8791, O8792, O8793, O8794, O8795, O8796, O8797, O8798, O8799, O8800, O8801, O8802, O8803, O8804, O8805, O8806, O8807, O8808, O8809, O8810, O8811, O8812, O8813, O8814, O8815, O8816, O8817, O8818, O8819, O8820, O8821, O8822, O8823, O8824, O8825, O8826, O8827, O8828, O8829, O8830, O8831, O8832, O8833, O8834, O8835, O8836, O8837, O8838, O8839, O8840, O8841, O8842, O8843, O8844, O8845, O8846, O8847, O8848, O8849, O8850, O8851, O8852, O8853, O8854, O8855, O8856, O8857, O8858, O8859, O8860, O8861, O8862, O8863, O8864, O8865, O8866, O8867, O8868, O8869, O8870, O8871, O8872, O8873, O8874, O8875, O8876, O8877, O8878, O8879, O8880, O8881, O8882, O8883, O8884, O8885, O8886, O8887, O8888, O8889, O8890, O8891, O8892, O8893, O8894, O8895, O8896, O8897, O8898, O8899, O8900, O8901, O8902, O8903, O8904, O8905, O8906, O8907, O8908, O8909, O8910, O8911, O8912, O8913, O8914, O8915, O8916, O8917, O8918, O8919, O8920, O8921, O8922, O8923, O8924, O8925, O8926, O8927, O8928, O8929, O8930, O8931, O8932, O8933, O8934, O8935, O8936, O8937, O8938, O8939, O8940, O8941, O8942, O8943, O8944, O8945, O8946, O8947, O8948, O8949, O8950, O8951, O8952, O8953, O8954, O8955, O8956, O8957, O8958, O8959, O8960, O8961, O8962, O8963, O8964, O8965, O8966, O8967, O8968, O8969, O8970, O8971, O8972, O8973, O8974, O8975, O8976, O8977, O8978, O8979, O8980, O8981, O8982, O8983, O8984, O8985, O8986, O8987, O8988, O8989, O8990, O8991, O8992, O8993, O8994, O8995, O8996, O8997, O8998, O8999, O9000, O9001, O9002, O9003, O9004, O9005, O9006, O9007, O9008, O9009, O9010, O9011, O9012, O9013, O9014, O9015, O9016, O9017, O9018, O9019, O9020, O9021, O9022, O9023, O9024, O9025, O9026, O9027, O9028, O9029, O9030, O9031, O9032, O9033, O9034, O9035, O9036, O9037, O9038, O9039, O9040, O9041, O9042, O9043, O9044, O9045, O9046, O9047, O9048, O9049, O9050, O9051, O9052, O9053, O9054, O9055, O9056, O9057, O9058, O9059, O9060, O9061, O9062, O9063, O9064, O9065, O9066, O9067, O9068, O9069, O9070, O9071, O9072, O9073, O9074, O9075, O9076, O9077, O9078, O9079, O9080, O9081, O9082, O9083, O9084, O9085, O9086, O9087, O9088, O9089, O9090, O9091, O9092, O9093, O9094, O9095, O9096, O9097, O9098, O9099, O9100, O9101, O9102, O9103, O9104, O9105, O9106, O9107, O9108, O9109, O9110, O9111, O9112, O9113, O9114, O9115, O9116, O9117, O9118, O9119, O9120, O9121, O9122, O9123, O9124, O9125, O9126, O9127, O9128, O9129, O9130, O9131, O9132, O9133, O9134, O9135, O9136, O9137, O9138, O9139, O9140, O9141, O9142, O9143, O9144, O9145, O9146, O9147, O9148, O9149, O9150, O9151, O9152, O9153, O9154, O9155, O9156, O9157, O9158, O9159, O9160, O9161, O9162, O9163, O9164, O9165, O9166, O9167, O9168, O9169, O9170, O9171, O9172, O9173, O9174, O9175, O9176, O9177, O9178, O9179, O9180, O9181, O9182, O9183, O9184, O9185, O9186, O9187, O9188, O9189, O9190, O9191, O9192, O9193, O9194, O9195, O9196, O9197, O9198, O9199, O9200, O9201, O9202, O9203, O9204, O9205, O9206, O9207, O9208, O9209, O9210, O9211, O9212, O9213, O9214, O9215, O9216, O9217, O9218, O9219, O9220, O9221, O9222, O9223, O9224, O9225, O9226, O9227, O9228, O9229, O9230, O9231, O9232, O9233, O9234, O9235, O9236, O9237, O9238, O9239, O9240, O9241, O9242, O9243, O9244, O9245, O9246, O9247, O9248, O9249, O9250, O9251, O9252, O9253, O9254, O9255, O9256, O9257, O9258, O9259, O9260, O9261, O9262, O9263, O9264, O9265, O9266, O9267, O9268, O9269, O9270, O9271, O9272, O9273, O9274, O9275, O9276, O9277, O9278, O9279, O9280, O9281, O9282, O9283, O9284, O9285, O9286, O9287, O9288, O9289, O9290, O9291, O9292, O9293, O9294, O9295, O9296, O9297, O9298, O9299, O9300, O9301, O9302, O9303, O9304, O9305, O9306, O9307, O9308, O9309, O9310, O9311, O9312, O9313, O9314, O9315, O9316, O9317, O9318, O9319, O9320, O9321, O9322, O9323, O9324, O9325, O9326, O9327, O9328, O9329, O9330, O9331, O9332, O9333, O9334, O9335, O9336, O9337, O9338, O9339, O9340, O9341, O9342, O9343, O9344, O9345, O9346, O9347, O9348, O9349, O9350, O9351, O9352, O9353, O9354, O9355, O9356, O9357, O9358, O9359, O9360, O9361, O9362, O9363, O9364, O9365, O9366, O9367, O9368, O9369, O9370, O9371, O9372, O9373, O9374, O9375, O9376, O9377, O9378, O9379, O9380, O9381, O9382, O9383, O9384, O9385, O9386, O9387, O9388, O9389, O9390, O9391, O9392, O9393, O9394, O9395, O9396, O9397, O9398, O9399, O9400, O9401, O9402, O9403, O9404, O9405, O9406, O9407, O9408, O9409, O9410, O9411, O9412, O9413, O9414, O9415, O9416, O9417, O9418, O9419, O9420, O9421, O9422, O9423, O9424, O9425, O9426, O9427, O9428, O9429, O9430, O9431, O9432, O9433, O9434, O9435, O9436, O9437, O9438, O9439, O9440, O9441, O9442, O9443, O9444, O9445, O9446, O9447, O9448, O9449, O9450, O9451, O9452, O9453, O9454, O9455, O9456, O9457, O9458, O9459, O9460, O9461, O9462, O9463, O9464, O9465, O9466, O9467, O9468, O9469, O9470, O9471, O9472, O9473, O9474, O9475, O9476, O9477, O9478, O9479, O9480, O9481, O9482, O9483, O9484, O9485, O9486, O9487, O9488, O9489, O9490, O9491, O9492, O9493, O9494, O9495, O9496, O9497, O9498, O9499, O9500, O9501, O9502, O9503, O9504, O9505, O9506, O9507, O9508, O9509, O9510, O9511, O9512, O9513, O9514, O9515, O9516, O9517, O9518, O9519, O9520, O9521, O9522, O9523, O9524, O9525, O9526, O9527, O9528, O9529, O9530, O9531, O9532, O9533, O9534, O9535, O9536, O9537, O9538, O9539, O9540, O9541, O9542, O9543, O9544, O9545, O9546, O9547, O9548, O9549, O9550, O9551, O9552, O9553, O9554, O9555, O9556, O9557, O9558, O9559, O9560, O9561, O9562, O9563, O9564, O9565, O9566, O9567, O9568, O9569, O9570, O9571, O9572, O9573, O9574, O9575, O9576, O9577, O9578, O9579, O9580, O9581, O9582, O9583, O9584, O9585, O9586, O9587, O9588, O9589, O9590, O9591, O9592, O9593, O9594, O9595, O9596, O9597, O9598, O9599, O9600, O9601, O9602, O9603, O9604, O9605, O9606, O9607, O9608, O9609, O9610, O9611, O9612, O9613, O9614, O9615, O9616, O9617, O9618, O9619, O9620, O9621, O9622, O9623, O9624, O9625, O9626, O9627, O9628, O9629, O9630, O9631, O9632, O9633, O9634, O9635, O9636, O9637, O9638, O9639, O9640, O9641, O9642, O9643, O9644, O9645, O9646, O9647, O9648, O9649, O9650, O9651, O9652, O9653, O9654, O9655, O9656, O9657, O9658, O9659, O9660, O9661, O9662, O9663, O9664, O9665, O9666, O9667, O9668, O9669, O9670, O9671, O9672, O9673, O9674, O9675, O9676, O9677, O9678, O9679, O9680, O9681, O9682, O9683, O9684, O9685, O9686, O9687, O9688, O9689, O9690, O9691, O9692, O9693, O9694, O9695, O9696, O9697, O9698, O9699, O9700, O9701, O9702, O9703, O9704, O9705, O9706, O9707, O9708, O9709, O9710, O9711, O9712, O9713, O9714, O9715, O9716, O9717, O9718, O9719, O9720, O9721, O9722, O9723, O9724, O9725, O9726, O9727, O9728, O9729, O9730, O9731, O9732, O9733, O9734, O9735, O9736, O9737, O9738, O9739, O9740, O9741, O9742, O9743, O9744, O9745, O9746, O9747, O9748, O9749, O9750, O9751, O9752, O9753, O9754, O9755, O9756, O9757, O9758, O9759, O9760, O9761, O9762, O9763, O9764, O9765, O9766, O9767, O9768, O9769, O9770, O9771, O9772, O9773, O9774, O9775, O9776, O9777, O9778, O9779, O9780, O9781, O9782, O9783, O9784, O9785, O9786, O9787, O9788, O9789, O9790, O9791, O9792, O9793, O9794, O9795, O9796, O9797, O9798, O9799, O9800, O9801, O9802, O9803, O9804, O9805, O9806, O9807, O9808, O9809, O9810, O9811, O9812, O9813, O9814, O9815, O9816, O9817, O9818, O9819, O9820, O9821, O9822, O9823, O9824, O9825, O9826, O9827, O9828, O9829, O9830, O9831, O9832, O9833, O9834, O9835, O9836, O9837, O9838, O9839, O9840, O9841, O9842, O9843, O9844, O9845, O9846, O9847, O9848, O9849, O9850, O9851, O9852, O9853, O9854, O9855, O9856, O9857, O9858, O9859, O9860, O9861, O9862, O9863, O9864, O9865, O9866, O9867, O9868, O9869, O9870, O9871, O9872, O9873, O9874, O9875, O9876, O9877, O9878, O9879, O9880, O9881, O9882, O9883, O9884, O9885, O9886, O9887, O9888, O9889, O9890, O9891, O9892, O9893, O9894, O9895, O9896, O9897, O9898, O9899, O9900, O9901, O9902, O9903, O9904, O9905, O9906, O9907, O9908, O9909, O9910, O9911, O9912, O9913, O9914, O9915, O9916, O9917, O9918, O9919, O9920, O9921, O9922, O9923, O9924, O9925, O9926, O9927, O9928, O9929, O9930, O9931, O9932, O9933, O9934, O9935, O9936, O9937, O9938, O9939, O9940, O9941, O9942, O9943, O9944, O9945, O9946, O9947, O9948, O9949, O9950, O9951, O9952, O9953, O9954, O9955, O9956, O9957, O9958, O9959, O9960, O9961, O9962, O9963, O9964, O9965, O9966, O9967, O9968, O9969, O9970, O9971, O9972, O9973, O9974, O9975, O9976, O9977, O9978, O9979, O9980, O9981, O9982, O9983, O9984, O9985, O9986, O9987, O9988, O9989, O9990, O9991, O9992, O9993, O9994, O9995, O9996, O9997, O9998, O9999, O10000, O10001, O10002, O10003, O10004, O10005, O10006, O10007, O10008, O10009, O10010, O10011, O10012, O10013, O10014, O10015, O10016, O10017, O10018, O10019, O10020, O10021, O10022, O10023, O10024, O10025, O10026, O10027, O10028, O10029, O10030, O10031, O10032, O10033, O10034, O10035, O10036, O10037, O10038, O10039, O10040, O10041, O10042, O10043, O10044, O10045, O10046, O10047, O10048, O10049, O10050, O10051, O10052, O10053, O10054, O10055, O10056, O10057, O10058, O10059, O10060, O10061, O10062, O10063, O10064, O10065, O10066, O10067, O10068, O10069, O10070, O10071, O10072, O10073, O10074, O10075, O10076, O10077, O10078, O10079, O10080, O10081, O10082, O10083, O10084, O10085, O10086, O10087, O10088, O10089, O10090, O10091, O10092, O10093, O10094, O10095, O10096, O10097, O10098, O10099, O10100, O10101, O10102, O10103, O10104, O10105, O10106, O10107, O10108, O10109, O10110, O10111, O10112, O10113, O10114, O10115, O10116, O10117, O10118, O10119, O10120, O10121, O10122, O10123, O10124, O10125, O10126, O10127, O10128, O10129, O10130, O10131, O10132, O10133, O10134, O10135, O10136, O10137, O10138, O10139, O10140, O10141, O10142, O10143, O10144, O10145, O10146, O10147, O10148, O10149, O10150, O10151, O10152, O10153, O10154, O10155, O10156, O10157, O10158, O10159, O10160, O10161, O10162, O10163, O10164, O10165, O10166, O10167, O10168, O10169, O10170, O10171, O10172, O10173, O10174, O10175, O10176, O10177, O10178, O10179, O10180, O10181, O10182, O10183, O10184, O10185, O10186, O10187, O10188, O10189, O10190, O10191, O10192, O10193, O10194, O10195, O10196, O10197, O10198, O10199, O10200, O10201, O10202, O10203, O10204, O10205, O10206, O10207, O10208, O10209, O10210, O10211, O10212, O10213, O10214, O10215, O10216, O10217, O10218, O10219, O10220, O10221, O10222, O10223, O10224, O10225, O10226, O10227, O10228, O10229, O10230, O10231, O10232, O10233, O10234, O10235, O10236, O10237, O10238, O10239, O10240, O10241, O10242, O10243, O10244, O10245, O10246, O10247, O10248, O10249, O10250, O10251, O10252, O10253, O10254, O10255, O10256, O10257, O10258, O10259, O10260, O10261, O10262, O10263, O10264, O10265, O10266, O10267, O10268, O10269, O10270, O10271, O10272, O10273, O10274, O10275, O10276, O10277, O10278, O10279, O10280, O10281, O10282, O10283, O10284, O10285, O10286, O10287, O10288, O10289, O10290, O10291, O10292, O10293, O10294, O10295, O10296, O10297, O10298, O10299, O10300, O10301, O10302, O10303, O10304, O10305, O10306, O10307, O10308, O10309, O10310, O10311, O10312, O10313, O10314, O10315, O10316, O10317, O10318, O10319, O10320, O10321, O10322, O10323, O10324, O10325, O10326, O10327, O10328, O10329, O10330, O10331, O10332, O10333, O10334, O10335, O10336, O10337, O10338, O10339, O10340, O10341, O10342, O10343, O10344, O10345, O10346, O10347, O10348, O10349, O10350, O10351, O10352, O10353, O10354, O10355, O10356, O10357, O10358, O10359, O10360, O10361, O10362, O10363, O10364, O10365, O10366, O10367, O10368, O10369, O10370, O10371, O10372, O10373, O10374, O10375, O10376, O10377, O10378, O10379, O10380, O10381, O10382, O10383, O10384, O10385, O10386, O10387, O10388, O10389, O10390, O10391, O10392, O10393, O10394, O10395, O10396, O10397, O10398, O10399, O10400, O10401, O10402, O10403, O10404, O10405, O10406, O10407, O10408, O10409, O10410, O10411, O10412, O10413, O10414, O10415, O10416, O10417, O10418, O10419, O10420, O10421, O10422, O10423, O10424, O10425, O10426, O10427, O10428, O10429, O10430, O10431, O10432, O10433, O10434, O10435, O10436, O10437, O10438, O10439, O10440, O10441, O10442, O10443, O10444, O10445, O10446, O10447, O10448, O10449, O10450, O10451, O10452, O10453, O10454, O10455, O10456, O10457, O10458, O10459, O10460, O10461, O10462, O10463, O10464, O10465, O10466, O10467, O10468, O10469, O10470, O10471, O10472, O10473, O10474, O10475, O10476, O10477, O10478, O10479, O10480, O10481, O10482, O10483, O10484, O10485, O10486, O10487, O10488, O10489, O10490, O10491, O10492, O10493, O10494, O10495, O10496, O10497, O10498, O10499, O10500, O10501, O10502, O10503, O10504, O10505, O10506, O10507, O10508, O10509, O10510, O10511, O10512, O10513, O10514, O10515, O10516, O10517, O10518, O10519, O10520, O10521, O10522, O10523, O10524, O10525, O10526, O10527, O10528, O10529, O10530, O10531, O10532, O10533, O10534, O10535, O10536, O10537, O10538, O10539, O10540, O10541, O10542, O10543, O10544, O10545, O10546, O10547, O10548, O10549, O10550, O10551, O10552, O10553, O10554, O10555, O10556, O10557, O10558, O10559, O10560, O10561, O10562, O10563, O10564, O10565, O10566, O10567, O10568, O10569, O10570, O10571, O10572, O10573, O10574, O10575, O10576, O10577, O10578, O10579, O10580, O10581, O10582, O10583, O10584, O10585, O10586, O10587, O10588, O10589, O10590, O10591, O10592, O10593, O10594, O10595, O10596, O10597, O10598, O10599, O10600, O10601, O10602, O10603, O10604, O10605, O10606, O10607, O10608, O10609, O10610, O10611, O10612, O10613, O10614, O10615, O10616, O10617, O10618, O10619, O10620, O10621, O10622, O10623, O10624, O10625, O10626, O10627, O10628, O10629, O10630, O10631, O10632, O10633, O10634, O10635, O10636, O10637, O10638, O10639, O10640, O10641, O10642, O10643, O10644, O10645, O10646, O10647, O10648, O10649, O10650, O10651, O10652, O10653, O10654, O10655, O10656, O10657, O10658, O10659, O10660, O10661, O10662, O10663, O10664, O10665, O10666, O10667, O10668, O10669, O10670, O10671, O10672, O10673, O10674, O10675, O10676, O10677, O10678, O10679, O10680, O10681, O10682, O10683, O10684, O10685, O10686, O10687, O10688, O10689, O10690, O10691, O10692, O10693, O10694, O10695, O10696, O10697, O10698, O10699, O10700, O10701, O10702, O10703, O10704, O10705, O10706, O10707, O10708, O10709, O10710, O10711, O10712, O10713, O10714, O10715, O10716, O10717, O10718, O10719, O10720, O10721, O10722, O10723, O10724, O10725, O10726, O10727, O10728, O10729, O10730, O10731, O10732, O10733, O10734, O10735, O10736, O10737, O10738, O10739, O10740, O10741, O10742, O10743, O10744, O10745, O10746, O10747, O10748, O10749, O10750, O10751, O10752, O10753, O10754, O10755, O10756, O10757, O10758, O10759, O10760, O10761, O10762, O10763, O10764, O10765, O10766, O10767, O10768, O10769, O10770, O10771, O10772, O10773, O10774, O10775, O10776, O10777, O10778, O10779, O10780, O10781, O10782, O10783, O10784, O10785, O10786, O10787, O10788, O10789, O10790, O10791, O10792, O10793, O10794, O10795, O10796, O10797, O10798, O10799, O10800, O10801, O10802, O10803, O10804, O10805, O10806, O10807, O10808, O10809, O10810, O10811, O10812, O10813, O10814, O10815, O10816, O10817, O10818, O10819, O10820, O10821, O10822, O10823, O10824, O10825, O10826, O10827, O10828, O10829, O10830, O10831, O10832, O10833, O10834, O10835, O10836, O10837, O10838, O10839, O10840, O10841, O10842, O10843, O10844, O10845, O10846, O10847, O10848, O10849, O10850, O10851, O10852, O10853, O10854, O10855, O10856, O10857, O10858, O10859, O10860, O10861, O10862, O10863, O10864, O10865, O10866, O10867, O10868, O10869, O10870, O10871, O10872, O10873, O10874, O10875, O10876, O10877, O10878, O10879, O10880, O10881, O10882, O10883, O10884, O10885, O10886, O10887, O10888, O10889, O10890, O10891, O10892, O10893, O10894, O10895, O10896, O10897, O10898, O10899, O10900, O10901, O10902, O10903, O10904, O10905, O10906, O10907, O10908, O10909, O10910, O10911, O10912, O10913, O10914, O10915, O10916, O10917, O10918, O10919, O10920, O10921, O10922, O10923, O10924, O10925, O10926, O10927, O10928, O10929, O10930, O10931, O10932, O10933, O10934, O10935, O10936, O10937, O10938, O10939, O10940, O10941, O10942, O10943, O10944, O10945, O10946, O10947, O10948, O10949, O10950, O10951, O10952, O10953, O10954, O10955, O10956, O10957, O10958, O10959, O10960, O10961, O10962, O10963, O10964, O10965, O10966, O10967, O10968, O10969, O10970, O10971, O10972, O10973, O10974, O10975, O10976, O10977, O10978, O10979, O10980, O10981, O10982, O10983, O10984, O10985, O10986, O10987, O10988, O10989, O10990, O10991, O10992, O10993, O10994, O10995, O10996, O10997, O10998, O10999, O11000, O11001, O11002, O11003, O11004, O11005, O11006, O11007, O11008, O11009, O11010, O11011, O11012, O11013, O11014, O11015, O11016, O11017, O11018, O11019, O11020, O11021, O11022, O11023, O11024, O11025, O11026, O11027, O11028, O11029, O11030, O11031, O11032, O11033, O11034, O11035, O11036, O11037, O11038, O11039, O11040, O11041, O11042, O11043, O11044, O11045, O11046, O11047, O11048, O11049, O11050, O11051, O11052, O11053, O11054, O11055, O11056, O11057, O11058, O11059, O11060, O11061, O11062, O11063, O11064, O11065, O11066, O11067, O11068, O11069, O11070, O11071, O11072, O11073, O11074, O11075, O11076, O11077, O11078, O11079, O11080, O11081, O11082, O11083, O11084, O11085, O11086, O11087, O11088, O11089, O11090, O11091, O11092, O11093, O11094, O11095, O11096, O11097, O11098, O11099, O11100, O11101, O11102, O11103, O11104, O11105, O11106, O11107, O11108, O11109, O11110, O11111, O11112, O11113, O11114, O11115, O11116, O11117, O11118, O11119, O11120, O11121, O11122, O11123, O11124, O11125, O11126, O11127, O11128, O11129, O11130, O11131, O11132, O11133, O11134, O11135, O11136, O11137, O11138, O11139, O11140, O11141, O11142, O11143, O11144, O11145, O11146, O11147, O11148, O11149, O11150, O11151, O11152, O11153, O11154, O11155, O11156, O11157, O11158, O11159, O11160, O11161, O11162, O11163, O11164, O11165, O11166, O11167, O11168, O11169, O11170, O11171, O11172, O11173, O11174, O11175, O11176, O11177, O11178, O11179, O11180, O11181, O11182, O11183, O11184, O11185, O11186, O11187, O11188, O11189, O11190, O11191, O11192, O11193, O11194, O11195, O11196, O11197, O11198, O11199, O11200, O11201, O11202, O11203, O11204, O11205, O11206, O11207, O11208, O11209, O11210, O11211, O11212, O11213, O11214, O11215, O11216, O11217, O11218, O11219, O11220, O11221, O11222, O11223, O11224, O11225, O11226, O11227, O11228, O11229, O11230, O11231, O11232, O11233, O11234, O11235, O11236, O11237, O11238, O11239, O11240, O11241, O11242, O11243, O11244, O11245, O11246, O11247, O11248, O11249, O11250, O11251, O11252, O11253, O11254, O11255, O11256, O11257, O11258, O11259, O11260, O11261, O11262, O11263, O11264, O11265, O11266, O11267, O11268, O11269, O11270, O11271, O11272, O11273, O11274, O11275, O11276, O11277, O11278, O11279, O11280, O11281, O11282, O11283, O11284, O11285, O11286, O11287, O11288, O11289, O11290, O11291, O11292, O11293, O11294, O11295, O11296, O11297, O11298, O11299, O11300, O11301, O11302, O11303, O11304, O11305, O11306, O11307, O11308, O11309, O11310, O11311, O11312, O11313, O11314, O11315, O11316, O11317, O11318, O11319, O11320, O11321, O11322, O11323, O11324, O11325, O11326, O11327, O11328, O11329, O11330, O11331, O11332, O11333, O11334, O11335, O11336, O11337, O11338, O11339, O11340, O11341, O11342, O11343, O11344, O11345, O11346, O11347, O11348, O11349, O11350, O11351, O11352, O11353, O11354, O11355, O11356, O11357, O11358, O11359, O11360, O11361, O11362, O11363, O11364, O11365, O11366, O11367, O11368, O11369, O11370, O11371, O11372, O11373, O11374, O11375, O11376, O11377, O11378, O11379, O11380, O11381, O11382, O11383, O11384, O11385, O11386, O11387, O11388, O11389, O11390, O11391, O11392, O11393, O11394, O11395, O11396, O11397, O11398, O11399, O11400, O11401, O11402, O11403, O11404, O11405, O11406, O11407, O11408, O11409, O11410, O11411, O11412, O11413, O11414, O11415, O11416, O11417, O11418, O11419, O11420, O11421, O11422, O11423, O11424, O11425, O11426, O11427, O11428, O11429, O11430, O11431, O11432, O11433, O11434, O11435, O11436, O11437, O11438, O11439, O11440, O11441, O11442, O11443, O11444, O11445, O11446, O11447, O11448, O11449, O11450, O11451, O11452, O11453, O11454, O11455, O11456, O11457, O11458, O11459, O11460, O11461, O11462, O11463, O11464, O11465, O11466, O11467, O11468, O11469, O11470, O11471, O11472, O11473, O11474, O11475, O11476, O11477, O11478, O11479, O11480, O11481, O11482, O11483, O11484, O11485, O11486, O11487, O11488, O11489, O11490, O11491, O11492, O11493, O11494, O11495, O11496, O11497, O11498, O11499, O11500, O11501, O11502, O11503, O11504, O11505, O11506, O11507, O11508, O11509, O11510, O11511, O11512, O11513, O11514, O11515, O11516, O11517, O11518, O11519, O11520, O11521, O11522, O11523, O11524, O11525, O11526, O11527, O11528, O11529, O11530, O11531, O11532, O11533, O11534, O11535, O11536, O11537, O11538, O11539, O11540, O11541, O11542, O11543, O11544, O11545, O11546, O11547, O11548, O11549, O11550, O11551, O11552, O11553, O11554, O11555, O11556, O11557, O11558, O11559, O11560, O11561, O11562, O11563, O11564, O11565, O11566, O11567, O11568, O11569, O11570, O11571, O11572, O11573, O11574, O11575, O11576, O11577, O11578, O11579, O11580, O11581, O11582, O11583, O11584, O11585, O11586, O11587, O11588, O11589, O11590, O11591, O11592, O11593, O11594, O11595, O11596, O11597, O11598, O11599, O11600, O11601, O11602, O11603, O11604, O11605, O11606, O11607, O11608, O11609, O11610, O11611, O11612, O11613, O11614, O11615, O11616, O11617, O11618, O11619, O11620, O11621, O11622, O11623, O11624, O11625, O11626, O11627, O11628, O11629, O11630, O11631, O11632, O11633, O11634, O11635, O11636, O11637, O11638, O11639, O11640, O11641, O11642, O11643, O11644, O11645, O11646, O11647, O11648, O11649, O11650, O11651, O11652, O11653, O11654, O11655, O11656, O11657, O11658, O11659, O11660, O11661, O11662, O11663, O11664, O11665, O11666, O11667, O11668, O11669, O11670, O11671, O11672, O11673, O11674, O11675, O11676, O11677, O11678, O11679, O11680, O11681, O11682, O11683, O11684, O11685, O11686, O11687, O11688, O11689, O11690, O11691, O11692, O11693, O11694, O11695, O11696, O11697, O11698, O11699, O11700, O11701, O11702, O11703, O11704, O11705, O11706, O11707, O11708, O11709, O11710, O11711, O11712, O11713, O11714, O11715, O11716, O11717, O11718, O11719, O11720, O11721, O11722, O11723, O11724, O11725, O11726, O11727, O11728, O11729, O11730, O11731, O11732, O11733, O11734, O11735, O11736, O11737, O11738, O11739, O11740, O11741, O11742, O11743, O11744, O11745, O11746, O11747, O11748, O11749, O11750, O11751, O11752, O11753, O11754, O11755, O11756, O11757, O11758, O11759, O11760, O11761, O11762, O11763, O11764, O11765, O11766, O11767, O11768, O11769, O11770, O11771, O11772, O11773, O11774, O11775, O11776, O11777, O11778, O11779, O11780, O11781, O11782, O11783, O11784, O11785, O11786, O11787, O11788, O11789, O11790, O11791, O11792, O11793, O11794, O11795, O11796, O11797, O11798, O11799, O11800, O11801, O11802, O11803, O11804, O11805, O11806, O11807, O11808, O11809, O11810, O11811, O11812, O11813, O11814, O11815, O11816, O11817, O11818, O11819, O11820, O11821, O11822, O11823, O11824, O11825, O11826, O11827, O11828, O11829, O11830, O11831, O11832, O11833, O11834, O11835, O11836, O11837, O11838, O11839, O11840, O11841, O11842, O11843, O11844, O11845, O11846, O11847, O11848, O11849, O11850, O11851, O11852, O11853, O11854, O11855, O11856, O11857, O11858, O11859, O11860, O11861, O11862, O11863, O11864, O11865, O11866, O11867, O11868, O11869, O11870, O11871, O11872, O11873, O11874, O11875, O11876, O11877, O11878, O11879, O11880, O11881, O11882, O11883, O11884, O11885, O11886, O11887, O11888, O11889, O11890, O11891, O11892, O11893, O11894, O11895, O11896, O11897, O11898, O11899, O11900, O11901, O11902, O11903, O11904, O11905, O11906, O11907, O11908, O11909, O11910, O11911, O11912, O11913, O11914, O11915, O11916, O11917, O11918, O11919, O11920, O11921, O11922, O11923, O11924, O11925, O11926, O11927, O11928, O11929, O11930, O11931, O11932, O11933, O11934, O11935, O11936, O11937, O11938, O11939, O11940, O11941, O11942, O11943, O11944, O11945, O11946, O11947, O11948, O11949, O11950, O11951, O11952, O11953, O11954, O11955, O11956, O11957, O11958, O11959, O11960, O11961, O11962, O11963, O11964, O11965, O11966, O11967, O11968, O11969, O11970, O11971, O11972, O11973, O11974, O11975, O11976, O11977, O11978, O11979, O11980, O11981, O11982, O11983, O11984, O11985, O11986, O11987, O11988, O11989, O11990, O11991, O11992, O11993, O11994, O11995, O11996, O11997, O11998, O11999, O12000, O12001, O12002, O12003, O12004, O12005, O12006, O12007, O12008, O12009, O12010, O12011, O12012, O12013, O12014, O12015, O12016, O12017, O12018, O12019, O12020, O12021, O12022, O12023, O12024, O12025, O12026, O12027, O12028, O12029, O12030, O12031, O12032, O12033, O12034, O12035, O12036, O12037, O12038, O12039, O12040, O12041, O12042, O12043, O12044, O12045, O12046, O12047, O12048, O12049, O12050, O12051, O12052, O12053, O12054, O12055, O12056, O12057, O12058, O12059, O12060, O12061, O12062, O12063, O12064, O12065, O12066, O12067, O12068, O12069, O12070, O12071, O12072, O12073, O12074, O12075, O12076, O12077, O12078, O12079, O12080, O12081, O12082, O12083, O12084, O12085, O12086, O12087, O12088, O12089, O12090, O12091, O12092, O12093, O12094, O12095, O12096, O12097, O12098, O12099, O12100, O12101, O12102, O12103, O12104, O12105, O12106, O12107, O12108, O12109, O12110, O12111, O12112, O12113, O12114, O12115, O12116, O12117, O12118, O12119, O12120, O12121, O12122, O12123, O12124, O12125, O12126, O12127, O12128, O12129, O12130, O12131, O12132, O12133, O12134, O12135, O12136, O12137, O12138, O12139, O12140, O12141, O12142, O12143, O12144, O12145, O12146, O12147, O12148, O12149, O12150, O12151, O12152, O12153, O12154, O12155, O12156, O12157, O12158, O12159, O12160, O12161, O12162, O12163, O12164, O12165, O12166, O12167, O12168, O12169, O12170, O12171, O12172, O12173, O12174, O12175, O12176, O12177, O12178, O12179, O12180, O12181, O12182, O12183, O12184, O12185, O12186, O12187, O12188, O12189, O12190, O12191, O12192, O12193, O12194, O12195, O12196, O12197, O12198, O12199, O12200, O12201, O12202, O12203, O12204, O12205, O12206, O12207, O12208, O12209, O12210, O12211, O12212, O12213, O12214, O12215, O12216, O12217, O12218, O12219, O12220, O12221, O12222, O12223, O12224, O12225, O12226, O12227, O12228, O12229, O12230, O12231, O12232, O12233, O12234, O12235, O12236, O12237, O12238, O12239, O12240, O12241, O12242, O12243, O12244, O12245, O12246, O12247, O12248, O12249, O12250, O12251, O12252, O12253, O12254, O12255, O12256, O12257, O12258, O12259, O12260, O12261, O12262, O12263, O12264, O12265, O12266, O12267, O12268, O12269, O12270, O12271, O12272, O12273, O12274, O12275, O12276, O12277, O12278, O12279, O12280, O12281, O12282, O12283, O12284, O12285, O12286, O12287, O12288, O12289, O12290, O12291, O12292, O12293, O12294, O12295, O12296, O12297, O12298, O12299, O12300, O12301, O12302, O12303, O12304, O12305, O12306, O12307, O12308, O12309, O12310, O12311, O12312, O12313, O12314, O12315, O12316, O12317, O12318, O12319, O12320, O12321, O12322, O12323, O12324, O12325, O12326, O12327, O12328, O12329, O12330, O12331, O12332, O12333, O12334, O12335, O12336, O12337, O12338, O12339, O12340, O12341, O12342, O12343, O12344, O12345, O12346, O12347, O12348, O12349, O12350, O12351, O12352, O12353, O12354, O12355, O12356, O12357, O12358, O12359, O12360, O12361, O12362, O12363, O12364, O12365, O12366, O12367, O12368, O12369, O12370, O12371, O12372, O12373, O12374, O12375, O12376, O12377, O12378, O12379, O12380, O12381, O12382, O12383, O12384, O12385, O12386, O12387, O12388, O12389, O12390, O12391, O12392, O12393, O12394, O12395, O12396, O12397, O12398, O12399, O12400, O12401, O12402, O12403, O12404, O12405, O12406, O12407, O12408, O12409, O12410, O12411, O12412, O12413, O12414, O12415, O12416, O12417, O12418, O12419, O12420, O12421, O12422, O12423, O12424, O12425, O12426, O12427, O12428, O12429, O12430, O12431, O12432, O12433, O12434, O12435, O12436, O12437, O12438, O12439, O12440, O12441, O12442, O12443, O12444, O12445, O12446, O12447, O12448, O12449, O12450, O12451, O12452, O12453, O12454, O12455, O12456, O12457, O12458, O12459, O12460, O12461, O12462, O12463, O12464, O12465, O12466, O12467, O12468, O12469, O12470, O12471, O12472, O12473, O12474, O12475, O12476, O12477, O12478, O12479, O12480, O12481, O12482, O12483, O12484, O12485, O12486, O12487, O12488, O12489, O12490, O12491, O12492, O12493, O12494, O12495, O12496, O12497, O12498, O12499, O12500, O12501, O12502, O12503, O12504, O12505, O12506, O12507, O12508, O12509, O12510, O12511, O12512, O12513, O12514, O12515, O12516, O12517, O12518, O12519, O12520, O12521, O12522, O12523, O12524, O12525, O12526, O12527, O12528, O12529, O12530, O12531, O12532, O12533, O12534, O12535, O12536, O12537, O12538, O12539, O12540, O12541, O12542, O12543, O12544, O12545, O12546, O12547, O12548, O12549, O12550, O12551, O12552, O12553, O12554, O12555, O12556, O12557, O12558, O12559, O12560, O12561, O12562, O12563, O12564, O12565, O12566, O12567, O12568, O12569, O12570, O12571, O12572, O12573, O12574, O12575, O12576, O12577, O12578, O12579, O12580, O12581, O12582, O12583, O12584, O12585, O12586, O12587, O12588, O12589, O12590, O12591, O12592, O12593, O12594, O12595, O12596, O12597, O12598, O12599, O12600, O12601, O12602, O12603, O12604, O12605, O12606, O12607, O12608, O12609, O12610, O12611, O12612, O12613, O12614, O12615, O12616, O12617, O12618, O12619, O12620, O12621, O12622, O12623, O12624, O12625, O12626, O12627, O12628, O12629, O12630, O12631, O12632, O12633, O12634, O12635, O12636, O12637, O12638, O12639, O12640, O12641, O12642, O12643, O12644, O12645, O12646, O12647, O12648, O12649, O12650, O12651, O12652, O12653, O12654, O12655, O12656, O12657, O12658, O12659, O12660, O12661, O12662, O12663, O12664, O12665, O12666, O12667, O12668, O12669, O12670, O12671, O12672, O12673, O12674, O12675, O12676, O12677, O12678, O12679, O12680, O12681, O12682, O12683, O12684, O12685, O12686, O12687, O12688, O12689, O12690, O12691, O12692, O12693, O12694, O12695, O12696, O12697, O12698, O12699, O12700, O12701, O12702, O12703, O12704, O12705, O12706, O12707, O12708, O12709, O12710, O12711, O12712, O12713, O12714, O12715, O12716, O12717, O12718, O12719, O12720, O12721, O12722, O12723, O12724, O12725, O12726, O12727, O12728, O12729, O12730, O12731, O12732, O12733, O12734, O12735, O12736, O12737, O12738, O12739, O12740, O12741, O12742, O12743, O12744, O12745, O12746, O12747, O12748, O12749, O12750, O12751, O12752, O12753, O12754, O12755, O12756, O12757, O12758, O12759, O12760, O12761, O12762, O12763, O12764, O12765, O12766, O12767, O12768, O12769, O12770, O12771, O12772, O12773, O12774, O12775, O12776, O12777, O12778, O12779, O12780, O12781, O12782, O12783, O12784, O12785, O12786, O12787, O12788, O12789, O12790, O12791, O12792, O12793, O12794, O12795, O12796, O12797, O12798, O12799, O12800, O12801, O12802, O12803, O12804, O12805, O12806, O12807, O12808, O12809, O12810, O12811, O12812, O12813, O12814, O12815, O12816, O12817, O12818, O12819, O12820, O12821, O12822, O12823, O12824, O12825, O12826, O12827, O12828, O12829, O12830, O12831, O12832, O12833, O12834, O12835, O12836, O12837, O12838, O12839, O12840, O12841, O12842, O12843, O12844, O12845, O12846, O12847, O12848, O12849, O12850, O12851, O12852, O12853, O12854, O12855, O12856, O12857, O12858, O12859, O12860, O12861, O12862, O12863, O12864, O12865, O12866, O12867, O12868, O12869, O12870, O12871, O12872, O12873, O12874, O12875, O12876, O12877, O12878, O12879, O12880, O12881, O12882, O12883, O12884, O12885, O12886, O12887, O12888, O12889, O12890, O12891, O12892, O12893, O12894, O12895, O12896, O12897, O12898, O12899, O12900, O12901, O12902, O12903, O12904, O12905, O12906, O12907, O12908, O12909, O12910, O12911, O12912, O12913, O12914, O12915, O12916, O12917, O12918, O12919, O12920, O12921, O12922, O12923, O12924, O12925, O12926, O12927, O12928, O12929, O12930, O12931, O12932, O12933, O12934, O12935, O12936, O12937, O12938, O12939, O12940, O12941, O12942, O12943, O12944, O12945, O12946, O12947, O12948, O12949, O12950, O12951, O12952, O12953, O12954, O12955, O12956, O12957, O12958, O12959, O12960, O12961, O12962, O12963, O12964, O12965, O12966, O12967, O12968, O12969, O12970, O12971, O12972, O12973, O12974, O12975, O12976, O12977, O12978, O12979, O12980, O12981, O12982, O12983, O12984, O12985, O12986, O12987, O12988, O12989, O12990, O12991, O12992, O12993, O12994, O12995, O12996, O12997, O12998, O12999, O13000, O13001, O13002, O13003, O13004, O13005, O13006, O13007, O13008, O13009, O13010, O13011, O13012, O13013, O13014, O13015, O13016, O13017, O13018, O13019, O13020, O13021, O13022, O13023, O13024, O13025, O13026, O13027, O13028, O13029, O13030, O13031, O13032, O13033, O13034, O13035, O13036, O13037, O13038, O13039, O13040, O13041, O13042, O13043, O13044, O13045, O13046, O13047, O13048, O13049, O13050, O13051, O13052, O13053, O13054, O13055, O13056, O13057, O13058, O13059, O13060, O13061, O13062, O13063, O13064, O13065, O13066, O13067, O13068, O13069, O13070, O13071, O13072, O13073, O13074, O13075, O13076, O13077, O13078, O13079, O13080, O13081, O13082, O13083, O13084, O13085, O13086, O13087, O13088, O13089, O13090, O13091, O13092, O13093, O13094, O13095, O13096, O13097, O13098, O13099, O13100, O13101, O13102, O13103, O13104, O13105, O13106, O13107, O13108, O13109, O13110, O13111, O13112, O13113, O13114, O13115, O13116, O13117, O13118, O13119, O13120, O13121, O13122, O13123, O13124, O13125, O13126, O13127, O13128, O13129, O13130, O13131, O13132, O13133, O13134, O13135, O13136, O13137, O13138, O13139, O13140, O13141, O13142, O13143, O13144, O13145, O13146, O13147, O13148, O13149, O13150, O13151, O13152, O13153, O13154, O13155, O13156, O13157, O13158, O13159, O13160, O13161, O13162, O13163, O13164, O13165, O13166, O13167, O13168, O13169, O13170, O13171, O13172, O13173, O13174, O13175, O13176, O13177, O13178, O13179, O13180, O13181, O13182, O13183, O13184, O13185, O13186, O13187, O13188, O13189, O13190, O13191, O13192, O13193, O13194, O13195, O13196, O13197, O13198, O13199, O13200, O13201, O13202, O13203, O13204, O13205, O13206, O13207, O13208, O13209, O13210, O13211, O13212, O13213, O13214, O13215, O13216, O13217, O13218, O13219, O13220, O13221, O13222, O13223, O13224, O13225, O13226, O13227, O13228, O13229, O13230, O13231, O13232, O13233, O13234, O13235, O13236, O13237, O13238, O13239, O13240, O13241, O13242, O13243, O13244, O13245, O13246, O13247, O13248, O13249, O13250, O13251, O13252, O13253, O13254, O13255, O13256, O13257, O13258, O13259, O13260, O13261, O13262, O13263, O13264, O13265, O13266, O13267, O13268, O13269, O13270, O13271, O13272, O13273, O13274, O13275, O13276, O13277, O13278, O13279, O13280, O13281, O13282, O13283, O13284, O13285, O13286, O13287, O13288, O13289, O13290, O13291, O13292, O13293, O13294, O13295, O13296, O13297, O13298, O13299, O13300, O13301, O13302, O13303, O13304, O13305, O13306, O13307, O13308, O13309, O13310, O13311, O13312, O13313, O13314, O13315, O13316, O13317, O13318, O13319, O13320, O13321, O13322, O13323, O13324, O13325, O13326, O13327, O13328, O13329, O13330, O13331, O13332, O13333, O13334, O13335, O13336, O13337, O13338, O13339, O13340, O13341, O13342, O13343, O13344, O13345, O13346, O13347, O13348, O13349, O13350, O13351, O13352, O13353, O13354, O13355, O13356, O13357, O13358, O13359, O13360, O13361, O13362, O13363, O13364, O13365, O13366, O13367, O13368, O13369, O13370, O13371, O13372, O13373, O13374, O13375, O13376, O13377, O13378, O13379, O13380, O13381, O13382, O13383, O13384, O13385, O13386, O13387, O13388, O13389, O13390, O13391, O13392, O13393, O13394, O13395, O13396, O13397, O13398, O13399, O13400, O13401, O13402, O13403, O13404, O13405, O13406, O13407, O13408, O13409, O13410, O13411, O13412, O13413, O13414, O13415, O13416, O13417, O13418, O13419, O13420, O13421, O13422, O13423, O13424, O13425, O13426, O13427, O13428, O13429, O13430, O13431, O13432, O13433, O13434, O13435, O13436, O13437, O13438, O13439, O13440, O13441, O13442, O13443, O13444, O13445, O13446, O13447, O13448, O13449, O13450, O13451, O13452, O13453, O13454, O13455, O13456, O13457, O13458, O13459, O13460, O13461, O13462, O13463, O13464, O13465, O13466, O13467, O13468, O13469, O13470, O13471, O13472, O13473, O13474, O13475, O13476, O13477, O13478, O13479, O13480, O13481, O13482, O13483, O13484, O13485, O13486, O13487, O13488, O13489, O13490, O13491, O13492, O13493, O13494, O13495, O13496, O13497, O13498, O13499, O13500, O13501, O13502, O13503, O13504, O13505, O13506, O13507, O13508, O13509, O13510, O13511, O13512, O13513, O13514, O13515, O13516, O13517, O13518, O13519, O13520, O13521, O13522, O13523, O13524, O13525, O13526, O13527, O13528, O13529, O13530, O13531, O13532, O13533, O13534, O13535, O13536, O13537, O13538, O13539, O13540, O13541, O13542, O13543, O13544, O13545, O13546, O13547, O13548, O13549, O13550, O13551, O13552, O13553, O13554, O13555, O13556, O13557, O13558, O13559, O13560, O13561, O13562, O13563, O13564, O13565, O13566, O13567, O13568, O13569, O13570, O13571, O13572, O13573, O13574, O13575, O13576, O13577, O13578, O13579, O13580, O13581, O13582, O13583, O13584, O13585, O13586, O13587, O13588, O13589, O13590, O13591, O13592, O13593, O13594, O13595, O13596, O13597, O13598, O13599, O13600, O13601, O13602, O13603, O13604, O13605, O13606, O13607, O13608, O13609, O13610, O13611, O13612, O13613, O13614, O13615, O13616, O13617, O13618, O13619, O13620, O13621, O13622, O13623, O13624, O13625, O13626, O13627, O13628, O13629, O13630, O13631, O13632, O13633, O13634, O13635, O13636, O13637, O13638, O13639, O13640, O13641, O13642, O13643, O13644, O13645, O13646, O13647, O13648, O13649, O13650, O13651, O13652, O13653, O13654, O13655, O13656, O13657, O13658, O13659, O13660, O13661, O13662, O13663, O13664, O13665, O13666, O13667, O13668, O13669, O13670, O13671, O13672, O13673, O13674, O13675, O13676, O13677, O13678, O13679, O13680, O13681, O13682, O13683, O13684, O13685, O13686, O13687, O13688, O13689, O13690, O13691, O13692, O13693, O13694, O13695, O13696, O13697, O13698, O13699, O13700, O13701, O13702, O13703, O13704, O13705, O13706, O13707, O13708, O13709, O13710, O13711, O13712, O13713, O13714, O13715, O13716, O13717, O13718, O13719, O13720, O13721, O13722, O13723, O13724, O13725, O13726, O13727, O13728, O13729, O13730, O13731, O13732, O13733, O13734, O13735, O13736, O13737, O13738, O13739, O13740, O13741, O13742, O13743, O13744, O13745, O13746, O13747, O13748, O13749, O13750, O13751, O13752, O13753, O13754, O13755, O13756, O13757, O13758, O13759, O13760, O13761, O13762, O13763, O13764, O13765, O13766, O13767, O13768, O13769, O13770, O13771, O13772, O13773, O13774, O13775, O13776, O13777, O13778, O13779, O13780, O13781, O13782, O13783, O13784, O13785, O13786, O13787, O13788, O13789, O13790, O13791, O13792, O13793, O13794, O13795, O13796, O13797, O13798, O13799, O13800, O13801, O13802, O13803, O13804, O13805, O13806, O13807, O13808, O13809, O13810, O13811, O13812, O13813, O13814, O13815, O13816, O13817, O13818, O13819, O13820, O13821, O13822, O13823, O13824, O13825, O13826, O13827, O13828, O13829, O13830, O13831, O13832, O13833, O13834, O13835, O13836, O13837, O13838, O13839, O13840, O13841, O13842, O13843, O13844, O13845, O13846, O13847, O13848, O13849, O13850, O13851, O13852, O13853, O13854, O13855, O13856, O13857, O13858, O13859, O13860, O13861, O13862, O13863, O13864, O13865, O13866, O13867, O13868, O13869, O13870, O13871, O13872, O13873, O13874, O13875, O13876, O13877, O13878, O13879, O13880, O13881, O13882, O13883, O13884, O13885, O13886, O13887, O13888, O13889, O13890, O13891, O13892, O13893, O13894, O13895, O13896, O13897, O13898, O13899, O13900, O13901, O13902, O13903, O13904, O13905, O13906, O13907, O13908, O13909, O13910, O13911, O13912, O13913, O13914, O13915, O13916, O13917, O13918, O13919, O13920, O13921, O13922, O13923, O13924, O13925, O13926, O13927, O13928, O13929, O13930, O13931, O13932, O13933, O13934, O13935, O13936, O13937, O13938, O13939, O13940, O13941, O13942, O13943, O13944, O13945, O13946, O13947, O13948, O13949, O13950, O13951, O13952, O13953, O13954, O13955, O13956, O13957, O13958, O13959, O13960, O13961, O13962, O13963, O13964, O13965, O13966, O13967, O13968, O13969, O13970, O13971, O13972, O13973, O13974, O13975, O13976, O13977, O13978, O13979, O13980, O13981, O13982, O13983, O13984, O13985, O13986, O13987, O13988, O13989, O13990, O13991, O13992, O13993, O13994, O13995, O13996, O13997, O13998, O13999, O14000, O14001, O14002, O14003, O14004, O14005, O14006, O14007, O14008, O14009, O14010, O14011, O14012, O14013, O14014, O14015, O14016, O14017, O14018, O14019, O14020, O14021, O14022, O14023, O14024, O14025, O14026, O14027, O14028, O14029, O14030, O14031, O14032, O14033, O14034, O14035, O14036, O14037, O14038, O14039, O14040, O14041, O14042, O14043, O14044, O14045, O14046, O14047, O14048, O14049, O14050, O14051, O14052, O14053, O14054, O14055, O14056, O14057, O14058, O14059, O14060, O14061, O14062, O14063, O14064, O14065, O14066, O14067, O14068, O14069, O14070, O14071, O14072, O14073, O14074, O14075, O14076, O14077, O14078, O14079, O14080, O14081, O14082, O14083, O14084, O14085, O14086, O14087, O14088, O14089, O14090, O14091, O14092, O14093, O14094, O14095, O14096, O14097, O14098, O14099, O14100, O14101, O14102, O14103, O14104, O14105, O14106, O14107, O14108, O14109, O14110, O14111, O14112, O14113, O14114, O14115, O14116, O14117, O14118, O14119, O14120, O14121, O14122, O14123, O14124, O14125, O14126, O14127, O14128, O14129, O14130, O14131, O14132, O14133, O14134, O14135, O14136, O14137, O14138, O14139, O14140, O14141, O14142, O14143, O14144, O14145, O14146, O14147, O14148, O14149, O14150, O14151, O14152, O14153, O14154, O14155, O14156, O14157, O14158, O14159, O14160, O14161, O14162, O14163, O14164, O14165, O14166, O14167, O14168, O14169, O14170, O14171, O14172, O14173, O14174, O14175, O14176, O14177, O14178, O14179, O14180, O14181, O14182, O14183, O14184, O14185, O14186, O14187, O14188, O14189, O14190, O14191, O14192, O14193, O14194, O14195, O14196, O14197, O14198, O14199, O14200, O14201, O14202, O14203, O14204, O14205, O14206, O14207, O14208, O14209, O14210, O14211, O14212, O14213, O14214, O14215, O14216, O14217, O14218, O14219, O14220, O14221, O14222, O14223, O14224, O14225, O14226, O14227, O14228, O14229, O14230, O14231, O14232, O14233, O14234, O14235, O14236, O14237, O14238, O14239, O14240, O14241, O14242, O14243, O14244, O14245, O14246, O14247, O14248, O14249, O14250, O14251, O14252, O14253, O14254, O14255, O14256, O14257, O14258, O14259, O14260, O14261, O14262, O14263, O14264, O14265, O14266, O14267, O14268, O14269, O14270, O14271, O14272, O14273, O14274, O14275, O14276, O14277, O14278, O14279, O14280, O14281, O14282, O14283, O14284, O14285, O14286, O14287, O14288, O14289, O14290, O14291, O14292, O14293, O14294, O14295, O14296, O14297, O14298, O14299, O14300, O14301, O14302, O14303, O14304, O14305, O14306, O14307, O14308, O14309, O14310, O14311, O14312, O14313, O14314, O14315, O14316, O14317, O14318, O14319, O14320, O14321, O14322, O14323, O14324, O14325, O14326, O14327, O14328, O14329, O14330, O14331, O14332, O14333, O14334, O14335, O14336, O14337, O14338, O14339, O14340, O14341, O14342, O14343, O14344, O14345, O14346, O14347, O14348, O14349, O14350, O14351, O14352, O14353, O14354, O14355, O14356, O14357, O14358, O14359, O14360, O14361, O14362, O14363, O14364, O14365, O14366, O14367, O14368, O14369, O14370, O14371, O14372, O14373, O14374, O14375, O14376, O14377, O14378, O14379, O14380, O14381, O14382, O14383, O14384, O14385, O14386, O14387, O14388, O14389, O14390, O14391, O14392, O14393, O14394, O14395, O14396, O14397, O14398, O14399, O14400, O14401, O14402, O14403, O14404, O14405, O14406, O14407, O14408, O14409, O14410, O14411, O14412, O14413, O14414, O14415, O14416, O14417, O14418, O14419, O14420, O14421, O14422, O14423, O14424, O14425, O14426, O14427, O14428, O14429, O14430, O14431, O14432, O14433, O14434, O14435, O14436, O14437, O14438, O14439, O14440, O14441, O14442, O14443, O14444, O14445, O14446, O14447, O14448, O14449, O14450, O14451, O14452, O14453, O14454, O14455, O14456, O14457, O14458, O14459, O14460, O14461, O14462, O14463, O14464, O14465, O14466, O14467, O14468, O14469, O14470, O14471, O14472, O14473, O14474, O14475, O14476, O14477, O14478, O14479, O14480, O14481, O14482, O14483, O14484, O14485, O14486, O14487, O14488, O14489, O14490, O14491, O14492, O14493, O14494, O14495, O14496, O14497, O14498, O14499, O14500, O14501, O14502, O14503, O14504, O14505, O14506, O14507, O14508, O14509, O14510, O14511, O14512, O14513, O14514, O14515, O14516, O14517, O14518, O14519, O14520, O14521, O14522, O14523, O14524, O14525, O14526, O14527, O14528, O14529, O14530, O14531, O14532, O14533, O14534, O14535, O14536, O14537, O14538, O14539, O14540, O14541, O14542, O14543, O14544, O14545, O14546, O14547, O14548, O14549, O14550, O14551, O14552, O14553, O14554, O14555, O14556, O14557, O14558, O14559, O14560, O14561, O14562, O14563, O14564, O14565, O14566, O14567, O14568, O14569, O14570, O14571, O14572, O14573, O14574, O14575, O14576, O14577, O14578, O14579, O14580, O14581, O14582, O14583, O14584, O14585, O14586, O14587, O14588, O14589, O14590, O14591, O14592, O14593, O14594, O14595, O14596, O14597, O14598, O14599, O14600, O14601, O14602, O14603, O14604, O14605, O14606, O14607, O14608, O14609, O14610, O14611, O14612, O14613, O14614, O14615, O14616, O14617, O14618, O14619, O14620, O14621, O14622, O14623, O14624, O14625, O14626, O14627, O14628, O14629, O14630, O14631, O14632, O14633, O14634, O14635, O14636, O14637, O14638, O14639, O14640, O14641, O14642, O14643, O14644, O14645, O14646, O14647, O14648, O14649, O14650, O14651, O14652, O14653, O14654, O14655, O14656, O14657, O14658, O14659, O14660, O14661, O14662, O14663, O14664, O14665, O14666, O14667, O14668, O14669, O14670, O14671, O14672, O14673, O14674, O14675, O14676, O14677, O14678, O14679, O14680, O14681, O14682, O14683, O14684, O14685, O14686, O14687, O14688, O14689, O14690, O14691, O14692, O14693, O14694, O14695, O14696, O14697, O14698, O14699, O14700, O14701, O14702, O14703, O14704, O14705, O14706, O14707, O14708, O14709, O14710, O14711, O14712, O14713, O14714, O14715, O14716, O14717, O14718, O14719, O14720, O14721, O14722, O14723, O14724, O14725, O14726, O14727, O14728, O14729, O14730, O14731, O14732, O14733, O14734, O14735, O14736, O14737, O14738, O14739, O14740, O14741, O14742, O14743, O14744, O14745, O14746, O14747, O14748, O14749, O14750, O14751, O14752, O14753, O14754, O14755, O14756, O14757, O14758, O14759, O14760, O14761, O14762, O14763, O14764, O14765, O14766, O14767, O14768, O14769, O14770, O14771, O14772, O14773, O14774, O14775, O14776, O14777, O14778, O14779, O14780, O14781, O14782, O14783, O14784, O14785, O14786, O14787, O14788, O14789, O14790, O14791, O14792, O14793, O14794, O14795, O14796, O14797, O14798, O14799, O14800, O14801, O14802, O14803, O14804, O14805, O14806, O14807, O14808, O14809, O14810, O14811, O14812, O14813, O14814, O14815, O14816, O14817, O14818, O14819, O14820, O14821, O14822, O14823, O14824, O14825, O14826, O14827, O14828, O14829, O14830, O14831, O14832, O14833, O14834, O14835, O14836, O14837, O14838, O14839, O14840, O14841, O14842, O14843, O14844, O14845, O14846, O14847, O14848, O14849, O14850, O14851, O14852, O14853, O14854, O14855, O14856, O14857, O14858, O14859, O14860, O14861, O14862, O14863, O14864, O14865, O14866, O14867, O14868, O14869, O14870, O14871, O14872, O14873, O14874, O14875, O14876, O14877, O14878, O14879, O14880, O14881, O14882, O14883, O14884, O14885, O14886, O14887, O14888, O14889, O14890, O14891, O14892, O14893, O14894, O14895, O14896, O14897, O14898, O14899, O14900, O14901, O14902, O14903, O14904, O14905, O14906, O14907, O14908, O14909, O14910, O14911, O14912, O14913, O14914, O14915, O14916, O14917, O14918, O14919, O14920, O14921, O14922, O14923, O14924, O14925, O14926, O14927, O14928, O14929, O14930, O14931, O14932, O14933, O14934, O14935, O14936, O14937, O14938, O14939, O14940, O14941, O14942, O14943, O14944, O14945, O14946, O14947, O14948, O14949, O14950, O14951, O14952, O14953, O14954, O14955, O14956, O14957, O14958, O14959, O14960, O14961, O14962, O14963, O14964, O14965, O14966, O14967, O14968, O14969, O14970, O14971, O14972, O14973, O14974, O14975, O14976, O14977, O14978, O14979, O14980, O14981, O14982, O14983, O14984, O14985, O14986, O14987, O14988, O14989, O14990, O14991, O14992, O14993, O14994, O14995, O14996, O14997, O14998, O14999, O15000, O15001, O15002, O15003, O15004, O15005, O15006, O15007, O15008, O15009, O15010, O15011, O15012, O15013, O15014, O15015, O15016, O15017, O15018, O15019, O15020, O15021, O15022, O15023, O15024, O15025, O15026, O15027, O15028, O15029, O15030, O15031, O15032, O15033, O15034, O15035, O15036, O15037, O15038, O15039, O15040, O15041, O15042, O15043, O15044, O15045, O15046, O15047, O15048, O15049, O15050, O15051, O15052, O15053, O15054, O15055, O15056, O15057, O15058, O15059, O15060, O15061, O15062, O15063, O15064, O15065, O15066, O15067, O15068, O15069, O15070, O15071, O15072, O15073, O15074, O15075, O15076, O15077, O15078, O15079, O15080, O15081, O15082, O15083, O15084, O15085, O15086, O15087, O15088, O15089, O15090, O15091, O15092, O15093, O15094, O15095, O15096, O15097, O15098, O15099, O15100, O15101, O15102, O15103, O15104, O15105, O15106, O15107, O15108, O15109, O15110, O15111, O15112, O15113, O15114, O15115, O15116, O15117, O15118, O15119, O15120, O15121, O15122, O15123, O15124, O15125, O15126, O15127, O15128, O15129, O15130, O15131, O15132, O15133, O15134, O15135, O15136, O15137, O15138, O15139, O15140, O15141, O15142, O15143, O15144, O15145, O15146, O15147, O15148, O15149, O15150, O15151, O15152, O15153, O15154, O15155, O15156, O15157, O15158, O15159, O15160, O15161, O15162, O15163, O15164, O15165, O15166, O15167, O15168, O15169, O15170, O15171, O15172, O15173, O15174, O15175, O15176, O15177, O15178, O15179, O15180, O15181, O15182, O15183, O15184, O15185, O15186, O15187, O15188, O15189, O15190, O15191, O15192, O15193, O15194, O15195, O15196, O15197, O15198, O15199, O15200, O15201, O15202, O15203, O15204, O15205, O15206, O15207, O15208, O15209, O15210, O15211, O15212, O15213, O15214, O15215, O15216, O15217, O15218, O15219, O15220, O15221, O15222, O15223, O15224, O15225, O15226, O15227, O15228, O15229, O15230, O15231, O15232, O15233, O15234, O15235, O15236, O15237, O15238, O15239, O15240, O15241, O15242, O15243, O15244, O15245, O15246, O15247, O15248, O15249, O15250, O15251, O15252, O15253, O15254, O15255, O15256, O15257, O15258, O15259, O15260, O15261, O15262, O15263, O15264, O15265, O15266, O15267, O15268, O15269, O15270, O15271, O15272, O15273, O15274, O15275, O15276, O15277, O15278, O15279, O15280, O15281, O15282, O15283, O15284, O15285, O15286, O15287, O15288, O15289, O15290, O15291, O15292, O15293, O15294, O15295, O15296, O15297, O15298, O15299, O15300, O15301, O15302, O15303, O15304, O15305, O15306, O15307, O15308, O15309, O15310, O15311, O15312, O15313, O15314, O15315, O15316, O15317, O15318, O15319, O15320, O15321, O15322, O15323, O15324, O15325, O15326, O15327, O15328, O15329, O15330, O15331, O15332, O15333, O15334, O15335, O15336, O15337, O15338, O15339, O15340, O15341, O15342, O15343, O15344, O15345, O15346, O15347, O15348, O15349, O15350, O15351, O15352, O15353, O15354, O15355, O15356, O15357, O15358, O15359, O15360, O15361, O15362, O15363, O15364, O15365, O15366, O15367, O15368, O15369, O15370, O15371, O15372, O15373, O15374, O15375, O15376, O15377, O15378, O15379, O15380, O15381, O15382, O15383, O15384, O15385, O15386, O15387, O15388, O15389, O15390, O15391, O15392, O15393, O15394, O15395, O15396, O15397, O15398, O15399, O15400, O15401, O15402, O15403, O15404, O15405, O15406, O15407, O15408, O15409, O15410, O15411, O15412, O15413, O15414, O15415, O15416, O15417, O15418, O15419, O15420, O15421, O15422, O15423, O15424, O15425, O15426, O15427, O15428, O15429, O15430, O15431, O15432, O15433, O15434, O15435, O15436, O15437, O15438, O15439, O15440, O15441, O15442, O15443, O15444, O15445, O15446, O15447, O15448, O15449, O15450, O15451, O15452, O15453, O15454, O15455, O15456, O15457, O15458, O15459, O15460, O15461, O15462, O15463, O15464, O15465, O15466, O15467, O15468, O15469, O15470, O15471, O15472, O15473, O15474, O15475, O15476, O15477, O15478, O15479, O15480, O15481, O15482, O15483, O15484, O15485, O15486, O15487, O15488, O15489, O15490, O15491, O15492, O15493, O15494, O15495, O15496, O15497, O15498, O15499, O15500, O15501, O15502, O15503, O15504, O15505, O15506, O15507, O15508, O15509, O15510, O15511, O15512, O15513, O15514, O15515, O15516, O15517, O15518, O15519, O15520, O15521, O15522, O15523, O15524, O15525, O15526, O15527, O15528, O15529, O15530, O15531, O15532, O15533, O15534, O15535, O15536, O15537, O15538, O15539, O15540, O15541, O15542, O15543, O15544, O15545, O15546, O15547, O15548, O15549, O15550, O15551, O15552, O15553, O15554, O15555, O15556, O15557, O15558, O15559, O15560, O15561, O15562, O15563, O15564, O15565, O15566, O15567, O15568, O15569, O15570, O15571, O15572, O15573, O15574, O15575, O15576, O15577, O15578, O15579, O15580, O15581, O15582, O15583, O15584, O15585, O15586, O15587, O15588, O15589, O15590, O15591, O15592, O15593, O15594, O15595, O15596, O15597, O15598, O15599, O15600, O15601, O15602, O15603, O15604, O15605, O15606, O15607, O15608, O15609, O15610, O15611, O15612, O15613, O15614, O15615, O15616, O15617, O15618, O15619, O15620, O15621, O15622, O15623, O15624, O15625, O15626, O15627, O15628, O15629, O15630, O15631, O15632, O15633, O15634, O15635, O15636, O15637, O15638, O15639, O15640, O15641, O15642, O15643, O15644, O15645, O15646, O15647, O15648, O15649, O15650, O15651, O15652, O15653, O15654, O15655, O15656, O15657, O15658, O15659, O15660, O15661, O15662, O15663, O15664, O15665, O15666, O15667, O15668, O15669, O15670, O15671, O15672, O15673, O15674, O15675, O15676, O15677, O15678, O15679, O15680, O15681, O15682, O15683, O15684, O15685, O15686, O15687, O15688, O15689, O15690, O15691, O15692, O15693, O15694, O15695, O15696, O15697, O15698, O15699, O15700, O15701, O15702, O15703, O15704, O15705, O15706, O15707, O15708, O15709, O15710, O15711, O15712, O15713, O15714, O15715, O15716, O15717, O15718, O15719, O15720, O15721, O15722, O15723, O15724, O15725, O15726, O15727, O15728, O15729, O15730, O15731, O15732, O15733, O15734, O15735, O15736, O15737, O15738, O15739, O15740, O15741, O15742, O15743, O15744, O15745, O15746, O15747, O15748, O15749, O15750, O15751, O15752, O15753, O15754, O15755, O15756, O15757, O15758, O15759, O15760, O15761, O15762, O15763, O15764, O15765, O15766, O15767, O15768, O15769, O15770, O15771, O15772, O15773, O15774, O15775, O15776, O15777, O15778, O15779, O15780, O15781, O15782, O15783, O15784, O15785, O15786, O15787, O15788, O15789, O15790, O15791, O15792, O15793, O15794, O15795, O15796, O15797, O15798, O15799, O15800, O15801, O15802, O15803, O15804, O15805, O15806, O15807, O15808, O15809, O15810, O15811, O15812, O15813, O15814, O15815, O15816, O15817, O15818, O15819, O15820, O15821, O15822, O15823, O15824, O15825, O15826, O15827, O15828, O15829, O15830, O15831, O15832, O15833, O15834, O15835, O15836, O15837, O15838, O15839, O15840, O15841, O15842, O15843, O15844, O15845, O15846, O15847, O15848, O15849, O15850, O15851, O15852, O15853, O15854, O15855, O15856, O15857, O15858, O15859, O15860, O15861, O15862, O15863, O15864, O15865, O15866, O15867, O15868, O15869, O15870, O15871, O15872, O15873, O15874, O15875, O15876, O15877, O15878, O15879, O15880, O15881, O15882, O15883, O15884, O15885, O15886, O15887, O15888, O15889, O15890, O15891, O15892, O15893, O15894, O15895, O15896, O15897, O15898, O15899, O15900, O15901, O15902, O15903, O15904, O15905, O15906, O15907, O15908, O15909, O15910, O15911, O15912, O15913, O15914, O15915, O15916, O15917, O15918, O15919, O15920, O15921, O15922, O15923, O15924, O15925, O15926, O15927, O15928, O15929, O15930, O15931, O15932, O15933, O15934, O15935, O15936, O15937, O15938, O15939, O15940, O15941, O15942, O15943, O15944, O15945, O15946, O15947, O15948, O15949, O15950, O15951, O15952, O15953, O15954, O15955, O15956, O15957, O15958, O15959, O15960, O15961, O15962, O15963, O15964, O15965, O15966, O15967, O15968, O15969, O15970, O15971, O15972, O15973, O15974, O15975, O15976, O15977, O15978, O15979, O15980, O15981, O15982, O15983, O15984, O15985, O15986, O15987, O15988, O15989, O15990, O15991, O15992, O15993, O15994, O15995, O15996, O15997, O15998, O15999, O16000, O16001, O16002, O16003, O16004, O16005, O16006, O16007, O16008, O16009, O16010, O16011, O16012, O16013, O16014, O16015, O16016, O16017, O16018, O16019, O16020, O16021, O16022, O16023, O16024, O16025, O16026, O16027, O16028, O16029, O16030, O16031, O16032, O16033, O16034, O16035, O16036, O16037, O16038, O16039, O16040, O16041, O16042, O16043, O16044, O16045, O16046, O16047, O16048, O16049, O16050, O16051, O16052, O16053, O16054, O16055, O16056, O16057, O16058, O16059, O16060, O16061, O16062, O16063, O16064, O16065, O16066, O16067, O16068, O16069, O16070, O16071, O16072, O16073, O16074, O16075, O16076, O16077, O16078, O16079, O16080, O16081, O16082, O16083, O16084, O16085, O16086, O16087, O16088, O16089, O16090, O16091, O16092, O16093, O16094, O16095, O16096, O16097, O16098, O16099, O16100, O16101, O16102, O16103, O16104, O16105, O16106, O16107, O16108, O16109, O16110, O16111, O16112, O16113, O16114, O16115, O16116, O16117, O16118, O16119, O16120, O16121, O16122, O16123, O16124, O16125, O16126, O16127, O16128, O16129, O16130, O16131, O16132, O16133, O16134, O16135, O16136, O16137, O16138, O16139, O16140, O16141, O16142, O16143, O16144, O16145, O16146, O16147, O16148, O16149, O16150, O16151, O16152, O16153, O16154, O16155, O16156, O16157, O16158, O16159, O16160, O16161, O16162, O16163, O16164, O16165, O16166, O16167, O16168, O16169, O16170, O16171, O16172, O16173, O16174, O16175, O16176, O16177, O16178, O16179, O16180, O16181, O16182, O16183, O16184, O16185, O16186, O16187, O16188, O16189, O16190, O16191, O16192, O16193, O16194, O16195, O16196, O16197, O16198, O16199, O16200, O16201, O16202, O16203, O16204, O16205, O16206, O16207, O16208, O16209, O16210, O16211, O16212, O16213, O16214, O16215, O16216, O16217, O16218, O16219, O16220, O16221, O16222, O16223, O16224, O16225, O16226, O16227, O16228, O16229, O16230, O16231, O16232, O16233, O16234, O16235, O16236, O16237, O16238, O16239, O16240, O16241, O16242, O16243, O16244, O16245, O16246, O16247, O16248, O16249, O16250, O16251, O16252, O16253, O16254, O16255, O16256, O16257, O16258, O16259, O16260, O16261, O16262, O16263, O16264, O16265, O16266, O16267, O16268, O16269, O16270, O16271, O16272, O16273, O16274, O16275, O16276, O16277, O16278, O16279, O16280, O16281, O16282, O16283, O16284, O16285, O16286, O16287, O16288, O16289, O16290, O16291, O16292, O16293, O16294, O16295, O16296, O16297, O16298, O16299, O16300, O16301, O16302, O16303, O16304, O16305, O16306, O16307, O16308, O16309, O16310, O16311, O16312, O16313, O16314, O16315, O16316, O16317, O16318, O16319, O16320, O16321, O16322, O16323, O16324, O16325, O16326, O16327, O16328, O16329, O16330, O16331, O16332, O16333, O16334, O16335, O16336, O16337, O16338, O16339, O16340, O16341, O16342, O16343, O16344, O16345, O16346, O16347, O16348, O16349, O16350, O16351, O16352, O16353, O16354, O16355, O16356, O16357, O16358, O16359, O16360, O16361, O16362, O16363, O16364, O16365, O16366, O16367, O16368, O16369, O16370, O16371, O16372, O16373, O16374, O16375, O16376, O16377, O16378, O16379, O16380, O16381, O16382, O16383, O16384, O16385, O16386, O16387, O16388, O16389, O16390, O16391, O16392, O16393, O16394, O16395, O16396, O16397, O16398, O16399, O16400, O16401, O16402, O16403, O16404, O16405, O16406, O16407, O16408, O16409, O16410, O16411, O16412, O16413, O16414, O16415, O16416, O16417, O16418, O16419, O16420, O16421, O16422, O16423, O16424, O16425, O16426, O16427, O16428, O16429, O16430, O16431, O16432, O16433, O16434, O16435, O16436, O16437, O16438, O16439, O16440, O16441, O16442, O16443, O16444, O16445, O16446, O16447, O16448, O16449, O16450, O16451, O16452, O16453, O16454, O16455, O16456, O16457, O16458, O16459, O16460, O16461, O16462, O16463, O16464, O16465, O16466, O16467, O16468, O16469, O16470, O16471, O16472, O16473, O16474, O16475, O16476, O16477, O16478, O16479, O16480, O16481, O16482, O16483, O16484, O16485, O16486, O16487, O16488, O16489, O16490, O16491, O16492, O16493, O16494, O16495, O16496, O16497, O16498, O16499, O16500, O16501, O16502, O16503, O16504, O16505, O16506, O16507, O16508, O16509, O16510, O16511, O16512, O16513, O16514, O16515, O16516, O16517, O16518, O16519, O16520, O16521, O16522, O16523, O16524, O16525, O16526, O16527, O16528, O16529, O16530, O16531, O16532, O16533, O16534, O16535, O16536, O16537, O16538, O16539, O16540, O16541, O16542, O16543, O16544, O16545, O16546, O16547, O16548, O16549, O16550, O16551, O16552, O16553, O16554, O16555, O16556, O16557, O16558, O16559, O16560, O16561, O16562, O16563, O16564, O16565, O16566, O16567, O16568, O16569, O16570, O16571, O16572, O16573, O16574, O16575, O16576, O16577, O16578, O16579, O16580, O16581, O16582, O16583, O16584, O16585, O16586, O16587, O16588, O16589, O16590, O16591, O16592, O16593, O16594, O16595, O16596, O16597, O16598, O16599, O16600, O16601, O16602, O16603, O16604, O16605, O16606, O16607, O16608, O16609, O16610, O16611, O16612, O16613, O16614, O16615, O16616, O16617, O16618, O16619, O16620, O16621, O16622, O16623, O16624, O16625, O16626, O16627, O16628, O16629, O16630, O16631, O16632, O16633, O16634, O16635, O16636, O16637, O16638, O16639, O16640, O16641, O16642, O16643, O16644, O16645, O16646, O16647, O16648, O16649, O16650, O16651, O16652, O16653, O16654, O16655, O16656, O16657, O16658, O16659, O16660, O16661, O16662, O16663, O16664, O16665, O16666, O16667, O16668, O16669, O16670, O16671, O16672, O16673, O16674, O16675, O16676, O16677, O16678, O16679, O16680, O16681, O16682, O16683, O16684, O16685, O16686, O16687, O16688, O16689, O16690, O16691, O16692, O16693, O16694, O16695, O16696, O16697, O16698, O16699, O16700, O16701, O16702, O16703, O16704, O16705, O16706, O16707, O16708, O16709, O16710, O16711, O16712, O16713, O16714, O16715, O16716, O16717, O16718, O16719, O16720, O16721, O16722, O16723, O16724, O16725, O16726, O16727, O16728, O16729, O16730, O16731, O16732, O16733, O16734, O16735, O16736, O16737, O16738, O16739, O16740, O16741, O16742, O16743, O16744, O16745, O16746, O16747, O16748, O16749, O16750, O16751, O16752, O16753, O16754, O16755, O16756, O16757, O16758, O16759, O16760, O16761, O16762, O16763, O16764, O16765, O16766, O16767, O16768, O16769, O16770, O16771, O16772, O16773, O16774, O16775, O16776, O16777, O16778, O16779, O16780, O16781, O16782, O16783, O16784, O16785, O16786, O16787, O16788, O16789, O16790, O16791, O16792, O16793, O16794, O16795, O16796, O16797, O16798, O16799, O16800, O16801, O16802, O16803, O16804, O16805, O16806, O16807, O16808, O16809, O16810, O16811, O16812, O16813, O16814, O16815, O16816, O16817, O16818, O16819, O16820, O16821, O16822, O16823, O16824, O16825, O16826, O16827, O16828, O16829, O16830, O16831, O16832, O16833, O16834, O16835, O16836, O16837, O16838, O16839, O16840, O16841, O16842, O16843, O16844, O16845, O16846, O16847, O16848, O16849, O16850, O16851, O16852, O16853, O16854, O16855, O16856, O16857, O16858, O16859, O16860, O16861, O16862, O16863, O16864, O16865, O16866, O16867, O16868, O16869, O16870, O16871, O16872, O16873, O16874, O16875, O16876, O16877, O16878, O16879, O16880, O16881, O16882, O16883, O16884, O16885, O16886, O16887, O16888, O16889, O16890, O16891, O16892, O16893, O16894, O16895, O16896, O16897, O16898, O16899, O16900, O16901, O16902, O16903, O16904, O16905, O16906, O16907, O16908, O16909, O16910, O16911, O16912, O16913, O16914, O16915, O16916, O16917, O16918, O16919, O16920, O16921, O16922, O16923, O16924, O16925, O16926, O16927, O16928, O16929, O16930, O16931, O16932, O16933, O16934, O16935, O16936, O16937, O16938, O16939, O16940, O16941, O16942, O16943, O16944, O16945, O16946, O16947, O16948, O16949, O16950, O16951, O16952, O16953, O16954, O16955, O16956, O16957, O16958, O16959, O16960, O16961, O16962, O16963, O16964, O16965, O16966, O16967, O16968, O16969, O16970, O16971, O16972, O16973, O16974, O16975, O16976, O16977, O16978, O16979, O16980, O16981, O16982, O16983, O16984, O16985, O16986, O16987, O16988, O16989, O16990, O16991, O16992, O16993, O16994, O16995, O16996, O16997, O16998, O16999, O17000, O17001, O17002, O17003, O17004, O17005, O17006, O17007, O17008, O17009, O17010, O17011, O17012, O17013, O17014, O17015, O17016, O17017, O17018, O17019, O17020, O17021, O17022, O17023, O17024, O17025, O17026, O17027, O17028, O17029, O17030, O17031, O17032, O17033, O17034, O17035, O17036, O17037, O17038, O17039, O17040, O17041, O17042, O17043, O17044, O17045, O17046, O17047, O17048, O17049, O17050, O17051, O17052, O17053, O17054, O17055, O17056, O17057, O17058, O17059, O17060, O17061, O17062, O17063, O17064, O17065, O17066, O17067, O17068, O17069, O17070, O17071, O17072, O17073, O17074, O17075, O17076, O17077, O17078, O17079, O17080, O17081, O17082, O17083, O17084, O17085, O17086, O17087, O17088, O17089, O17090, O17091, O17092, O17093, O17094, O17095, O17096, O17097, O17098, O17099, O17100, O17101, O17102, O17103, O17104, O17105, O17106, O17107, O17108, O17109, O17110, O17111, O17112, O17113, O17114, O17115, O17116, O17117, O17118, O17119, O17120, O17121, O17122, O17123, O17124, O17125, O17126, O17127, O17128, O17129, O17130, O17131, O17132, O17133, O17134, O17135, O17136, O17137, O17138, O17139, O17140, O17141, O17142, O17143, O17144, O17145, O17146, O17147, O17148, O17149, O17150, O17151, O17152, O17153, O17154, O17155, O17156, O17157, O17158, O17159, O17160, O17161, O17162, O17163, O17164, O17165, O17166, O17167, O17168, O17169, O17170, O17171, O17172, O17173, O17174, O17175, O17176, O17177, O17178, O17179, O17180, O17181, O17182, O17183, O17184, O17185, O17186, O17187, O17188, O17189, O17190, O17191, O17192, O17193, O17194, O17195, O17196, O17197, O17198, O17199, O17200, O17201, O17202, O17203, O17204, O17205, O17206, O17207, O17208, O17209, O17210, O17211, O17212, O17213, O17214, O17215, O17216, O17217, O17218, O17219, O17220, O17221, O17222, O17223, O17224, O17225, O17226, O17227, O17228, O17229, O17230, O17231, O17232, O17233, O17234, O17235, O17236, O17237, O17238, O17239, O17240, O17241, O17242, O17243, O17244, O17245, O17246, O17247, O17248, O17249, O17250, O17251, O17252, O17253, O17254, O17255, O17256, O17257, O17258, O17259, O17260, O17261, O17262, O17263, O17264, O17265, O17266, O17267, O17268, O17269, O17270, O17271, O17272, O17273, O17274, O17275, O17276, O17277, O17278, O17279, O17280, O17281, O17282, O17283, O17284, O17285, O17286, O17287, O17288, O17289, O17290, O17291, O17292, O17293, O17294, O17295, O17296, O17297, O17298, O17299, O17300, O17301, O17302, O17303, O17304, O17305, O17306, O17307, O17308, O17309, O17310, O17311, O17312, O17313, O17314, O17315, O17316, O17317, O17318, O17319, O17320, O17321, O17322, O17323, O17324, O17325, O17326, O17327, O17328, O17329, O17330, O17331, O17332, O17333, O17334, O17335, O17336, O17337, O17338, O17339, O17340, O17341, O17342, O17343, O17344, O17345, O17346, O17347, O17348, O17349, O17350, O17351, O17352, O17353, O17354, O17355, O17356, O17357, O17358, O17359, O17360, O17361, O17362, O17363, O17364, O17365, O17366, O17367, O17368, O17369, O17370, O17371, O17372, O17373, O17374, O17375, O17376, O17377, O17378, O17379, O17380, O17381, O17382, O17383, O17384, O17385, O17386, O17387, O17388, O17389, O17390, O17391, O17392, O17393, O17394, O17395, O17396, O17397, O17398, O17399, O17400, O17401, O17402, O17403, O17404, O17405, O17406, O17407, O17408, O17409, O17410, O17411, O17412, O17413, O17414, O17415, O17416, O17417, O17418, O17419, O17420, O17421, O17422, O17423, O17424, O17425, O17426, O17427, O17428, O17429, O17430, O17431, O17432, O17433, O17434, O17435, O17436, O17437, O17438, O17439, O17440, O17441, O17442, O17443, O17444, O17445, O17446, O17447, O17448, O17449, O17450, O17451, O17452, O17453, O17454, O17455, O17456, O17457, O17458, O17459, O17460, O17461, O17462, O17463, O17464, O17465, O17466, O17467, O17468, O17469, O17470, O17471, O17472, O17473, O17474, O17475, O17476, O17477, O17478, O17479, O17480, O17481, O17482, O17483, O17484, O17485, O17486, O17487, O17488, O17489, O17490, O17491, O17492, O17493, O17494, O17495, O17496, O17497, O17498, O17499, O17500, O17501, O17502, O17503, O17504, O17505, O17506, O17507, O17508, O17509, O17510, O17511, O17512, O17513, O17514, O17515, O17516, O17517, O17518, O17519, O17520, O17521, O17522, O17523, O17524, O17525, O17526, O17527, O17528, O17529, O17530, O17531, O17532, O17533, O17534, O17535, O17536, O17537, O17538, O17539, O17540, O17541, O17542, O17543, O17544, O17545, O17546, O17547, O17548, O17549, O17550, O17551, O17552, O17553, O17554, O17555, O17556, O17557, O17558, O17559, O17560, O17561, O17562, O17563, O17564, O17565, O17566, O17567, O17568, O17569, O17570, O17571, O17572, O17573, O17574, O17575, O17576, O17577, O17578, O17579, O17580, O17581, O17582, O17583, O17584, O17585, O17586, O17587, O17588, O17589, O17590, O17591, O17592, O17593, O17594, O17595, O17596, O17597, O17598, O17599, O17600, O17601, O17602, O17603, O17604, O17605, O17606, O17607, O17608, O17609, O17610, O17611, O17612, O17613, O17614, O17615, O17616, O17617, O17618, O17619, O17620, O17621, O17622, O17623, O17624, O17625, O17626, O17627, O17628, O17629, O17630, O17631, O17632, O17633, O17634, O17635, O17636, O17637, O17638, O17639, O17640, O17641, O17642, O17643, O17644, O17645, O17646, O17647, O17648, O17649, O17650, O17651, O17652, O17653, O17654, O17655, O17656, O17657, O17658, O17659, O17660, O17661, O17662, O17663, O17664, O17665, O17666, O17667, O17668, O17669, O17670, O17671, O17672, O17673, O17674, O17675, O17676, O17677, O17678, O17679, O17680, O17681, O17682, O17683, O17684, O17685, O17686, O17687, O17688, O17689, O17690, O17691, O17692, O17693, O17694, O17695, O17696, O17697, O17698, O17699, O17700, O17701, O17702, O17703, O17704, O17705, O17706, O17707, O17708, O17709, O17710, O17711, O17712, O17713, O17714, O17715, O17716, O17717, O17718, O17719, O17720, O17721, O17722, O17723, O17724, O17725, O17726, O17727, O17728, O17729, O17730, O17731, O17732, O17733, O17734, O17735, O17736, O17737, O17738, O17739, O17740, O17741, O17742, O17743, O17744, O17745, O17746, O17747, O17748, O17749, O17750, O17751, O17752, O17753, O17754, O17755, O17756, O17757, O17758, O17759, O17760, O17761, O17762, O17763, O17764, O17765, O17766, O17767, O17768, O17769, O17770, O17771, O17772, O17773, O17774, O17775, O17776, O17777, O17778, O17779, O17780, O17781, O17782, O17783, O17784, O17785, O17786, O17787, O17788, O17789, O17790, O17791, O17792, O17793, O17794, O17795, O17796, O17797, O17798, O17799, O17800, O17801, O17802, O17803, O17804, O17805, O17806, O17807, O17808, O17809, O17810, O17811, O17812, O17813, O17814, O17815, O17816, O17817, O17818, O17819, O17820, O17821, O17822, O17823, O17824, O17825, O17826, O17827, O17828, O17829, O17830, O17831, O17832, O17833, O17834, O17835, O17836, O17837, O17838, O17839, O17840, O17841, O17842, O17843, O17844, O17845, O17846, O17847, O17848, O17849, O17850, O17851, O17852, O17853, O17854, O17855, O17856, O17857, O17858, O17859, O17860, O17861, O17862, O17863, O17864, O17865, O17866, O17867, O17868, O17869, O17870, O17871, O17872, O17873, O17874, O17875, O17876, O17877, O17878, O17879, O17880, O17881, O17882, O17883, O17884, O17885, O17886, O17887, O17888, O17889, O17890, O17891, O17892, O17893, O17894, O17895, O17896, O17897, O17898, O17899, O17900, O17901, O17902, O17903, O17904, O17905, O17906, O17907, O17908, O17909, O17910, O17911, O17912, O17913, O17914, O17915, O17916, O17917, O17918, O17919, O17920, O17921, O17922, O17923, O17924, O17925, O17926, O17927, O17928, O17929, O17930, O17931, O17932, O17933, O17934, O17935, O17936, O17937, O17938, O17939, O17940, O17941, O17942, O17943, O17944, O17945, O17946, O17947, O17948, O17949, O17950, O17951, O17952, O17953, O17954, O17955, O17956, O17957, O17958, O17959, O17960, O17961, O17962, O17963, O17964, O17965, O17966, O17967, O17968, O17969, O17970, O17971, O17972, O17973, O17974, O17975, O17976, O17977, O17978, O17979, O17980, O17981, O17982, O17983, O17984, O17985, O17986, O17987, O17988, O17989, O17990, O17991, O17992, O17993, O17994, O17995, O17996, O17997, O17998, O17999, O18000, O18001, O18002, O18003, O18004, O18005, O18006, O18007, O18008, O18009, O18010, O18011, O18012, O18013, O18014, O18015, O18016, O18017, O18018, O18019, O18020, O18021, O18022, O18023, O18024, O18025, O18026, O18027, O18028, O18029, O18030, O18031, O18032, O18033, O18034, O18035, O18036, O18037, O18038, O18039, O18040, O18041, O18042, O18043, O18044, O18045, O18046, O18047, O18048, O18049, O18050, O18051, O18052, O18053, O18054, O18055, O18056, O18057, O18058, O18059, O18060, O18061, O18062, O18063, O18064, O18065, O18066, O18067, O18068, O18069, O18070, O18071, O18072, O18073, O18074, O18075, O18076, O18077, O18078, O18079, O18080, O18081, O18082, O18083, O18084, O18085, O18086, O18087, O18088, O18089, O18090, O18091, O18092, O18093, O18094, O18095, O18096, O18097, O18098, O18099, O18100, O18101, O18102, O18103, O18104, O18105, O18106, O18107, O18108, O18109, O18110, O18111, O18112, O18113, O18114, O18115, O18116, O18117, O18118, O18119, O18120, O18121, O18122, O18123, O18124, O18125, O18126, O18127, O18128, O18129, O18130, O18131, O18132, O18133, O18134, O18135, O18136, O18137, O18138, O18139, O18140, O18141, O18142, O18143, O18144, O18145, O18146, O18147, O18148, O18149, O18150, O18151, O18152, O18153, O18154, O18155, O18156, O18157, O18158, O18159, O18160, O18161, O18162, O18163, O18164, O18165, O18166, O18167, O18168, O18169, O18170, O18171, O18172, O18173, O18174, O18175, O18176, O18177, O18178, O18179, O18180, O18181, O18182, O18183, O18184, O18185, O18186, O18187, O18188, O18189, O18190, O18191, O18192, O18193, O18194, O18195, O18196, O18197, O18198, O18199, O18200, O18201, O18202, O18203, O18204, O18205, O18206, O18207, O18208, O18209, O18210, O18211, O18212, O18213, O18214, O18215, O18216, O18217, O18218, O18219, O18220, O18221, O18222, O18223, O18224, O18225, O18226, O18227, O18228, O18229, O18230, O18231, O18232, O18233, O18234, O18235, O18236, O18237, O18238, O18239, O18240, O18241, O18242, O18243, O18244, O18245, O18246, O18247, O18248, O18249, O18250, O18251, O18252, O18253, O18254, O18255, O18256, O18257, O18258, O18259, O18260, O18261, O18262, O18263, O18264, O18265, O18266, O18267, O18268, O18269, O18270, O18271, O18272, O18273, O18274, O18275, O18276, O18277, O18278, O18279, O18280, O18281, O18282, O18283, O18284, O18285, O18286, O18287, O18288, O18289, O18290, O18291, O18292, O18293, O18294, O18295, O18296, O18297, O18298, O18299, O18300, O18301, O18302, O18303, O18304, O18305, O18306, O18307, O18308, O18309, O18310, O18311, O18312, O18313, O18314, O18315, O18316, O18317, O18318, O18319, O18320, O18321, O18322, O18323, O18324, O18325, O18326, O18327, O18328, O18329, O18330, O18331, O18332, O18333, O18334, O18335, O18336, O18337, O18338, O18339, O18340, O18341, O18342, O18343, O18344, O18345, O18346, O18347, O18348, O18349, O18350, O18351, O18352, O18353, O18354, O18355, O18356, O18357, O18358, O18359, O18360, O18361, O18362, O18363, O18364, O18365, O18366, O18367, O18368, O18369, O18370, O18371, O18372, O18373, O18374, O18375, O18376, O18377, O18378, O18379, O18380, O18381, O18382, O18383, O18384, O18385, O18386, O18387, O18388, O18389, O18390, O18391, O18392, O18393, O18394, O18395, O18396, O18397, O18398, O18399, O18400, O18401, O18402, O18403, O18404, O18405, O18406, O18407, O18408, O18409, O18410, O18411, O18412, O18413, O18414, O18415, O18416, O18417, O18418, O18419, O18420, O18421, O18422, O18423, O18424, O18425, O18426, O18427, O18428, O18429, O18430, O18431, O18432, O18433, O18434, O18435, O18436, O18437, O18438, O18439, O18440, O18441, O18442, O18443, O18444, O18445, O18446, O18447, O18448, O18449, O18450, O18451, O18452, O18453, O18454, O18455, O18456, O18457, O18458, O18459, O18460, O18461, O18462, O18463, O18464, O18465, O18466, O18467, O18468, O18469, O18470, O18471, O18472, O18473, O18474, O18475, O18476, O18477, O18478, O18479, O18480, O18481, O18482, O18483, O18484, O18485, O18486, O18487, O18488, O18489, O18490, O18491, O18492, O18493, O18494, O18495, O18496, O18497, O18498, O18499, O18500, O18501, O18502, O18503, O18504, O18505, O18506, O18507, O18508, O18509, O18510, O18511, O18512, O18513, O18514, O18515, O18516, O18517, O18518, O18519, O18520, O18521, O18522, O18523, O18524, O18525, O18526, O18527, O18528, O18529, O18530, O18531, O18532, O18533, O18534, O18535, O18536, O18537, O18538, O18539, O18540, O18541, O18542, O18543, O18544, O18545, O18546, O18547, O18548, O18549, O18550, O18551, O18552, O18553, O18554, O18555, O18556, O18557, O18558, O18559, O18560, O18561, O18562, O18563, O18564, O18565, O18566, O18567, O18568, O18569, O18570, O18571, O18572, O18573, O18574, O18575, O18576, O18577, O18578, O18579, O18580, O18581, O18582, O18583, O18584, O18585, O18586, O18587, O18588, O18589, O18590, O18591, O18592, O18593, O18594, O18595, O18596, O18597, O18598, O18599, O18600, O18601, O18602, O18603, O18604, O18605, O18606, O18607, O18608, O18609, O18610, O18611, O18612, O18613, O18614, O18615, O18616, O18617, O18618, O18619, O18620, O18621, O18622, O18623, O18624, O18625, O18626, O18627, O18628, O18629, O18630, O18631, O18632, O18633, O18634, O18635, O18636, O18637, O18638, O18639, O18640, O18641, O18642, O18643, O18644, O18645, O18646, O18647, O18648, O18649, O18650, O18651, O18652, O18653, O18654, O18655, O18656, O18657, O18658, O18659, O18660, O18661, O18662, O18663, O18664, O18665, O18666, O18667, O18668, O18669, O18670, O18671, O18672, O18673, O18674, O18675, O18676, O18677, O18678, O18679, O18680, O18681, O18682, O18683, O18684, O18685, O18686, O18687, O18688, O18689, O18690, O18691, O18692, O18693, O18694, O18695, O18696, O18697, O18698, O18699, O18700, O18701, O18702, O18703, O18704, O18705, O18706, O18707, O18708, O18709, O18710, O18711, O18712, O18713, O18714, O18715, O18716, O18717, O18718, O18719, O18720, O18721, O18722, O18723, O18724, O18725, O18726, O18727, O18728, O18729, O18730, O18731, O18732, O18733, O18734, O18735, O18736, O18737, O18738, O18739, O18740, O18741, O18742, O18743, O18744, O18745, O18746, O18747, O18748, O18749, O18750, O18751, O18752, O18753, O18754, O18755, O18756, O18757, O18758, O18759, O18760, O18761, O18762, O18763, O18764, O18765, O18766, O18767, O18768, O18769, O18770, O18771, O18772, O18773, O18774, O18775, O18776, O18777, O18778, O18779, O18780, O18781, O18782, O18783, O18784, O18785, O18786, O18787, O18788, O18789, O18790, O18791, O18792, O18793, O18794, O18795, O18796, O18797, O18798, O18799, O18800, O18801, O18802, O18803, O18804, O18805, O18806, O18807, O18808, O18809, O18810, O18811, O18812, O18813, O18814, O18815, O18816, O18817, O18818, O18819, O18820, O18821, O18822, O18823, O18824, O18825, O18826, O18827, O18828, O18829, O18830, O18831, O18832, O18833, O18834, O18835, O18836, O18837, O18838, O18839, O18840, O18841, O18842, O18843, O18844, O18845, O18846, O18847, O18848, O18849, O18850, O18851, O18852, O18853, O18854, O18855, O18856, O18857, O18858, O18859, O18860, O18861, O18862, O18863, O18864, O18865, O18866, O18867, O18868, O18869, O18870, O18871, O18872, O18873, O18874, O18875, O18876, O18877, O18878, O18879, O18880, O18881, O18882, O18883, O18884, O18885, O18886, O18887, O18888, O18889, O18890, O18891, O18892, O18893, O18894, O18895, O18896, O18897, O18898, O18899, O18900, O18901, O18902, O18903, O18904, O18905, O18906, O18907, O18908, O18909, O18910, O18911, O18912, O18913, O18914, O18915, O18916, O18917, O18918, O18919, O18920, O18921, O18922, O18923, O18924, O18925, O18926, O18927, O18928, O18929, O18930, O18931, O18932, O18933, O18934, O18935, O18936, O18937, O18938, O18939, O18940, O18941, O18942, O18943, O18944, O18945, O18946, O18947, O18948, O18949, O18950, O18951, O18952, O18953, O18954, O18955, O18956, O18957, O18958, O18959, O18960, O18961, O18962, O18963, O18964, O18965, O18966, O18967, O18968, O18969, O18970, O18971, O18972, O18973, O18974, O18975, O18976, O18977, O18978, O18979, O18980, O18981, O18982, O18983, O18984, O18985, O18986, O18987, O18988, O18989, O18990, O18991, O18992, O18993, O18994, O18995, O18996, O18997, O18998, O18999, O19000, O19001, O19002, O19003, O19004, O19005, O19006, O19007, O19008, O19009, O19010, O19011, O19012, O19013, O19014, O19015, O19016, O19017, O19018, O19019, O19020, O19021, O19022, O19023, O19024, O19025, O19026, O19027, O19028, O19029, O19030, O19031, O19032, O19033, O19034, O19035, O19036, O19037, O19038, O19039, O19040, O19041, O19042, O19043, O19044, O19045, O19046, O19047, O19048, O19049, O19050, O19051, O19052, O19053, O19054, O19055, O19056, O19057, O19058, O19059, O19060, O19061, O19062, O19063, O19064, O19065, O19066, O19067, O19068, O19069, O19070, O19071, O19072, O19073, O19074, O19075, O19076, O19077, O19078, O19079, O19080, O19081, O19082, O19083, O19084, O19085, O19086, O19087, O19088, O19089, O19090, O19091, O19092, O19093, O19094, O19095, O19096, O19097, O19098, O19099, O19100, O19101, O19102, O19103, O19104, O19105, O19106, O19107, O19108, O19109, O19110, O19111, O19112, O19113, O19114, O19115, O19116, O19117, O19118, O19119, O19120, O19121, O19122, O19123, O19124, O19125, O19126, O19127, O19128, O19129, O19130, O19131, O19132, O19133, O19134, O19135, O19136, O19137, O19138, O19139, O19140, O19141, O19142, O19143, O19144, O19145, O19146, O19147, O19148, O19149, O19150, O19151, O19152, O19153, O19154, O19155, O19156, O19157, O19158, O19159, O19160, O19161, O19162, O19163, O19164, O19165, O19166, O19167, O19168, O19169, O19170, O19171, O19172, O19173, O19174, O19175, O19176, O19177, O19178, O19179, O19180, O19181, O19182, O19183, O19184, O19185, O19186, O19187, O19188, O19189, O19190, O19191, O19192, O19193, O19194, O19195, O19196, O19197, O19198, O19199, O19200, O19201, O19202, O19203, O19204, O19205, O19206, O19207, O19208, O19209, O19210, O19211, O19212, O19213, O19214, O19215, O19216, O19217, O19218, O19219, O19220, O19221, O19222, O19223, O19224, O19225, O19226, O19227, O19228, O19229, O19230, O19231, O19232, O19233, O19234, O19235, O19236, O19237, O19238, O19239, O19240, O19241, O19242, O19243, O19244, O19245, O19246, O19247, O19248, O19249, O19250, O19251, O19252, O19253, O19254, O19255, O19256, O19257, O19258, O19259, O19260, O19261, O19262, O19263, O19264, O19265, O19266, O19267, O19268, O19269, O19270, O19271, O19272, O19273, O19274, O19275, O19276, O19277, O19278, O19279, O19280, O19281, O19282, O19283, O19284, O19285, O19286, O19287, O19288, O19289, O19290, O19291, O19292, O19293, O19294, O19295, O19296, O19297, O19298, O19299, O19300, O19301, O19302, O19303, O19304, O19305, O19306, O19307, O19308, O19309, O19310, O19311, O19312, O19313, O19314, O19315, O19316, O19317, O19318, O19319, O19320, O19321, O19322, O19323, O19324, O19325, O19326, O19327, O19328, O19329, O19330, O19331, O19332, O19333, O19334, O19335, O19336, O19337, O19338, O19339, O19340, O19341, O19342, O19343, O19344, O19345, O19346, O19347, O19348, O19349, O19350, O19351, O19352, O19353, O19354, O19355, O19356, O19357, O19358, O19359, O19360, O19361, O19362, O19363, O19364, O19365, O19366, O19367, O19368, O19369, O19370, O19371, O19372, O19373, O19374, O19375, O19376, O19377, O19378, O19379, O19380, O19381, O19382, O19383, O19384, O19385, O19386, O19387, O19388, O19389, O19390, O19391, O19392, O19393, O19394, O19395, O19396, O19397, O19398, O19399, O19400, O19401, O19402, O19403, O19404, O19405, O19406, O19407, O19408, O19409, O19410, O19411, O19412, O19413, O19414, O19415, O19416, O19417, O19418, O19419, O19420, O19421, O19422, O19423, O19424, O19425, O19426, O19427, O19428, O19429, O19430, O19431, O19432, O19433, O19434, O19435, O19436, O19437, O19438, O19439, O19440, O19441, O19442, O19443, O19444, O19445, O19446, O19447, O19448, O19449, O19450, O19451, O19452, O19453, O19454, O19455, O19456, O19457, O19458, O19459, O19460, O19461, O19462, O19463, O19464, O19465, O19466, O19467, O19468, O19469, O19470, O19471, O19472, O19473, O19474, O19475, O19476, O19477, O19478, O19479, O19480, O19481, O19482, O19483, O19484, O19485, O19486, O19487, O19488, O19489, O19490, O19491, O19492, O19493, O19494, O19495, O19496, O19497, O19498, O19499, O19500, O19501, O19502, O19503, O19504, O19505, O19506, O19507, O19508, O19509, O19510, O19511, O19512, O19513, O19514, O19515, O19516, O19517, O19518, O19519, O19520, O19521, O19522, O19523, O19524, O19525, O19526, O19527, O19528, O19529, O19530, O19531, O19532, O19533, O19534, O19535, O19536, O19537, O19538, O19539, O19540, O19541, O19542, O19543, O19544, O19545, O19546, O19547, O19548, O19549, O19550, O19551, O19552, O19553, O19554, O19555, O19556, O19557, O19558, O19559, O19560, O19561, O19562, O19563, O19564, O19565, O19566, O19567, O19568, O19569, O19570, O19571, O19572, O19573, O19574, O19575, O19576, O19577, O19578, O19579, O19580, O19581, O19582, O19583, O19584, O19585, O19586, O19587, O19588, O19589, O19590, O19591, O19592, O19593, O19594, O19595, O19596, O19597, O19598, O19599, O19600, O19601, O19602, O19603, O19604, O19605, O19606, O19607, O19608, O19609, O19610, O19611, O19612, O19613, O19614, O19615, O19616, O19617, O19618, O19619, O19620, O19621, O19622, O19623, O19624, O19625, O19626, O19627, O19628, O19629, O19630, O19631, O19632, O19633, O19634, O19635, O19636, O19637, O19638, O19639, O19640, O19641, O19642, O19643, O19644, O19645, O19646, O19647, O19648, O19649, O19650, O19651, O19652, O19653, O19654, O19655, O19656, O19657, O19658, O19659, O19660, O19661, O19662, O19663, O19664, O19665, O19666, O19667, O19668, O19669, O19670, O19671, O19672, O19673, O19674, O19675, O19676, O19677, O19678, O19679, O19680, O19681, O19682, O19683, O19684, O19685, O19686, O19687, O19688, O19689, O19690, O19691, O19692, O19693, O19694, O19695, O19696, O19697, O19698, O19699, O19700, O19701, O19702, O19703, O19704, O19705, O19706, O19707, O19708, O19709, O19710, O19711, O19712, O19713, O19714, O19715, O19716, O19717, O19718, O19719, O19720, O19721, O19722, O19723, O19724, O19725, O19726, O19727, O19728, O19729, O19730, O19731, O19732, O19733, O19734, O19735, O19736, O19737, O19738, O19739, O19740, O19741, O19742, O19743, O19744, O19745, O19746, O19747, O19748, O19749, O19750, O19751, O19752, O19753, O19754, O19755, O19756, O19757, O19758, O19759, O19760, O19761, O19762);
  input I0, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I16, I17, I18, I19, I20, I21, I22, I23, I24, I26, I27, I28, I29, I30, I31, I32, I34, I36, I38, I39, I40, I42, I43, I44, I45, I46, I48, I49, I50, I51, I52, I54, I55, I56, I57, I58, I60, I61, I62, I64, I65, I66, I68, I70, I71, I72, I74, I75, I76, I78, I79, I80, I81, I82, I84, I85, I86, I88, I90, I91, I92, I94, I95, I96, I98, I100, I102, I103, I104, I106, I108, I109, I110, I111, I112, I113, I114, I115, I116, I117, I118, I120, I121, I122, I123, I124, I126, I128, I130, I132, I134, I135, I136, I137, I138, I140, I142, I144, I145, I146, I147, I148, I150, I151, I152, I153, I154, I156, I157, I158, I160, I161, I162, I163, I164, I165, I166, I168, I169, I170, I171, I172, I174, I175, I176, I178, I179, I180, I181, I182, I184, I185, I186, I188, I190, I191, I192, I193, I194, I195, I196, I197, I198, I200, I202, I203, I204, I206, I207, I208, I209, I210, I212, I213, I214, I215, I216, I217, I218, I219, I220, I221, I222, I223, I224, I225, I226, I227, I228, I229, I230, I231, I232, I233, I234, I235, I236, I237, I238, I239, I240, I241, I242, I243, I244, I245, I246, I247, I248, I249, I250, I252, I253, I254, I255, I256, I257, I258, I259, I260, I261, I262, I263, I264, I266, I267, I268, I269, I270, I271, I272, I274, I276, I277, I278, I280, I282, I283, I284, I285, I286, I288, I289, I290, I291, I292, I294, I296, I297, I298, I299, I300, I301, I302, I303, I304, I305, I306, I308, I309, I310, I312, I313, I314, I315, I316, I317, I318, I319, I320, I322, I323, I324, I326, I328, I329, I330, I331, I332, I334, I335, I336, I337, I338, I339, I340, I342, I344, I346, I347, I348, I349, I350, I351, I352, I353, I354, I355, I356, I357, I358, I360, I361, I362, I364, I365, I366, I368, I370, I371, I372, I374, I375, I376, I378, I380, I382, I384, I385, I386, I387, I388, I389, I390, I391, I392, I393, I394, I396, I398, I400, I401, I402, I404, I405, I406, I407, I408, I409, I410, I412, I413, I414, I415, I416, I417, I418, I420, I421, I422, I423, I424, I426, I428, I429, I430, I431, I432, I433, I434, I435, I436, I437, I438, I439, I440, I441, I442, I443, I444, I445, I446, I447, I448, I450, I451, I452, I454, I455, I456, I457, I458, I459, I460, I462, I463, I464, I466, I467, I468, I469, I470, I471, I472, I474, I475, I476, I477, I478, I479, I480, I481, I482, I483, I484, I485, I486, I488, I489, I490, I491, I492, I493, I494, I495, I496, I498, I499, I500, I501, I502, I503, I504, I505, I506, I507, I508, I509, I510, I511, I512, I514, I516, I517, I518, I519, I520, I521, I522, I524, I525, I526, I527, I528, I530, I531, I532, I533, I534, I535, I536, I537, I538, I539, I540, I541, I542, I543, I544, I546, I547, I548, I549, I550, I551, I552, I554, I555, I556, I557, I558, I559, I560, I562, I563, I564, I565, I566, I567, I568, I570, I572, I574, I575, I576, I578, I579, I580, I581, I582, I583, I584, I586, I587, I588, I590, I592, I594, I595, I596, I597, I598, I600, I601, I602, I603, I604, I605, I606, I607, I608, I609, I610, I612, I613, I614, I615, I616, I618, I619, I620, I621, I622, I623, I624, I625, I626, I628, I629, I630, I631, I632, I633, I634, I635, I636, I637, I638, I639, I640, I641, I642, I643, I644, I646, I647, I648, I649, I650, I652, I654, I655, I656, I657, I658, I659, I660, I661, I662, I664, I665, I666, I668, I669, I670, I671, I672, I673, I674, I675, I676, I677, I678, I679, I680, I681, I682, I683, I684, I685, I686, I687, I688, I690, I691, I692, I693, I694, I695, I696, I697, I698, I700, I701, I702, I704, I705, I706, I707, I708, I710, I711, I712, I713, I714, I715, I716, I718, I719, I720, I721, I722, I723, I724, I725, I726, I727, I728, I729, I730, I731, I732, I734, I735, I736, I737, I738, I740, I741, I742, I743, I744, I745, I746, I747, I748, I750, I752, I753, I754, I755, I756, I758, I759, I760, I762, I764, I765, I766, I767, I768, I770, I771, I772, I773, I774, I776, I777, I778, I779, I780, I781, I782, I784, I785, I786, I787, I788, I790, I791, I792, I793, I794, I796, I797, I798, I799, I800, I802, I804, I806, I808, I809, I810, I811, I812, I813, I814, I815, I816, I817, I818, I819, I820, I821, I822, I824, I825, I826, I827, I828, I829, I830, I831, I832, I833, I834, I836, I838, I839, I840, I842, I843, I844, I846, I848, I849, I850, I852, I853, I854, I856, I857, I858, I859, I860, I861, I862, I863, I864, I866, I868, I870, I871, I872, I873, I874, I875, I876, I877, I878, I879, I880, I881, I882, I884, I885, I886, I887, I888, I889, I890, I892, I893, I894, I895, I896, I898, I900, I901, I902, I903, I904, I905, I906, I907, I908, I909, I910, I911, I912, I913, I914, I915, I916, I917, I918, I919, I920, I921, I922, I923, I924, I925, I926, I927, I928, I929, I930, I932, I933, I934, I936, I937, I938, I939, I940, I941, I942, I943, I944, I945, I946, I947, I948, I950, I952, I953, I954, I956, I957, I958, I960, I962, I963, I964, I965, I966, I967, I968, I969, I970, I972, I973, I974, I975, I976, I977, I978, I980, I981, I982, I983, I984, I986, I987, I988, I989, I990, I991, I992, I993, I994, I995, I996, I998, I999, I1000, I1001, I1002, I1003, I1004, I1005, I1006, I1008, I1010, I1011, I1012, I1013, I1014, I1015, I1016, I1018, I1019, I1020, I1021, I1022, I1024, I1025, I1026, I1027, I1028, I1029, I1030, I1031, I1032, I1033, I1034, I1036, I1038, I1040, I1041, I1042, I1043, I1044, I1045, I1046, I1047, I1048, I1049, I1050, I1051, I1052, I1053, I1054, I1055, I1056, I1058, I1059, I1060, I1062, I1064, I1065, I1066, I1067, I1068, I1069, I1070, I1072, I1073, I1074, I1075, I1076, I1078, I1079, I1080, I1082, I1084, I1086, I1087, I1088, I1089, I1090, I1091, I1092, I1094, I1095, I1096, I1098, I1100, I1102, I1103, I1104, I1105, I1106, I1107, I1108, I1110, I1111, I1112, I1113, I1114, I1115, I1116, I1117, I1118, I1119, I1120, I1121, I1122, I1123, I1124, I1126, I1127, I1128, I1129, I1130, I1131, I1132, I1133, I1134, I1135, I1136, I1138, I1139, I1140, I1141, I1142, I1143, I1144, I1145, I1146, I1147, I1148, I1149, I1150, I1151, I1152, I1153, I1154, I1156, I1157, I1158, I1159, I1160, I1161, I1162, I1163, I1164, I1165, I1166, I1167, I1168, I1170, I1171, I1172, I1173, I1174, I1175, I1176, I1177, I1178, I1179, I1180, I1181, I1182, I1184, I1186, I1187, I1188, I1189, I1190, I1192, I1193, I1194, I1195, I1196, I1197, I1198, I1199, I1200, I1201, I1202, I1204, I1206, I1208, I1209, I1210, I1211, I1212, I1213, I1214, I1215, I1216, I1217, I1218, I1219, I1220, I1221, I1222, I1224, I1225, I1226, I1228, I1229, I1230, I1231, I1232, I1233, I1234, I1235, I1236, I1238, I1239, I1240, I1242, I1243, I1244, I1245, I1246, I1247, I1248, I1250, I1251, I1252, I1253, I1254, I1255, I1256, I1258, I1259, I1260, I1261, I1262, I1263, I1264, I1265, I1266, I1267, I1268, I1270, I1271, I1272, I1273, I1274, I1276, I1277, I1278, I1280, I1281, I1282, I1283, I1284, I1286, I1287, I1288, I1289, I1290, I1292, I1293, I1294, I1296, I1298, I1299, I1300, I1301, I1302, I1303, I1304, I1305, I1306, I1307, I1308, I1310, I1312, I1314, I1316, I1317, I1318, I1319, I1320, I1321, I1322, I1323, I1324, I1325, I1326, I1328, I1329, I1330, I1331, I1332, I1333, I1334, I1336, I1337, I1338, I1339, I1340, I1341, I1342, I1343, I1344, I1345, I1346, I1347, I1348, I1350, I1352, I1353, I1354, I1355, I1356, I1357, I1358, I1360, I1361, I1362, I1364, I1365, I1366, I1367, I1368, I1370, I1372, I1373, I1374, I1375, I1376, I1377, I1378, I1380, I1381, I1382, I1384, I1385, I1386, I1388, I1389, I1390, I1391, I1392, I1393, I1394, I1395, I1396, I1398, I1399, I1400, I1401, I1402, I1403, I1404, I1406, I1407, I1408, I1409, I1410, I1411, I1412, I1414, I1415, I1416, I1418, I1419, I1420, I1421, I1422, I1423, I1424, I1425, I1426, I1427, I1428, I1429, I1430, I1431, I1432, I1434, I1435, I1436, I1437, I1438, I1439, I1440, I1441, I1442, I1444, I1445, I1446, I1447, I1448, I1449, I1450, I1452, I1453, I1454, I1455, I1456, I1457, I1458, I1459, I1460, I1461, I1462, I1463, I1464, I1465, I1466, I1467, I1468, I1470, I1471, I1472, I1473, I1474, I1475, I1476, I1477, I1478, I1480, I1482, I1483, I1484, I1486, I1488, I1489, I1490, I1491, I1492, I1493, I1494, I1495, I1496, I1497, I1498, I1500, I1501, I1502, I1503, I1504, I1505, I1506, I1507, I1508, I1509, I1510, I1512, I1513, I1514, I1516, I1518, I1519, I1520, I1522, I1523, I1524, I1526, I1528, I1529, I1530, I1531, I1532, I1533, I1534, I1535, I1536, I1538, I1540, I1541, I1542, I1544, I1545, I1546, I1547, I1548, I1550, I1552, I1553, I1554, I1556, I1557, I1558, I1560, I1561, I1562, I1563, I1564, I1565, I1566, I1568, I1569, I1570, I1571, I1572, I1573, I1574, I1575, I1576, I1577, I1578, I1579, I1580, I1582, I1584, I1585, I1586, I1588, I1589, I1590, I1591, I1592, I1593, I1594, I1596, I1597, I1598, I1599, I1600, I1602, I1603, I1604, I1606, I1608, I1609, I1610, I1611, I1612, I1614, I1616, I1617, I1618, I1619, I1620, I1621, I1622, I1624, I1626, I1628, I1629, I1630, I1632, I1633, I1634, I1636, I1637, I1638, I1639, I1640, I1642, I1644, I1646, I1647, I1648, I1649, I1650, I1651, I1652, I1653, I1654, I1656, I1657, I1658, I1659, I1660, I1662, I1663, I1664, I1665, I1666, I1667, I1668, I1669, I1670, I1671, I1672, I1674, I1675, I1676, I1677, I1678, I1679, I1680, I1681, I1682, I1684, I1685, I1686, I1687, I1688, I1689, I1690, I1692, I1694, I1695, I1696, I1697, I1698, I1700, I1701, I1702, I1703, I1704, I1706, I1707, I1708, I1709, I1710, I1711, I1712, I1714, I1715, I1716, I1717, I1718, I1719, I1720, I1722, I1724, I1725, I1726, I1727, I1728, I1729, I1730, I1731, I1732, I1733, I1734, I1736, I1737, I1738, I1739, I1740, I1742, I1743, I1744, I1746, I1747, I1748, I1749, I1750, I1751, I1752, I1753, I1754, I1755, I1756, I1758, I1759, I1760, I1761, I1762, I1763, I1764, I1766, I1768, I1769, I1770, I1772, I1773, I1774, I1775, I1776, I1777, I1778, I1779, I1780, I1782, I1783, I1784, I1786, I1788, I1790, I1792, I1793, I1794, I1795, I1796, I1798, I1799, I1800, I1801, I1802, I1803, I1804, I1806, I1807, I1808, I1809, I1810, I1811, I1812, I1813, I1814, I1815, I1816, I1818, I1819, I1820, I1822, I1824, I1825, I1826, I1828, I1830, I1831, I1832, I1834, I1835, I1836, I1837, I1838, I1839, I1840, I1841, I1842, I1843, I1844, I1846, I1847, I1848, I1850, I1851, I1852, I1853, I1854, I1856, I1858, I1859, I1860, I1861, I1862, I1863, I1864, I1865, I1866, I1868, I1870, I1872, I1873, I1874, I1875, I1876, I1877, I1878, I1880, I1881, I1882, I1883, I1884, I1886, I1887, I1888, I1889, I1890, I1892, I1893, I1894, I1895, I1896, I1898, I1900, I1901, I1902, I1903, I1904, I1906, I1907, I1908, I1909, I1910, I1911, I1912, I1913, I1914, I1915, I1916, I1917, I1918, I1919, I1920, I1921, I1922, I1923, I1924, I1925, I1926, I1927, I1928, I1930, I1931, I1932, I1933, I1934, I1935, I1936, I1937, I1938, I1939, I1940, I1941, I1942, I1943, I1944, I1945, I1946, I1948, I1949, I1950, I1952, I1953, I1954, I1955, I1956, I1957, I1958, I1959, I1960, I1962, I1963, I1964, I1965, I1966, I1968, I1969, I1970, I1972, I1974, I1975, I1976, I1977, I1978, I1979, I1980, I1981, I1982, I1983, I1984, I1985, I1986, I1987, I1988, I1990, I1991, I1992, I1993, I1994, I1996, I1997, I1998;
  output O0, O1, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15, O16, O17, O18, O19, O20, O21, O22, O23, O24, O25, O26, O27, O28, O29, O30, O31, O32, O33, O34, O35, O36, O37, O38, O39, O40, O41, O42, O43, O44, O45, O46, O47, O48, O49, O50, O51, O52, O53, O54, O55, O56, O57, O58, O59, O60, O61, O62, O63, O64, O65, O66, O67, O68, O69, O70, O71, O72, O73, O74, O75, O76, O77, O78, O79, O80, O81, O82, O83, O84, O85, O86, O87, O88, O89, O90, O91, O92, O93, O94, O95, O96, O97, O98, O99, O100, O101, O102, O103, O104, O105, O106, O107, O108, O109, O110, O111, O112, O113, O114, O115, O116, O117, O118, O119, O120, O121, O122, O123, O124, O125, O126, O127, O128, O129, O130, O131, O132, O133, O134, O135, O136, O137, O138, O139, O140, O141, O142, O143, O144, O145, O146, O147, O148, O149, O150, O151, O152, O153, O154, O155, O156, O157, O158, O159, O160, O161, O162, O163, O164, O165, O166, O167, O168, O169, O170, O171, O172, O173, O174, O175, O176, O177, O178, O179, O180, O181, O182, O183, O184, O185, O186, O187, O188, O189, O190, O191, O192, O193, O194, O195, O196, O197, O198, O199, O200, O201, O202, O203, O204, O205, O206, O207, O208, O209, O210, O211, O212, O213, O214, O215, O216, O217, O218, O219, O220, O221, O222, O223, O224, O225, O226, O227, O228, O229, O230, O231, O232, O233, O234, O235, O236, O237, O238, O239, O240, O241, O242, O243, O244, O245, O246, O247, O248, O249, O250, O251, O252, O253, O254, O255, O256, O257, O258, O259, O260, O261, O262, O263, O264, O265, O266, O267, O268, O269, O270, O271, O272, O273, O274, O275, O276, O277, O278, O279, O280, O281, O282, O283, O284, O285, O286, O287, O288, O289, O290, O291, O292, O293, O294, O295, O296, O297, O298, O299, O300, O301, O302, O303, O304, O305, O306, O307, O308, O309, O310, O311, O312, O313, O314, O315, O316, O317, O318, O319, O320, O321, O322, O323, O324, O325, O326, O327, O328, O329, O330, O331, O332, O333, O334, O335, O336, O337, O338, O339, O340, O341, O342, O343, O344, O345, O346, O347, O348, O349, O350, O351, O352, O353, O354, O355, O356, O357, O358, O359, O360, O361, O362, O363, O364, O365, O366, O367, O368, O369, O370, O371, O372, O373, O374, O375, O376, O377, O378, O379, O380, O381, O382, O383, O384, O385, O386, O387, O388, O389, O390, O391, O392, O393, O394, O395, O396, O397, O398, O399, O400, O401, O402, O403, O404, O405, O406, O407, O408, O409, O410, O411, O412, O413, O414, O415, O416, O417, O418, O419, O420, O421, O422, O423, O424, O425, O426, O427, O428, O429, O430, O431, O432, O433, O434, O435, O436, O437, O438, O439, O440, O441, O442, O443, O444, O445, O446, O447, O448, O449, O450, O451, O452, O453, O454, O455, O456, O457, O458, O459, O460, O461, O462, O463, O464, O465, O466, O467, O468, O469, O470, O471, O472, O473, O474, O475, O476, O477, O478, O479, O480, O481, O482, O483, O484, O485, O486, O487, O488, O489, O490, O491, O492, O493, O494, O495, O496, O497, O498, O499, O500, O501, O502, O503, O504, O505, O506, O507, O508, O509, O510, O511, O512, O513, O514, O515, O516, O517, O518, O519, O520, O521, O522, O523, O524, O525, O526, O527, O528, O529, O530, O531, O532, O533, O534, O535, O536, O537, O538, O539, O540, O541, O542, O543, O544, O545, O546, O547, O548, O549, O550, O551, O552, O553, O554, O555, O556, O557, O558, O559, O560, O561, O562, O563, O564, O565, O566, O567, O568, O569, O570, O571, O572, O573, O574, O575, O576, O577, O578, O579, O580, O581, O582, O583, O584, O585, O586, O587, O588, O589, O590, O591, O592, O593, O594, O595, O596, O597, O598, O599, O600, O601, O602, O603, O604, O605, O606, O607, O608, O609, O610, O611, O612, O613, O614, O615, O616, O617, O618, O619, O620, O621, O622, O623, O624, O625, O626, O627, O628, O629, O630, O631, O632, O633, O634, O635, O636, O637, O638, O639, O640, O641, O642, O643, O644, O645, O646, O647, O648, O649, O650, O651, O652, O653, O654, O655, O656, O657, O658, O659, O660, O661, O662, O663, O664, O665, O666, O667, O668, O669, O670, O671, O672, O673, O674, O675, O676, O677, O678, O679, O680, O681, O682, O683, O684, O685, O686, O687, O688, O689, O690, O691, O692, O693, O694, O695, O696, O697, O698, O699, O700, O701, O702, O703, O704, O705, O706, O707, O708, O709, O710, O711, O712, O713, O714, O715, O716, O717, O718, O719, O720, O721, O722, O723, O724, O725, O726, O727, O728, O729, O730, O731, O732, O733, O734, O735, O736, O737, O738, O739, O740, O741, O742, O743, O744, O745, O746, O747, O748, O749, O750, O751, O752, O753, O754, O755, O756, O757, O758, O759, O760, O761, O762, O763, O764, O765, O766, O767, O768, O769, O770, O771, O772, O773, O774, O775, O776, O777, O778, O779, O780, O781, O782, O783, O784, O785, O786, O787, O788, O789, O790, O791, O792, O793, O794, O795, O796, O797, O798, O799, O800, O801, O802, O803, O804, O805, O806, O807, O808, O809, O810, O811, O812, O813, O814, O815, O816, O817, O818, O819, O820, O821, O822, O823, O824, O825, O826, O827, O828, O829, O830, O831, O832, O833, O834, O835, O836, O837, O838, O839, O840, O841, O842, O843, O844, O845, O846, O847, O848, O849, O850, O851, O852, O853, O854, O855, O856, O857, O858, O859, O860, O861, O862, O863, O864, O865, O866, O867, O868, O869, O870, O871, O872, O873, O874, O875, O876, O877, O878, O879, O880, O881, O882, O883, O884, O885, O886, O887, O888, O889, O890, O891, O892, O893, O894, O895, O896, O897, O898, O899, O900, O901, O902, O903, O904, O905, O906, O907, O908, O909, O910, O911, O912, O913, O914, O915, O916, O917, O918, O919, O920, O921, O922, O923, O924, O925, O926, O927, O928, O929, O930, O931, O932, O933, O934, O935, O936, O937, O938, O939, O940, O941, O942, O943, O944, O945, O946, O947, O948, O949, O950, O951, O952, O953, O954, O955, O956, O957, O958, O959, O960, O961, O962, O963, O964, O965, O966, O967, O968, O969, O970, O971, O972, O973, O974, O975, O976, O977, O978, O979, O980, O981, O982, O983, O984, O985, O986, O987, O988, O989, O990, O991, O992, O993, O994, O995, O996, O997, O998, O999, O1000, O1001, O1002, O1003, O1004, O1005, O1006, O1007, O1008, O1009, O1010, O1011, O1012, O1013, O1014, O1015, O1016, O1017, O1018, O1019, O1020, O1021, O1022, O1023, O1024, O1025, O1026, O1027, O1028, O1029, O1030, O1031, O1032, O1033, O1034, O1035, O1036, O1037, O1038, O1039, O1040, O1041, O1042, O1043, O1044, O1045, O1046, O1047, O1048, O1049, O1050, O1051, O1052, O1053, O1054, O1055, O1056, O1057, O1058, O1059, O1060, O1061, O1062, O1063, O1064, O1065, O1066, O1067, O1068, O1069, O1070, O1071, O1072, O1073, O1074, O1075, O1076, O1077, O1078, O1079, O1080, O1081, O1082, O1083, O1084, O1085, O1086, O1087, O1088, O1089, O1090, O1091, O1092, O1093, O1094, O1095, O1096, O1097, O1098, O1099, O1100, O1101, O1102, O1103, O1104, O1105, O1106, O1107, O1108, O1109, O1110, O1111, O1112, O1113, O1114, O1115, O1116, O1117, O1118, O1119, O1120, O1121, O1122, O1123, O1124, O1125, O1126, O1127, O1128, O1129, O1130, O1131, O1132, O1133, O1134, O1135, O1136, O1137, O1138, O1139, O1140, O1141, O1142, O1143, O1144, O1145, O1146, O1147, O1148, O1149, O1150, O1151, O1152, O1153, O1154, O1155, O1156, O1157, O1158, O1159, O1160, O1161, O1162, O1163, O1164, O1165, O1166, O1167, O1168, O1169, O1170, O1171, O1172, O1173, O1174, O1175, O1176, O1177, O1178, O1179, O1180, O1181, O1182, O1183, O1184, O1185, O1186, O1187, O1188, O1189, O1190, O1191, O1192, O1193, O1194, O1195, O1196, O1197, O1198, O1199, O1200, O1201, O1202, O1203, O1204, O1205, O1206, O1207, O1208, O1209, O1210, O1211, O1212, O1213, O1214, O1215, O1216, O1217, O1218, O1219, O1220, O1221, O1222, O1223, O1224, O1225, O1226, O1227, O1228, O1229, O1230, O1231, O1232, O1233, O1234, O1235, O1236, O1237, O1238, O1239, O1240, O1241, O1242, O1243, O1244, O1245, O1246, O1247, O1248, O1249, O1250, O1251, O1252, O1253, O1254, O1255, O1256, O1257, O1258, O1259, O1260, O1261, O1262, O1263, O1264, O1265, O1266, O1267, O1268, O1269, O1270, O1271, O1272, O1273, O1274, O1275, O1276, O1277, O1278, O1279, O1280, O1281, O1282, O1283, O1284, O1285, O1286, O1287, O1288, O1289, O1290, O1291, O1292, O1293, O1294, O1295, O1296, O1297, O1298, O1299, O1300, O1301, O1302, O1303, O1304, O1305, O1306, O1307, O1308, O1309, O1310, O1311, O1312, O1313, O1314, O1315, O1316, O1317, O1318, O1319, O1320, O1321, O1322, O1323, O1324, O1325, O1326, O1327, O1328, O1329, O1330, O1331, O1332, O1333, O1334, O1335, O1336, O1337, O1338, O1339, O1340, O1341, O1342, O1343, O1344, O1345, O1346, O1347, O1348, O1349, O1350, O1351, O1352, O1353, O1354, O1355, O1356, O1357, O1358, O1359, O1360, O1361, O1362, O1363, O1364, O1365, O1366, O1367, O1368, O1369, O1370, O1371, O1372, O1373, O1374, O1375, O1376, O1377, O1378, O1379, O1380, O1381, O1382, O1383, O1384, O1385, O1386, O1387, O1388, O1389, O1390, O1391, O1392, O1393, O1394, O1395, O1396, O1397, O1398, O1399, O1400, O1401, O1402, O1403, O1404, O1405, O1406, O1407, O1408, O1409, O1410, O1411, O1412, O1413, O1414, O1415, O1416, O1417, O1418, O1419, O1420, O1421, O1422, O1423, O1424, O1425, O1426, O1427, O1428, O1429, O1430, O1431, O1432, O1433, O1434, O1435, O1436, O1437, O1438, O1439, O1440, O1441, O1442, O1443, O1444, O1445, O1446, O1447, O1448, O1449, O1450, O1451, O1452, O1453, O1454, O1455, O1456, O1457, O1458, O1459, O1460, O1461, O1462, O1463, O1464, O1465, O1466, O1467, O1468, O1469, O1470, O1471, O1472, O1473, O1474, O1475, O1476, O1477, O1478, O1479, O1480, O1481, O1482, O1483, O1484, O1485, O1486, O1487, O1488, O1489, O1490, O1491, O1492, O1493, O1494, O1495, O1496, O1497, O1498, O1499, O1500, O1501, O1502, O1503, O1504, O1505, O1506, O1507, O1508, O1509, O1510, O1511, O1512, O1513, O1514, O1515, O1516, O1517, O1518, O1519, O1520, O1521, O1522, O1523, O1524, O1525, O1526, O1527, O1528, O1529, O1530, O1531, O1532, O1533, O1534, O1535, O1536, O1537, O1538, O1539, O1540, O1541, O1542, O1543, O1544, O1545, O1546, O1547, O1548, O1549, O1550, O1551, O1552, O1553, O1554, O1555, O1556, O1557, O1558, O1559, O1560, O1561, O1562, O1563, O1564, O1565, O1566, O1567, O1568, O1569, O1570, O1571, O1572, O1573, O1574, O1575, O1576, O1577, O1578, O1579, O1580, O1581, O1582, O1583, O1584, O1585, O1586, O1587, O1588, O1589, O1590, O1591, O1592, O1593, O1594, O1595, O1596, O1597, O1598, O1599, O1600, O1601, O1602, O1603, O1604, O1605, O1606, O1607, O1608, O1609, O1610, O1611, O1612, O1613, O1614, O1615, O1616, O1617, O1618, O1619, O1620, O1621, O1622, O1623, O1624, O1625, O1626, O1627, O1628, O1629, O1630, O1631, O1632, O1633, O1634, O1635, O1636, O1637, O1638, O1639, O1640, O1641, O1642, O1643, O1644, O1645, O1646, O1647, O1648, O1649, O1650, O1651, O1652, O1653, O1654, O1655, O1656, O1657, O1658, O1659, O1660, O1661, O1662, O1663, O1664, O1665, O1666, O1667, O1668, O1669, O1670, O1671, O1672, O1673, O1674, O1675, O1676, O1677, O1678, O1679, O1680, O1681, O1682, O1683, O1684, O1685, O1686, O1687, O1688, O1689, O1690, O1691, O1692, O1693, O1694, O1695, O1696, O1697, O1698, O1699, O1700, O1701, O1702, O1703, O1704, O1705, O1706, O1707, O1708, O1709, O1710, O1711, O1712, O1713, O1714, O1715, O1716, O1717, O1718, O1719, O1720, O1721, O1722, O1723, O1724, O1725, O1726, O1727, O1728, O1729, O1730, O1731, O1732, O1733, O1734, O1735, O1736, O1737, O1738, O1739, O1740, O1741, O1742, O1743, O1744, O1745, O1746, O1747, O1748, O1749, O1750, O1751, O1752, O1753, O1754, O1755, O1756, O1757, O1758, O1759, O1760, O1761, O1762, O1763, O1764, O1765, O1766, O1767, O1768, O1769, O1770, O1771, O1772, O1773, O1774, O1775, O1776, O1777, O1778, O1779, O1780, O1781, O1782, O1783, O1784, O1785, O1786, O1787, O1788, O1789, O1790, O1791, O1792, O1793, O1794, O1795, O1796, O1797, O1798, O1799, O1800, O1801, O1802, O1803, O1804, O1805, O1806, O1807, O1808, O1809, O1810, O1811, O1812, O1813, O1814, O1815, O1816, O1817, O1818, O1819, O1820, O1821, O1822, O1823, O1824, O1825, O1826, O1827, O1828, O1829, O1830, O1831, O1832, O1833, O1834, O1835, O1836, O1837, O1838, O1839, O1840, O1841, O1842, O1843, O1844, O1845, O1846, O1847, O1848, O1849, O1850, O1851, O1852, O1853, O1854, O1855, O1856, O1857, O1858, O1859, O1860, O1861, O1862, O1863, O1864, O1865, O1866, O1867, O1868, O1869, O1870, O1871, O1872, O1873, O1874, O1875, O1876, O1877, O1878, O1879, O1880, O1881, O1882, O1883, O1884, O1885, O1886, O1887, O1888, O1889, O1890, O1891, O1892, O1893, O1894, O1895, O1896, O1897, O1898, O1899, O1900, O1901, O1902, O1903, O1904, O1905, O1906, O1907, O1908, O1909, O1910, O1911, O1912, O1913, O1914, O1915, O1916, O1917, O1918, O1919, O1920, O1921, O1922, O1923, O1924, O1925, O1926, O1927, O1928, O1929, O1930, O1931, O1932, O1933, O1934, O1935, O1936, O1937, O1938, O1939, O1940, O1941, O1942, O1943, O1944, O1945, O1946, O1947, O1948, O1949, O1950, O1951, O1952, O1953, O1954, O1955, O1956, O1957, O1958, O1959, O1960, O1961, O1962, O1963, O1964, O1965, O1966, O1967, O1968, O1969, O1970, O1971, O1972, O1973, O1974, O1975, O1976, O1977, O1978, O1979, O1980, O1981, O1982, O1983, O1984, O1985, O1986, O1987, O1988, O1989, O1990, O1991, O1992, O1993, O1994, O1995, O1996, O1997, O1998, O1999, O2000, O2001, O2002, O2003, O2004, O2005, O2006, O2007, O2008, O2009, O2010, O2011, O2012, O2013, O2014, O2015, O2016, O2017, O2018, O2019, O2020, O2021, O2022, O2023, O2024, O2025, O2026, O2027, O2028, O2029, O2030, O2031, O2032, O2033, O2034, O2035, O2036, O2037, O2038, O2039, O2040, O2041, O2042, O2043, O2044, O2045, O2046, O2047, O2048, O2049, O2050, O2051, O2052, O2053, O2054, O2055, O2056, O2057, O2058, O2059, O2060, O2061, O2062, O2063, O2064, O2065, O2066, O2067, O2068, O2069, O2070, O2071, O2072, O2073, O2074, O2075, O2076, O2077, O2078, O2079, O2080, O2081, O2082, O2083, O2084, O2085, O2086, O2087, O2088, O2089, O2090, O2091, O2092, O2093, O2094, O2095, O2096, O2097, O2098, O2099, O2100, O2101, O2102, O2103, O2104, O2105, O2106, O2107, O2108, O2109, O2110, O2111, O2112, O2113, O2114, O2115, O2116, O2117, O2118, O2119, O2120, O2121, O2122, O2123, O2124, O2125, O2126, O2127, O2128, O2129, O2130, O2131, O2132, O2133, O2134, O2135, O2136, O2137, O2138, O2139, O2140, O2141, O2142, O2143, O2144, O2145, O2146, O2147, O2148, O2149, O2150, O2151, O2152, O2153, O2154, O2155, O2156, O2157, O2158, O2159, O2160, O2161, O2162, O2163, O2164, O2165, O2166, O2167, O2168, O2169, O2170, O2171, O2172, O2173, O2174, O2175, O2176, O2177, O2178, O2179, O2180, O2181, O2182, O2183, O2184, O2185, O2186, O2187, O2188, O2189, O2190, O2191, O2192, O2193, O2194, O2195, O2196, O2197, O2198, O2199, O2200, O2201, O2202, O2203, O2204, O2205, O2206, O2207, O2208, O2209, O2210, O2211, O2212, O2213, O2214, O2215, O2216, O2217, O2218, O2219, O2220, O2221, O2222, O2223, O2224, O2225, O2226, O2227, O2228, O2229, O2230, O2231, O2232, O2233, O2234, O2235, O2236, O2237, O2238, O2239, O2240, O2241, O2242, O2243, O2244, O2245, O2246, O2247, O2248, O2249, O2250, O2251, O2252, O2253, O2254, O2255, O2256, O2257, O2258, O2259, O2260, O2261, O2262, O2263, O2264, O2265, O2266, O2267, O2268, O2269, O2270, O2271, O2272, O2273, O2274, O2275, O2276, O2277, O2278, O2279, O2280, O2281, O2282, O2283, O2284, O2285, O2286, O2287, O2288, O2289, O2290, O2291, O2292, O2293, O2294, O2295, O2296, O2297, O2298, O2299, O2300, O2301, O2302, O2303, O2304, O2305, O2306, O2307, O2308, O2309, O2310, O2311, O2312, O2313, O2314, O2315, O2316, O2317, O2318, O2319, O2320, O2321, O2322, O2323, O2324, O2325, O2326, O2327, O2328, O2329, O2330, O2331, O2332, O2333, O2334, O2335, O2336, O2337, O2338, O2339, O2340, O2341, O2342, O2343, O2344, O2345, O2346, O2347, O2348, O2349, O2350, O2351, O2352, O2353, O2354, O2355, O2356, O2357, O2358, O2359, O2360, O2361, O2362, O2363, O2364, O2365, O2366, O2367, O2368, O2369, O2370, O2371, O2372, O2373, O2374, O2375, O2376, O2377, O2378, O2379, O2380, O2381, O2382, O2383, O2384, O2385, O2386, O2387, O2388, O2389, O2390, O2391, O2392, O2393, O2394, O2395, O2396, O2397, O2398, O2399, O2400, O2401, O2402, O2403, O2404, O2405, O2406, O2407, O2408, O2409, O2410, O2411, O2412, O2413, O2414, O2415, O2416, O2417, O2418, O2419, O2420, O2421, O2422, O2423, O2424, O2425, O2426, O2427, O2428, O2429, O2430, O2431, O2432, O2433, O2434, O2435, O2436, O2437, O2438, O2439, O2440, O2441, O2442, O2443, O2444, O2445, O2446, O2447, O2448, O2449, O2450, O2451, O2452, O2453, O2454, O2455, O2456, O2457, O2458, O2459, O2460, O2461, O2462, O2463, O2464, O2465, O2466, O2467, O2468, O2469, O2470, O2471, O2472, O2473, O2474, O2475, O2476, O2477, O2478, O2479, O2480, O2481, O2482, O2483, O2484, O2485, O2486, O2487, O2488, O2489, O2490, O2491, O2492, O2493, O2494, O2495, O2496, O2497, O2498, O2499, O2500, O2501, O2502, O2503, O2504, O2505, O2506, O2507, O2508, O2509, O2510, O2511, O2512, O2513, O2514, O2515, O2516, O2517, O2518, O2519, O2520, O2521, O2522, O2523, O2524, O2525, O2526, O2527, O2528, O2529, O2530, O2531, O2532, O2533, O2534, O2535, O2536, O2537, O2538, O2539, O2540, O2541, O2542, O2543, O2544, O2545, O2546, O2547, O2548, O2549, O2550, O2551, O2552, O2553, O2554, O2555, O2556, O2557, O2558, O2559, O2560, O2561, O2562, O2563, O2564, O2565, O2566, O2567, O2568, O2569, O2570, O2571, O2572, O2573, O2574, O2575, O2576, O2577, O2578, O2579, O2580, O2581, O2582, O2583, O2584, O2585, O2586, O2587, O2588, O2589, O2590, O2591, O2592, O2593, O2594, O2595, O2596, O2597, O2598, O2599, O2600, O2601, O2602, O2603, O2604, O2605, O2606, O2607, O2608, O2609, O2610, O2611, O2612, O2613, O2614, O2615, O2616, O2617, O2618, O2619, O2620, O2621, O2622, O2623, O2624, O2625, O2626, O2627, O2628, O2629, O2630, O2631, O2632, O2633, O2634, O2635, O2636, O2637, O2638, O2639, O2640, O2641, O2642, O2643, O2644, O2645, O2646, O2647, O2648, O2649, O2650, O2651, O2652, O2653, O2654, O2655, O2656, O2657, O2658, O2659, O2660, O2661, O2662, O2663, O2664, O2665, O2666, O2667, O2668, O2669, O2670, O2671, O2672, O2673, O2674, O2675, O2676, O2677, O2678, O2679, O2680, O2681, O2682, O2683, O2684, O2685, O2686, O2687, O2688, O2689, O2690, O2691, O2692, O2693, O2694, O2695, O2696, O2697, O2698, O2699, O2700, O2701, O2702, O2703, O2704, O2705, O2706, O2707, O2708, O2709, O2710, O2711, O2712, O2713, O2714, O2715, O2716, O2717, O2718, O2719, O2720, O2721, O2722, O2723, O2724, O2725, O2726, O2727, O2728, O2729, O2730, O2731, O2732, O2733, O2734, O2735, O2736, O2737, O2738, O2739, O2740, O2741, O2742, O2743, O2744, O2745, O2746, O2747, O2748, O2749, O2750, O2751, O2752, O2753, O2754, O2755, O2756, O2757, O2758, O2759, O2760, O2761, O2762, O2763, O2764, O2765, O2766, O2767, O2768, O2769, O2770, O2771, O2772, O2773, O2774, O2775, O2776, O2777, O2778, O2779, O2780, O2781, O2782, O2783, O2784, O2785, O2786, O2787, O2788, O2789, O2790, O2791, O2792, O2793, O2794, O2795, O2796, O2797, O2798, O2799, O2800, O2801, O2802, O2803, O2804, O2805, O2806, O2807, O2808, O2809, O2810, O2811, O2812, O2813, O2814, O2815, O2816, O2817, O2818, O2819, O2820, O2821, O2822, O2823, O2824, O2825, O2826, O2827, O2828, O2829, O2830, O2831, O2832, O2833, O2834, O2835, O2836, O2837, O2838, O2839, O2840, O2841, O2842, O2843, O2844, O2845, O2846, O2847, O2848, O2849, O2850, O2851, O2852, O2853, O2854, O2855, O2856, O2857, O2858, O2859, O2860, O2861, O2862, O2863, O2864, O2865, O2866, O2867, O2868, O2869, O2870, O2871, O2872, O2873, O2874, O2875, O2876, O2877, O2878, O2879, O2880, O2881, O2882, O2883, O2884, O2885, O2886, O2887, O2888, O2889, O2890, O2891, O2892, O2893, O2894, O2895, O2896, O2897, O2898, O2899, O2900, O2901, O2902, O2903, O2904, O2905, O2906, O2907, O2908, O2909, O2910, O2911, O2912, O2913, O2914, O2915, O2916, O2917, O2918, O2919, O2920, O2921, O2922, O2923, O2924, O2925, O2926, O2927, O2928, O2929, O2930, O2931, O2932, O2933, O2934, O2935, O2936, O2937, O2938, O2939, O2940, O2941, O2942, O2943, O2944, O2945, O2946, O2947, O2948, O2949, O2950, O2951, O2952, O2953, O2954, O2955, O2956, O2957, O2958, O2959, O2960, O2961, O2962, O2963, O2964, O2965, O2966, O2967, O2968, O2969, O2970, O2971, O2972, O2973, O2974, O2975, O2976, O2977, O2978, O2979, O2980, O2981, O2982, O2983, O2984, O2985, O2986, O2987, O2988, O2989, O2990, O2991, O2992, O2993, O2994, O2995, O2996, O2997, O2998, O2999, O3000, O3001, O3002, O3003, O3004, O3005, O3006, O3007, O3008, O3009, O3010, O3011, O3012, O3013, O3014, O3015, O3016, O3017, O3018, O3019, O3020, O3021, O3022, O3023, O3024, O3025, O3026, O3027, O3028, O3029, O3030, O3031, O3032, O3033, O3034, O3035, O3036, O3037, O3038, O3039, O3040, O3041, O3042, O3043, O3044, O3045, O3046, O3047, O3048, O3049, O3050, O3051, O3052, O3053, O3054, O3055, O3056, O3057, O3058, O3059, O3060, O3061, O3062, O3063, O3064, O3065, O3066, O3067, O3068, O3069, O3070, O3071, O3072, O3073, O3074, O3075, O3076, O3077, O3078, O3079, O3080, O3081, O3082, O3083, O3084, O3085, O3086, O3087, O3088, O3089, O3090, O3091, O3092, O3093, O3094, O3095, O3096, O3097, O3098, O3099, O3100, O3101, O3102, O3103, O3104, O3105, O3106, O3107, O3108, O3109, O3110, O3111, O3112, O3113, O3114, O3115, O3116, O3117, O3118, O3119, O3120, O3121, O3122, O3123, O3124, O3125, O3126, O3127, O3128, O3129, O3130, O3131, O3132, O3133, O3134, O3135, O3136, O3137, O3138, O3139, O3140, O3141, O3142, O3143, O3144, O3145, O3146, O3147, O3148, O3149, O3150, O3151, O3152, O3153, O3154, O3155, O3156, O3157, O3158, O3159, O3160, O3161, O3162, O3163, O3164, O3165, O3166, O3167, O3168, O3169, O3170, O3171, O3172, O3173, O3174, O3175, O3176, O3177, O3178, O3179, O3180, O3181, O3182, O3183, O3184, O3185, O3186, O3187, O3188, O3189, O3190, O3191, O3192, O3193, O3194, O3195, O3196, O3197, O3198, O3199, O3200, O3201, O3202, O3203, O3204, O3205, O3206, O3207, O3208, O3209, O3210, O3211, O3212, O3213, O3214, O3215, O3216, O3217, O3218, O3219, O3220, O3221, O3222, O3223, O3224, O3225, O3226, O3227, O3228, O3229, O3230, O3231, O3232, O3233, O3234, O3235, O3236, O3237, O3238, O3239, O3240, O3241, O3242, O3243, O3244, O3245, O3246, O3247, O3248, O3249, O3250, O3251, O3252, O3253, O3254, O3255, O3256, O3257, O3258, O3259, O3260, O3261, O3262, O3263, O3264, O3265, O3266, O3267, O3268, O3269, O3270, O3271, O3272, O3273, O3274, O3275, O3276, O3277, O3278, O3279, O3280, O3281, O3282, O3283, O3284, O3285, O3286, O3287, O3288, O3289, O3290, O3291, O3292, O3293, O3294, O3295, O3296, O3297, O3298, O3299, O3300, O3301, O3302, O3303, O3304, O3305, O3306, O3307, O3308, O3309, O3310, O3311, O3312, O3313, O3314, O3315, O3316, O3317, O3318, O3319, O3320, O3321, O3322, O3323, O3324, O3325, O3326, O3327, O3328, O3329, O3330, O3331, O3332, O3333, O3334, O3335, O3336, O3337, O3338, O3339, O3340, O3341, O3342, O3343, O3344, O3345, O3346, O3347, O3348, O3349, O3350, O3351, O3352, O3353, O3354, O3355, O3356, O3357, O3358, O3359, O3360, O3361, O3362, O3363, O3364, O3365, O3366, O3367, O3368, O3369, O3370, O3371, O3372, O3373, O3374, O3375, O3376, O3377, O3378, O3379, O3380, O3381, O3382, O3383, O3384, O3385, O3386, O3387, O3388, O3389, O3390, O3391, O3392, O3393, O3394, O3395, O3396, O3397, O3398, O3399, O3400, O3401, O3402, O3403, O3404, O3405, O3406, O3407, O3408, O3409, O3410, O3411, O3412, O3413, O3414, O3415, O3416, O3417, O3418, O3419, O3420, O3421, O3422, O3423, O3424, O3425, O3426, O3427, O3428, O3429, O3430, O3431, O3432, O3433, O3434, O3435, O3436, O3437, O3438, O3439, O3440, O3441, O3442, O3443, O3444, O3445, O3446, O3447, O3448, O3449, O3450, O3451, O3452, O3453, O3454, O3455, O3456, O3457, O3458, O3459, O3460, O3461, O3462, O3463, O3464, O3465, O3466, O3467, O3468, O3469, O3470, O3471, O3472, O3473, O3474, O3475, O3476, O3477, O3478, O3479, O3480, O3481, O3482, O3483, O3484, O3485, O3486, O3487, O3488, O3489, O3490, O3491, O3492, O3493, O3494, O3495, O3496, O3497, O3498, O3499, O3500, O3501, O3502, O3503, O3504, O3505, O3506, O3507, O3508, O3509, O3510, O3511, O3512, O3513, O3514, O3515, O3516, O3517, O3518, O3519, O3520, O3521, O3522, O3523, O3524, O3525, O3526, O3527, O3528, O3529, O3530, O3531, O3532, O3533, O3534, O3535, O3536, O3537, O3538, O3539, O3540, O3541, O3542, O3543, O3544, O3545, O3546, O3547, O3548, O3549, O3550, O3551, O3552, O3553, O3554, O3555, O3556, O3557, O3558, O3559, O3560, O3561, O3562, O3563, O3564, O3565, O3566, O3567, O3568, O3569, O3570, O3571, O3572, O3573, O3574, O3575, O3576, O3577, O3578, O3579, O3580, O3581, O3582, O3583, O3584, O3585, O3586, O3587, O3588, O3589, O3590, O3591, O3592, O3593, O3594, O3595, O3596, O3597, O3598, O3599, O3600, O3601, O3602, O3603, O3604, O3605, O3606, O3607, O3608, O3609, O3610, O3611, O3612, O3613, O3614, O3615, O3616, O3617, O3618, O3619, O3620, O3621, O3622, O3623, O3624, O3625, O3626, O3627, O3628, O3629, O3630, O3631, O3632, O3633, O3634, O3635, O3636, O3637, O3638, O3639, O3640, O3641, O3642, O3643, O3644, O3645, O3646, O3647, O3648, O3649, O3650, O3651, O3652, O3653, O3654, O3655, O3656, O3657, O3658, O3659, O3660, O3661, O3662, O3663, O3664, O3665, O3666, O3667, O3668, O3669, O3670, O3671, O3672, O3673, O3674, O3675, O3676, O3677, O3678, O3679, O3680, O3681, O3682, O3683, O3684, O3685, O3686, O3687, O3688, O3689, O3690, O3691, O3692, O3693, O3694, O3695, O3696, O3697, O3698, O3699, O3700, O3701, O3702, O3703, O3704, O3705, O3706, O3707, O3708, O3709, O3710, O3711, O3712, O3713, O3714, O3715, O3716, O3717, O3718, O3719, O3720, O3721, O3722, O3723, O3724, O3725, O3726, O3727, O3728, O3729, O3730, O3731, O3732, O3733, O3734, O3735, O3736, O3737, O3738, O3739, O3740, O3741, O3742, O3743, O3744, O3745, O3746, O3747, O3748, O3749, O3750, O3751, O3752, O3753, O3754, O3755, O3756, O3757, O3758, O3759, O3760, O3761, O3762, O3763, O3764, O3765, O3766, O3767, O3768, O3769, O3770, O3771, O3772, O3773, O3774, O3775, O3776, O3777, O3778, O3779, O3780, O3781, O3782, O3783, O3784, O3785, O3786, O3787, O3788, O3789, O3790, O3791, O3792, O3793, O3794, O3795, O3796, O3797, O3798, O3799, O3800, O3801, O3802, O3803, O3804, O3805, O3806, O3807, O3808, O3809, O3810, O3811, O3812, O3813, O3814, O3815, O3816, O3817, O3818, O3819, O3820, O3821, O3822, O3823, O3824, O3825, O3826, O3827, O3828, O3829, O3830, O3831, O3832, O3833, O3834, O3835, O3836, O3837, O3838, O3839, O3840, O3841, O3842, O3843, O3844, O3845, O3846, O3847, O3848, O3849, O3850, O3851, O3852, O3853, O3854, O3855, O3856, O3857, O3858, O3859, O3860, O3861, O3862, O3863, O3864, O3865, O3866, O3867, O3868, O3869, O3870, O3871, O3872, O3873, O3874, O3875, O3876, O3877, O3878, O3879, O3880, O3881, O3882, O3883, O3884, O3885, O3886, O3887, O3888, O3889, O3890, O3891, O3892, O3893, O3894, O3895, O3896, O3897, O3898, O3899, O3900, O3901, O3902, O3903, O3904, O3905, O3906, O3907, O3908, O3909, O3910, O3911, O3912, O3913, O3914, O3915, O3916, O3917, O3918, O3919, O3920, O3921, O3922, O3923, O3924, O3925, O3926, O3927, O3928, O3929, O3930, O3931, O3932, O3933, O3934, O3935, O3936, O3937, O3938, O3939, O3940, O3941, O3942, O3943, O3944, O3945, O3946, O3947, O3948, O3949, O3950, O3951, O3952, O3953, O3954, O3955, O3956, O3957, O3958, O3959, O3960, O3961, O3962, O3963, O3964, O3965, O3966, O3967, O3968, O3969, O3970, O3971, O3972, O3973, O3974, O3975, O3976, O3977, O3978, O3979, O3980, O3981, O3982, O3983, O3984, O3985, O3986, O3987, O3988, O3989, O3990, O3991, O3992, O3993, O3994, O3995, O3996, O3997, O3998, O3999, O4000, O4001, O4002, O4003, O4004, O4005, O4006, O4007, O4008, O4009, O4010, O4011, O4012, O4013, O4014, O4015, O4016, O4017, O4018, O4019, O4020, O4021, O4022, O4023, O4024, O4025, O4026, O4027, O4028, O4029, O4030, O4031, O4032, O4033, O4034, O4035, O4036, O4037, O4038, O4039, O4040, O4041, O4042, O4043, O4044, O4045, O4046, O4047, O4048, O4049, O4050, O4051, O4052, O4053, O4054, O4055, O4056, O4057, O4058, O4059, O4060, O4061, O4062, O4063, O4064, O4065, O4066, O4067, O4068, O4069, O4070, O4071, O4072, O4073, O4074, O4075, O4076, O4077, O4078, O4079, O4080, O4081, O4082, O4083, O4084, O4085, O4086, O4087, O4088, O4089, O4090, O4091, O4092, O4093, O4094, O4095, O4096, O4097, O4098, O4099, O4100, O4101, O4102, O4103, O4104, O4105, O4106, O4107, O4108, O4109, O4110, O4111, O4112, O4113, O4114, O4115, O4116, O4117, O4118, O4119, O4120, O4121, O4122, O4123, O4124, O4125, O4126, O4127, O4128, O4129, O4130, O4131, O4132, O4133, O4134, O4135, O4136, O4137, O4138, O4139, O4140, O4141, O4142, O4143, O4144, O4145, O4146, O4147, O4148, O4149, O4150, O4151, O4152, O4153, O4154, O4155, O4156, O4157, O4158, O4159, O4160, O4161, O4162, O4163, O4164, O4165, O4166, O4167, O4168, O4169, O4170, O4171, O4172, O4173, O4174, O4175, O4176, O4177, O4178, O4179, O4180, O4181, O4182, O4183, O4184, O4185, O4186, O4187, O4188, O4189, O4190, O4191, O4192, O4193, O4194, O4195, O4196, O4197, O4198, O4199, O4200, O4201, O4202, O4203, O4204, O4205, O4206, O4207, O4208, O4209, O4210, O4211, O4212, O4213, O4214, O4215, O4216, O4217, O4218, O4219, O4220, O4221, O4222, O4223, O4224, O4225, O4226, O4227, O4228, O4229, O4230, O4231, O4232, O4233, O4234, O4235, O4236, O4237, O4238, O4239, O4240, O4241, O4242, O4243, O4244, O4245, O4246, O4247, O4248, O4249, O4250, O4251, O4252, O4253, O4254, O4255, O4256, O4257, O4258, O4259, O4260, O4261, O4262, O4263, O4264, O4265, O4266, O4267, O4268, O4269, O4270, O4271, O4272, O4273, O4274, O4275, O4276, O4277, O4278, O4279, O4280, O4281, O4282, O4283, O4284, O4285, O4286, O4287, O4288, O4289, O4290, O4291, O4292, O4293, O4294, O4295, O4296, O4297, O4298, O4299, O4300, O4301, O4302, O4303, O4304, O4305, O4306, O4307, O4308, O4309, O4310, O4311, O4312, O4313, O4314, O4315, O4316, O4317, O4318, O4319, O4320, O4321, O4322, O4323, O4324, O4325, O4326, O4327, O4328, O4329, O4330, O4331, O4332, O4333, O4334, O4335, O4336, O4337, O4338, O4339, O4340, O4341, O4342, O4343, O4344, O4345, O4346, O4347, O4348, O4349, O4350, O4351, O4352, O4353, O4354, O4355, O4356, O4357, O4358, O4359, O4360, O4361, O4362, O4363, O4364, O4365, O4366, O4367, O4368, O4369, O4370, O4371, O4372, O4373, O4374, O4375, O4376, O4377, O4378, O4379, O4380, O4381, O4382, O4383, O4384, O4385, O4386, O4387, O4388, O4389, O4390, O4391, O4392, O4393, O4394, O4395, O4396, O4397, O4398, O4399, O4400, O4401, O4402, O4403, O4404, O4405, O4406, O4407, O4408, O4409, O4410, O4411, O4412, O4413, O4414, O4415, O4416, O4417, O4418, O4419, O4420, O4421, O4422, O4423, O4424, O4425, O4426, O4427, O4428, O4429, O4430, O4431, O4432, O4433, O4434, O4435, O4436, O4437, O4438, O4439, O4440, O4441, O4442, O4443, O4444, O4445, O4446, O4447, O4448, O4449, O4450, O4451, O4452, O4453, O4454, O4455, O4456, O4457, O4458, O4459, O4460, O4461, O4462, O4463, O4464, O4465, O4466, O4467, O4468, O4469, O4470, O4471, O4472, O4473, O4474, O4475, O4476, O4477, O4478, O4479, O4480, O4481, O4482, O4483, O4484, O4485, O4486, O4487, O4488, O4489, O4490, O4491, O4492, O4493, O4494, O4495, O4496, O4497, O4498, O4499, O4500, O4501, O4502, O4503, O4504, O4505, O4506, O4507, O4508, O4509, O4510, O4511, O4512, O4513, O4514, O4515, O4516, O4517, O4518, O4519, O4520, O4521, O4522, O4523, O4524, O4525, O4526, O4527, O4528, O4529, O4530, O4531, O4532, O4533, O4534, O4535, O4536, O4537, O4538, O4539, O4540, O4541, O4542, O4543, O4544, O4545, O4546, O4547, O4548, O4549, O4550, O4551, O4552, O4553, O4554, O4555, O4556, O4557, O4558, O4559, O4560, O4561, O4562, O4563, O4564, O4565, O4566, O4567, O4568, O4569, O4570, O4571, O4572, O4573, O4574, O4575, O4576, O4577, O4578, O4579, O4580, O4581, O4582, O4583, O4584, O4585, O4586, O4587, O4588, O4589, O4590, O4591, O4592, O4593, O4594, O4595, O4596, O4597, O4598, O4599, O4600, O4601, O4602, O4603, O4604, O4605, O4606, O4607, O4608, O4609, O4610, O4611, O4612, O4613, O4614, O4615, O4616, O4617, O4618, O4619, O4620, O4621, O4622, O4623, O4624, O4625, O4626, O4627, O4628, O4629, O4630, O4631, O4632, O4633, O4634, O4635, O4636, O4637, O4638, O4639, O4640, O4641, O4642, O4643, O4644, O4645, O4646, O4647, O4648, O4649, O4650, O4651, O4652, O4653, O4654, O4655, O4656, O4657, O4658, O4659, O4660, O4661, O4662, O4663, O4664, O4665, O4666, O4667, O4668, O4669, O4670, O4671, O4672, O4673, O4674, O4675, O4676, O4677, O4678, O4679, O4680, O4681, O4682, O4683, O4684, O4685, O4686, O4687, O4688, O4689, O4690, O4691, O4692, O4693, O4694, O4695, O4696, O4697, O4698, O4699, O4700, O4701, O4702, O4703, O4704, O4705, O4706, O4707, O4708, O4709, O4710, O4711, O4712, O4713, O4714, O4715, O4716, O4717, O4718, O4719, O4720, O4721, O4722, O4723, O4724, O4725, O4726, O4727, O4728, O4729, O4730, O4731, O4732, O4733, O4734, O4735, O4736, O4737, O4738, O4739, O4740, O4741, O4742, O4743, O4744, O4745, O4746, O4747, O4748, O4749, O4750, O4751, O4752, O4753, O4754, O4755, O4756, O4757, O4758, O4759, O4760, O4761, O4762, O4763, O4764, O4765, O4766, O4767, O4768, O4769, O4770, O4771, O4772, O4773, O4774, O4775, O4776, O4777, O4778, O4779, O4780, O4781, O4782, O4783, O4784, O4785, O4786, O4787, O4788, O4789, O4790, O4791, O4792, O4793, O4794, O4795, O4796, O4797, O4798, O4799, O4800, O4801, O4802, O4803, O4804, O4805, O4806, O4807, O4808, O4809, O4810, O4811, O4812, O4813, O4814, O4815, O4816, O4817, O4818, O4819, O4820, O4821, O4822, O4823, O4824, O4825, O4826, O4827, O4828, O4829, O4830, O4831, O4832, O4833, O4834, O4835, O4836, O4837, O4838, O4839, O4840, O4841, O4842, O4843, O4844, O4845, O4846, O4847, O4848, O4849, O4850, O4851, O4852, O4853, O4854, O4855, O4856, O4857, O4858, O4859, O4860, O4861, O4862, O4863, O4864, O4865, O4866, O4867, O4868, O4869, O4870, O4871, O4872, O4873, O4874, O4875, O4876, O4877, O4878, O4879, O4880, O4881, O4882, O4883, O4884, O4885, O4886, O4887, O4888, O4889, O4890, O4891, O4892, O4893, O4894, O4895, O4896, O4897, O4898, O4899, O4900, O4901, O4902, O4903, O4904, O4905, O4906, O4907, O4908, O4909, O4910, O4911, O4912, O4913, O4914, O4915, O4916, O4917, O4918, O4919, O4920, O4921, O4922, O4923, O4924, O4925, O4926, O4927, O4928, O4929, O4930, O4931, O4932, O4933, O4934, O4935, O4936, O4937, O4938, O4939, O4940, O4941, O4942, O4943, O4944, O4945, O4946, O4947, O4948, O4949, O4950, O4951, O4952, O4953, O4954, O4955, O4956, O4957, O4958, O4959, O4960, O4961, O4962, O4963, O4964, O4965, O4966, O4967, O4968, O4969, O4970, O4971, O4972, O4973, O4974, O4975, O4976, O4977, O4978, O4979, O4980, O4981, O4982, O4983, O4984, O4985, O4986, O4987, O4988, O4989, O4990, O4991, O4992, O4993, O4994, O4995, O4996, O4997, O4998, O4999, O5000, O5001, O5002, O5003, O5004, O5005, O5006, O5007, O5008, O5009, O5010, O5011, O5012, O5013, O5014, O5015, O5016, O5017, O5018, O5019, O5020, O5021, O5022, O5023, O5024, O5025, O5026, O5027, O5028, O5029, O5030, O5031, O5032, O5033, O5034, O5035, O5036, O5037, O5038, O5039, O5040, O5041, O5042, O5043, O5044, O5045, O5046, O5047, O5048, O5049, O5050, O5051, O5052, O5053, O5054, O5055, O5056, O5057, O5058, O5059, O5060, O5061, O5062, O5063, O5064, O5065, O5066, O5067, O5068, O5069, O5070, O5071, O5072, O5073, O5074, O5075, O5076, O5077, O5078, O5079, O5080, O5081, O5082, O5083, O5084, O5085, O5086, O5087, O5088, O5089, O5090, O5091, O5092, O5093, O5094, O5095, O5096, O5097, O5098, O5099, O5100, O5101, O5102, O5103, O5104, O5105, O5106, O5107, O5108, O5109, O5110, O5111, O5112, O5113, O5114, O5115, O5116, O5117, O5118, O5119, O5120, O5121, O5122, O5123, O5124, O5125, O5126, O5127, O5128, O5129, O5130, O5131, O5132, O5133, O5134, O5135, O5136, O5137, O5138, O5139, O5140, O5141, O5142, O5143, O5144, O5145, O5146, O5147, O5148, O5149, O5150, O5151, O5152, O5153, O5154, O5155, O5156, O5157, O5158, O5159, O5160, O5161, O5162, O5163, O5164, O5165, O5166, O5167, O5168, O5169, O5170, O5171, O5172, O5173, O5174, O5175, O5176, O5177, O5178, O5179, O5180, O5181, O5182, O5183, O5184, O5185, O5186, O5187, O5188, O5189, O5190, O5191, O5192, O5193, O5194, O5195, O5196, O5197, O5198, O5199, O5200, O5201, O5202, O5203, O5204, O5205, O5206, O5207, O5208, O5209, O5210, O5211, O5212, O5213, O5214, O5215, O5216, O5217, O5218, O5219, O5220, O5221, O5222, O5223, O5224, O5225, O5226, O5227, O5228, O5229, O5230, O5231, O5232, O5233, O5234, O5235, O5236, O5237, O5238, O5239, O5240, O5241, O5242, O5243, O5244, O5245, O5246, O5247, O5248, O5249, O5250, O5251, O5252, O5253, O5254, O5255, O5256, O5257, O5258, O5259, O5260, O5261, O5262, O5263, O5264, O5265, O5266, O5267, O5268, O5269, O5270, O5271, O5272, O5273, O5274, O5275, O5276, O5277, O5278, O5279, O5280, O5281, O5282, O5283, O5284, O5285, O5286, O5287, O5288, O5289, O5290, O5291, O5292, O5293, O5294, O5295, O5296, O5297, O5298, O5299, O5300, O5301, O5302, O5303, O5304, O5305, O5306, O5307, O5308, O5309, O5310, O5311, O5312, O5313, O5314, O5315, O5316, O5317, O5318, O5319, O5320, O5321, O5322, O5323, O5324, O5325, O5326, O5327, O5328, O5329, O5330, O5331, O5332, O5333, O5334, O5335, O5336, O5337, O5338, O5339, O5340, O5341, O5342, O5343, O5344, O5345, O5346, O5347, O5348, O5349, O5350, O5351, O5352, O5353, O5354, O5355, O5356, O5357, O5358, O5359, O5360, O5361, O5362, O5363, O5364, O5365, O5366, O5367, O5368, O5369, O5370, O5371, O5372, O5373, O5374, O5375, O5376, O5377, O5378, O5379, O5380, O5381, O5382, O5383, O5384, O5385, O5386, O5387, O5388, O5389, O5390, O5391, O5392, O5393, O5394, O5395, O5396, O5397, O5398, O5399, O5400, O5401, O5402, O5403, O5404, O5405, O5406, O5407, O5408, O5409, O5410, O5411, O5412, O5413, O5414, O5415, O5416, O5417, O5418, O5419, O5420, O5421, O5422, O5423, O5424, O5425, O5426, O5427, O5428, O5429, O5430, O5431, O5432, O5433, O5434, O5435, O5436, O5437, O5438, O5439, O5440, O5441, O5442, O5443, O5444, O5445, O5446, O5447, O5448, O5449, O5450, O5451, O5452, O5453, O5454, O5455, O5456, O5457, O5458, O5459, O5460, O5461, O5462, O5463, O5464, O5465, O5466, O5467, O5468, O5469, O5470, O5471, O5472, O5473, O5474, O5475, O5476, O5477, O5478, O5479, O5480, O5481, O5482, O5483, O5484, O5485, O5486, O5487, O5488, O5489, O5490, O5491, O5492, O5493, O5494, O5495, O5496, O5497, O5498, O5499, O5500, O5501, O5502, O5503, O5504, O5505, O5506, O5507, O5508, O5509, O5510, O5511, O5512, O5513, O5514, O5515, O5516, O5517, O5518, O5519, O5520, O5521, O5522, O5523, O5524, O5525, O5526, O5527, O5528, O5529, O5530, O5531, O5532, O5533, O5534, O5535, O5536, O5537, O5538, O5539, O5540, O5541, O5542, O5543, O5544, O5545, O5546, O5547, O5548, O5549, O5550, O5551, O5552, O5553, O5554, O5555, O5556, O5557, O5558, O5559, O5560, O5561, O5562, O5563, O5564, O5565, O5566, O5567, O5568, O5569, O5570, O5571, O5572, O5573, O5574, O5575, O5576, O5577, O5578, O5579, O5580, O5581, O5582, O5583, O5584, O5585, O5586, O5587, O5588, O5589, O5590, O5591, O5592, O5593, O5594, O5595, O5596, O5597, O5598, O5599, O5600, O5601, O5602, O5603, O5604, O5605, O5606, O5607, O5608, O5609, O5610, O5611, O5612, O5613, O5614, O5615, O5616, O5617, O5618, O5619, O5620, O5621, O5622, O5623, O5624, O5625, O5626, O5627, O5628, O5629, O5630, O5631, O5632, O5633, O5634, O5635, O5636, O5637, O5638, O5639, O5640, O5641, O5642, O5643, O5644, O5645, O5646, O5647, O5648, O5649, O5650, O5651, O5652, O5653, O5654, O5655, O5656, O5657, O5658, O5659, O5660, O5661, O5662, O5663, O5664, O5665, O5666, O5667, O5668, O5669, O5670, O5671, O5672, O5673, O5674, O5675, O5676, O5677, O5678, O5679, O5680, O5681, O5682, O5683, O5684, O5685, O5686, O5687, O5688, O5689, O5690, O5691, O5692, O5693, O5694, O5695, O5696, O5697, O5698, O5699, O5700, O5701, O5702, O5703, O5704, O5705, O5706, O5707, O5708, O5709, O5710, O5711, O5712, O5713, O5714, O5715, O5716, O5717, O5718, O5719, O5720, O5721, O5722, O5723, O5724, O5725, O5726, O5727, O5728, O5729, O5730, O5731, O5732, O5733, O5734, O5735, O5736, O5737, O5738, O5739, O5740, O5741, O5742, O5743, O5744, O5745, O5746, O5747, O5748, O5749, O5750, O5751, O5752, O5753, O5754, O5755, O5756, O5757, O5758, O5759, O5760, O5761, O5762, O5763, O5764, O5765, O5766, O5767, O5768, O5769, O5770, O5771, O5772, O5773, O5774, O5775, O5776, O5777, O5778, O5779, O5780, O5781, O5782, O5783, O5784, O5785, O5786, O5787, O5788, O5789, O5790, O5791, O5792, O5793, O5794, O5795, O5796, O5797, O5798, O5799, O5800, O5801, O5802, O5803, O5804, O5805, O5806, O5807, O5808, O5809, O5810, O5811, O5812, O5813, O5814, O5815, O5816, O5817, O5818, O5819, O5820, O5821, O5822, O5823, O5824, O5825, O5826, O5827, O5828, O5829, O5830, O5831, O5832, O5833, O5834, O5835, O5836, O5837, O5838, O5839, O5840, O5841, O5842, O5843, O5844, O5845, O5846, O5847, O5848, O5849, O5850, O5851, O5852, O5853, O5854, O5855, O5856, O5857, O5858, O5859, O5860, O5861, O5862, O5863, O5864, O5865, O5866, O5867, O5868, O5869, O5870, O5871, O5872, O5873, O5874, O5875, O5876, O5877, O5878, O5879, O5880, O5881, O5882, O5883, O5884, O5885, O5886, O5887, O5888, O5889, O5890, O5891, O5892, O5893, O5894, O5895, O5896, O5897, O5898, O5899, O5900, O5901, O5902, O5903, O5904, O5905, O5906, O5907, O5908, O5909, O5910, O5911, O5912, O5913, O5914, O5915, O5916, O5917, O5918, O5919, O5920, O5921, O5922, O5923, O5924, O5925, O5926, O5927, O5928, O5929, O5930, O5931, O5932, O5933, O5934, O5935, O5936, O5937, O5938, O5939, O5940, O5941, O5942, O5943, O5944, O5945, O5946, O5947, O5948, O5949, O5950, O5951, O5952, O5953, O5954, O5955, O5956, O5957, O5958, O5959, O5960, O5961, O5962, O5963, O5964, O5965, O5966, O5967, O5968, O5969, O5970, O5971, O5972, O5973, O5974, O5975, O5976, O5977, O5978, O5979, O5980, O5981, O5982, O5983, O5984, O5985, O5986, O5987, O5988, O5989, O5990, O5991, O5992, O5993, O5994, O5995, O5996, O5997, O5998, O5999, O6000, O6001, O6002, O6003, O6004, O6005, O6006, O6007, O6008, O6009, O6010, O6011, O6012, O6013, O6014, O6015, O6016, O6017, O6018, O6019, O6020, O6021, O6022, O6023, O6024, O6025, O6026, O6027, O6028, O6029, O6030, O6031, O6032, O6033, O6034, O6035, O6036, O6037, O6038, O6039, O6040, O6041, O6042, O6043, O6044, O6045, O6046, O6047, O6048, O6049, O6050, O6051, O6052, O6053, O6054, O6055, O6056, O6057, O6058, O6059, O6060, O6061, O6062, O6063, O6064, O6065, O6066, O6067, O6068, O6069, O6070, O6071, O6072, O6073, O6074, O6075, O6076, O6077, O6078, O6079, O6080, O6081, O6082, O6083, O6084, O6085, O6086, O6087, O6088, O6089, O6090, O6091, O6092, O6093, O6094, O6095, O6096, O6097, O6098, O6099, O6100, O6101, O6102, O6103, O6104, O6105, O6106, O6107, O6108, O6109, O6110, O6111, O6112, O6113, O6114, O6115, O6116, O6117, O6118, O6119, O6120, O6121, O6122, O6123, O6124, O6125, O6126, O6127, O6128, O6129, O6130, O6131, O6132, O6133, O6134, O6135, O6136, O6137, O6138, O6139, O6140, O6141, O6142, O6143, O6144, O6145, O6146, O6147, O6148, O6149, O6150, O6151, O6152, O6153, O6154, O6155, O6156, O6157, O6158, O6159, O6160, O6161, O6162, O6163, O6164, O6165, O6166, O6167, O6168, O6169, O6170, O6171, O6172, O6173, O6174, O6175, O6176, O6177, O6178, O6179, O6180, O6181, O6182, O6183, O6184, O6185, O6186, O6187, O6188, O6189, O6190, O6191, O6192, O6193, O6194, O6195, O6196, O6197, O6198, O6199, O6200, O6201, O6202, O6203, O6204, O6205, O6206, O6207, O6208, O6209, O6210, O6211, O6212, O6213, O6214, O6215, O6216, O6217, O6218, O6219, O6220, O6221, O6222, O6223, O6224, O6225, O6226, O6227, O6228, O6229, O6230, O6231, O6232, O6233, O6234, O6235, O6236, O6237, O6238, O6239, O6240, O6241, O6242, O6243, O6244, O6245, O6246, O6247, O6248, O6249, O6250, O6251, O6252, O6253, O6254, O6255, O6256, O6257, O6258, O6259, O6260, O6261, O6262, O6263, O6264, O6265, O6266, O6267, O6268, O6269, O6270, O6271, O6272, O6273, O6274, O6275, O6276, O6277, O6278, O6279, O6280, O6281, O6282, O6283, O6284, O6285, O6286, O6287, O6288, O6289, O6290, O6291, O6292, O6293, O6294, O6295, O6296, O6297, O6298, O6299, O6300, O6301, O6302, O6303, O6304, O6305, O6306, O6307, O6308, O6309, O6310, O6311, O6312, O6313, O6314, O6315, O6316, O6317, O6318, O6319, O6320, O6321, O6322, O6323, O6324, O6325, O6326, O6327, O6328, O6329, O6330, O6331, O6332, O6333, O6334, O6335, O6336, O6337, O6338, O6339, O6340, O6341, O6342, O6343, O6344, O6345, O6346, O6347, O6348, O6349, O6350, O6351, O6352, O6353, O6354, O6355, O6356, O6357, O6358, O6359, O6360, O6361, O6362, O6363, O6364, O6365, O6366, O6367, O6368, O6369, O6370, O6371, O6372, O6373, O6374, O6375, O6376, O6377, O6378, O6379, O6380, O6381, O6382, O6383, O6384, O6385, O6386, O6387, O6388, O6389, O6390, O6391, O6392, O6393, O6394, O6395, O6396, O6397, O6398, O6399, O6400, O6401, O6402, O6403, O6404, O6405, O6406, O6407, O6408, O6409, O6410, O6411, O6412, O6413, O6414, O6415, O6416, O6417, O6418, O6419, O6420, O6421, O6422, O6423, O6424, O6425, O6426, O6427, O6428, O6429, O6430, O6431, O6432, O6433, O6434, O6435, O6436, O6437, O6438, O6439, O6440, O6441, O6442, O6443, O6444, O6445, O6446, O6447, O6448, O6449, O6450, O6451, O6452, O6453, O6454, O6455, O6456, O6457, O6458, O6459, O6460, O6461, O6462, O6463, O6464, O6465, O6466, O6467, O6468, O6469, O6470, O6471, O6472, O6473, O6474, O6475, O6476, O6477, O6478, O6479, O6480, O6481, O6482, O6483, O6484, O6485, O6486, O6487, O6488, O6489, O6490, O6491, O6492, O6493, O6494, O6495, O6496, O6497, O6498, O6499, O6500, O6501, O6502, O6503, O6504, O6505, O6506, O6507, O6508, O6509, O6510, O6511, O6512, O6513, O6514, O6515, O6516, O6517, O6518, O6519, O6520, O6521, O6522, O6523, O6524, O6525, O6526, O6527, O6528, O6529, O6530, O6531, O6532, O6533, O6534, O6535, O6536, O6537, O6538, O6539, O6540, O6541, O6542, O6543, O6544, O6545, O6546, O6547, O6548, O6549, O6550, O6551, O6552, O6553, O6554, O6555, O6556, O6557, O6558, O6559, O6560, O6561, O6562, O6563, O6564, O6565, O6566, O6567, O6568, O6569, O6570, O6571, O6572, O6573, O6574, O6575, O6576, O6577, O6578, O6579, O6580, O6581, O6582, O6583, O6584, O6585, O6586, O6587, O6588, O6589, O6590, O6591, O6592, O6593, O6594, O6595, O6596, O6597, O6598, O6599, O6600, O6601, O6602, O6603, O6604, O6605, O6606, O6607, O6608, O6609, O6610, O6611, O6612, O6613, O6614, O6615, O6616, O6617, O6618, O6619, O6620, O6621, O6622, O6623, O6624, O6625, O6626, O6627, O6628, O6629, O6630, O6631, O6632, O6633, O6634, O6635, O6636, O6637, O6638, O6639, O6640, O6641, O6642, O6643, O6644, O6645, O6646, O6647, O6648, O6649, O6650, O6651, O6652, O6653, O6654, O6655, O6656, O6657, O6658, O6659, O6660, O6661, O6662, O6663, O6664, O6665, O6666, O6667, O6668, O6669, O6670, O6671, O6672, O6673, O6674, O6675, O6676, O6677, O6678, O6679, O6680, O6681, O6682, O6683, O6684, O6685, O6686, O6687, O6688, O6689, O6690, O6691, O6692, O6693, O6694, O6695, O6696, O6697, O6698, O6699, O6700, O6701, O6702, O6703, O6704, O6705, O6706, O6707, O6708, O6709, O6710, O6711, O6712, O6713, O6714, O6715, O6716, O6717, O6718, O6719, O6720, O6721, O6722, O6723, O6724, O6725, O6726, O6727, O6728, O6729, O6730, O6731, O6732, O6733, O6734, O6735, O6736, O6737, O6738, O6739, O6740, O6741, O6742, O6743, O6744, O6745, O6746, O6747, O6748, O6749, O6750, O6751, O6752, O6753, O6754, O6755, O6756, O6757, O6758, O6759, O6760, O6761, O6762, O6763, O6764, O6765, O6766, O6767, O6768, O6769, O6770, O6771, O6772, O6773, O6774, O6775, O6776, O6777, O6778, O6779, O6780, O6781, O6782, O6783, O6784, O6785, O6786, O6787, O6788, O6789, O6790, O6791, O6792, O6793, O6794, O6795, O6796, O6797, O6798, O6799, O6800, O6801, O6802, O6803, O6804, O6805, O6806, O6807, O6808, O6809, O6810, O6811, O6812, O6813, O6814, O6815, O6816, O6817, O6818, O6819, O6820, O6821, O6822, O6823, O6824, O6825, O6826, O6827, O6828, O6829, O6830, O6831, O6832, O6833, O6834, O6835, O6836, O6837, O6838, O6839, O6840, O6841, O6842, O6843, O6844, O6845, O6846, O6847, O6848, O6849, O6850, O6851, O6852, O6853, O6854, O6855, O6856, O6857, O6858, O6859, O6860, O6861, O6862, O6863, O6864, O6865, O6866, O6867, O6868, O6869, O6870, O6871, O6872, O6873, O6874, O6875, O6876, O6877, O6878, O6879, O6880, O6881, O6882, O6883, O6884, O6885, O6886, O6887, O6888, O6889, O6890, O6891, O6892, O6893, O6894, O6895, O6896, O6897, O6898, O6899, O6900, O6901, O6902, O6903, O6904, O6905, O6906, O6907, O6908, O6909, O6910, O6911, O6912, O6913, O6914, O6915, O6916, O6917, O6918, O6919, O6920, O6921, O6922, O6923, O6924, O6925, O6926, O6927, O6928, O6929, O6930, O6931, O6932, O6933, O6934, O6935, O6936, O6937, O6938, O6939, O6940, O6941, O6942, O6943, O6944, O6945, O6946, O6947, O6948, O6949, O6950, O6951, O6952, O6953, O6954, O6955, O6956, O6957, O6958, O6959, O6960, O6961, O6962, O6963, O6964, O6965, O6966, O6967, O6968, O6969, O6970, O6971, O6972, O6973, O6974, O6975, O6976, O6977, O6978, O6979, O6980, O6981, O6982, O6983, O6984, O6985, O6986, O6987, O6988, O6989, O6990, O6991, O6992, O6993, O6994, O6995, O6996, O6997, O6998, O6999, O7000, O7001, O7002, O7003, O7004, O7005, O7006, O7007, O7008, O7009, O7010, O7011, O7012, O7013, O7014, O7015, O7016, O7017, O7018, O7019, O7020, O7021, O7022, O7023, O7024, O7025, O7026, O7027, O7028, O7029, O7030, O7031, O7032, O7033, O7034, O7035, O7036, O7037, O7038, O7039, O7040, O7041, O7042, O7043, O7044, O7045, O7046, O7047, O7048, O7049, O7050, O7051, O7052, O7053, O7054, O7055, O7056, O7057, O7058, O7059, O7060, O7061, O7062, O7063, O7064, O7065, O7066, O7067, O7068, O7069, O7070, O7071, O7072, O7073, O7074, O7075, O7076, O7077, O7078, O7079, O7080, O7081, O7082, O7083, O7084, O7085, O7086, O7087, O7088, O7089, O7090, O7091, O7092, O7093, O7094, O7095, O7096, O7097, O7098, O7099, O7100, O7101, O7102, O7103, O7104, O7105, O7106, O7107, O7108, O7109, O7110, O7111, O7112, O7113, O7114, O7115, O7116, O7117, O7118, O7119, O7120, O7121, O7122, O7123, O7124, O7125, O7126, O7127, O7128, O7129, O7130, O7131, O7132, O7133, O7134, O7135, O7136, O7137, O7138, O7139, O7140, O7141, O7142, O7143, O7144, O7145, O7146, O7147, O7148, O7149, O7150, O7151, O7152, O7153, O7154, O7155, O7156, O7157, O7158, O7159, O7160, O7161, O7162, O7163, O7164, O7165, O7166, O7167, O7168, O7169, O7170, O7171, O7172, O7173, O7174, O7175, O7176, O7177, O7178, O7179, O7180, O7181, O7182, O7183, O7184, O7185, O7186, O7187, O7188, O7189, O7190, O7191, O7192, O7193, O7194, O7195, O7196, O7197, O7198, O7199, O7200, O7201, O7202, O7203, O7204, O7205, O7206, O7207, O7208, O7209, O7210, O7211, O7212, O7213, O7214, O7215, O7216, O7217, O7218, O7219, O7220, O7221, O7222, O7223, O7224, O7225, O7226, O7227, O7228, O7229, O7230, O7231, O7232, O7233, O7234, O7235, O7236, O7237, O7238, O7239, O7240, O7241, O7242, O7243, O7244, O7245, O7246, O7247, O7248, O7249, O7250, O7251, O7252, O7253, O7254, O7255, O7256, O7257, O7258, O7259, O7260, O7261, O7262, O7263, O7264, O7265, O7266, O7267, O7268, O7269, O7270, O7271, O7272, O7273, O7274, O7275, O7276, O7277, O7278, O7279, O7280, O7281, O7282, O7283, O7284, O7285, O7286, O7287, O7288, O7289, O7290, O7291, O7292, O7293, O7294, O7295, O7296, O7297, O7298, O7299, O7300, O7301, O7302, O7303, O7304, O7305, O7306, O7307, O7308, O7309, O7310, O7311, O7312, O7313, O7314, O7315, O7316, O7317, O7318, O7319, O7320, O7321, O7322, O7323, O7324, O7325, O7326, O7327, O7328, O7329, O7330, O7331, O7332, O7333, O7334, O7335, O7336, O7337, O7338, O7339, O7340, O7341, O7342, O7343, O7344, O7345, O7346, O7347, O7348, O7349, O7350, O7351, O7352, O7353, O7354, O7355, O7356, O7357, O7358, O7359, O7360, O7361, O7362, O7363, O7364, O7365, O7366, O7367, O7368, O7369, O7370, O7371, O7372, O7373, O7374, O7375, O7376, O7377, O7378, O7379, O7380, O7381, O7382, O7383, O7384, O7385, O7386, O7387, O7388, O7389, O7390, O7391, O7392, O7393, O7394, O7395, O7396, O7397, O7398, O7399, O7400, O7401, O7402, O7403, O7404, O7405, O7406, O7407, O7408, O7409, O7410, O7411, O7412, O7413, O7414, O7415, O7416, O7417, O7418, O7419, O7420, O7421, O7422, O7423, O7424, O7425, O7426, O7427, O7428, O7429, O7430, O7431, O7432, O7433, O7434, O7435, O7436, O7437, O7438, O7439, O7440, O7441, O7442, O7443, O7444, O7445, O7446, O7447, O7448, O7449, O7450, O7451, O7452, O7453, O7454, O7455, O7456, O7457, O7458, O7459, O7460, O7461, O7462, O7463, O7464, O7465, O7466, O7467, O7468, O7469, O7470, O7471, O7472, O7473, O7474, O7475, O7476, O7477, O7478, O7479, O7480, O7481, O7482, O7483, O7484, O7485, O7486, O7487, O7488, O7489, O7490, O7491, O7492, O7493, O7494, O7495, O7496, O7497, O7498, O7499, O7500, O7501, O7502, O7503, O7504, O7505, O7506, O7507, O7508, O7509, O7510, O7511, O7512, O7513, O7514, O7515, O7516, O7517, O7518, O7519, O7520, O7521, O7522, O7523, O7524, O7525, O7526, O7527, O7528, O7529, O7530, O7531, O7532, O7533, O7534, O7535, O7536, O7537, O7538, O7539, O7540, O7541, O7542, O7543, O7544, O7545, O7546, O7547, O7548, O7549, O7550, O7551, O7552, O7553, O7554, O7555, O7556, O7557, O7558, O7559, O7560, O7561, O7562, O7563, O7564, O7565, O7566, O7567, O7568, O7569, O7570, O7571, O7572, O7573, O7574, O7575, O7576, O7577, O7578, O7579, O7580, O7581, O7582, O7583, O7584, O7585, O7586, O7587, O7588, O7589, O7590, O7591, O7592, O7593, O7594, O7595, O7596, O7597, O7598, O7599, O7600, O7601, O7602, O7603, O7604, O7605, O7606, O7607, O7608, O7609, O7610, O7611, O7612, O7613, O7614, O7615, O7616, O7617, O7618, O7619, O7620, O7621, O7622, O7623, O7624, O7625, O7626, O7627, O7628, O7629, O7630, O7631, O7632, O7633, O7634, O7635, O7636, O7637, O7638, O7639, O7640, O7641, O7642, O7643, O7644, O7645, O7646, O7647, O7648, O7649, O7650, O7651, O7652, O7653, O7654, O7655, O7656, O7657, O7658, O7659, O7660, O7661, O7662, O7663, O7664, O7665, O7666, O7667, O7668, O7669, O7670, O7671, O7672, O7673, O7674, O7675, O7676, O7677, O7678, O7679, O7680, O7681, O7682, O7683, O7684, O7685, O7686, O7687, O7688, O7689, O7690, O7691, O7692, O7693, O7694, O7695, O7696, O7697, O7698, O7699, O7700, O7701, O7702, O7703, O7704, O7705, O7706, O7707, O7708, O7709, O7710, O7711, O7712, O7713, O7714, O7715, O7716, O7717, O7718, O7719, O7720, O7721, O7722, O7723, O7724, O7725, O7726, O7727, O7728, O7729, O7730, O7731, O7732, O7733, O7734, O7735, O7736, O7737, O7738, O7739, O7740, O7741, O7742, O7743, O7744, O7745, O7746, O7747, O7748, O7749, O7750, O7751, O7752, O7753, O7754, O7755, O7756, O7757, O7758, O7759, O7760, O7761, O7762, O7763, O7764, O7765, O7766, O7767, O7768, O7769, O7770, O7771, O7772, O7773, O7774, O7775, O7776, O7777, O7778, O7779, O7780, O7781, O7782, O7783, O7784, O7785, O7786, O7787, O7788, O7789, O7790, O7791, O7792, O7793, O7794, O7795, O7796, O7797, O7798, O7799, O7800, O7801, O7802, O7803, O7804, O7805, O7806, O7807, O7808, O7809, O7810, O7811, O7812, O7813, O7814, O7815, O7816, O7817, O7818, O7819, O7820, O7821, O7822, O7823, O7824, O7825, O7826, O7827, O7828, O7829, O7830, O7831, O7832, O7833, O7834, O7835, O7836, O7837, O7838, O7839, O7840, O7841, O7842, O7843, O7844, O7845, O7846, O7847, O7848, O7849, O7850, O7851, O7852, O7853, O7854, O7855, O7856, O7857, O7858, O7859, O7860, O7861, O7862, O7863, O7864, O7865, O7866, O7867, O7868, O7869, O7870, O7871, O7872, O7873, O7874, O7875, O7876, O7877, O7878, O7879, O7880, O7881, O7882, O7883, O7884, O7885, O7886, O7887, O7888, O7889, O7890, O7891, O7892, O7893, O7894, O7895, O7896, O7897, O7898, O7899, O7900, O7901, O7902, O7903, O7904, O7905, O7906, O7907, O7908, O7909, O7910, O7911, O7912, O7913, O7914, O7915, O7916, O7917, O7918, O7919, O7920, O7921, O7922, O7923, O7924, O7925, O7926, O7927, O7928, O7929, O7930, O7931, O7932, O7933, O7934, O7935, O7936, O7937, O7938, O7939, O7940, O7941, O7942, O7943, O7944, O7945, O7946, O7947, O7948, O7949, O7950, O7951, O7952, O7953, O7954, O7955, O7956, O7957, O7958, O7959, O7960, O7961, O7962, O7963, O7964, O7965, O7966, O7967, O7968, O7969, O7970, O7971, O7972, O7973, O7974, O7975, O7976, O7977, O7978, O7979, O7980, O7981, O7982, O7983, O7984, O7985, O7986, O7987, O7988, O7989, O7990, O7991, O7992, O7993, O7994, O7995, O7996, O7997, O7998, O7999, O8000, O8001, O8002, O8003, O8004, O8005, O8006, O8007, O8008, O8009, O8010, O8011, O8012, O8013, O8014, O8015, O8016, O8017, O8018, O8019, O8020, O8021, O8022, O8023, O8024, O8025, O8026, O8027, O8028, O8029, O8030, O8031, O8032, O8033, O8034, O8035, O8036, O8037, O8038, O8039, O8040, O8041, O8042, O8043, O8044, O8045, O8046, O8047, O8048, O8049, O8050, O8051, O8052, O8053, O8054, O8055, O8056, O8057, O8058, O8059, O8060, O8061, O8062, O8063, O8064, O8065, O8066, O8067, O8068, O8069, O8070, O8071, O8072, O8073, O8074, O8075, O8076, O8077, O8078, O8079, O8080, O8081, O8082, O8083, O8084, O8085, O8086, O8087, O8088, O8089, O8090, O8091, O8092, O8093, O8094, O8095, O8096, O8097, O8098, O8099, O8100, O8101, O8102, O8103, O8104, O8105, O8106, O8107, O8108, O8109, O8110, O8111, O8112, O8113, O8114, O8115, O8116, O8117, O8118, O8119, O8120, O8121, O8122, O8123, O8124, O8125, O8126, O8127, O8128, O8129, O8130, O8131, O8132, O8133, O8134, O8135, O8136, O8137, O8138, O8139, O8140, O8141, O8142, O8143, O8144, O8145, O8146, O8147, O8148, O8149, O8150, O8151, O8152, O8153, O8154, O8155, O8156, O8157, O8158, O8159, O8160, O8161, O8162, O8163, O8164, O8165, O8166, O8167, O8168, O8169, O8170, O8171, O8172, O8173, O8174, O8175, O8176, O8177, O8178, O8179, O8180, O8181, O8182, O8183, O8184, O8185, O8186, O8187, O8188, O8189, O8190, O8191, O8192, O8193, O8194, O8195, O8196, O8197, O8198, O8199, O8200, O8201, O8202, O8203, O8204, O8205, O8206, O8207, O8208, O8209, O8210, O8211, O8212, O8213, O8214, O8215, O8216, O8217, O8218, O8219, O8220, O8221, O8222, O8223, O8224, O8225, O8226, O8227, O8228, O8229, O8230, O8231, O8232, O8233, O8234, O8235, O8236, O8237, O8238, O8239, O8240, O8241, O8242, O8243, O8244, O8245, O8246, O8247, O8248, O8249, O8250, O8251, O8252, O8253, O8254, O8255, O8256, O8257, O8258, O8259, O8260, O8261, O8262, O8263, O8264, O8265, O8266, O8267, O8268, O8269, O8270, O8271, O8272, O8273, O8274, O8275, O8276, O8277, O8278, O8279, O8280, O8281, O8282, O8283, O8284, O8285, O8286, O8287, O8288, O8289, O8290, O8291, O8292, O8293, O8294, O8295, O8296, O8297, O8298, O8299, O8300, O8301, O8302, O8303, O8304, O8305, O8306, O8307, O8308, O8309, O8310, O8311, O8312, O8313, O8314, O8315, O8316, O8317, O8318, O8319, O8320, O8321, O8322, O8323, O8324, O8325, O8326, O8327, O8328, O8329, O8330, O8331, O8332, O8333, O8334, O8335, O8336, O8337, O8338, O8339, O8340, O8341, O8342, O8343, O8344, O8345, O8346, O8347, O8348, O8349, O8350, O8351, O8352, O8353, O8354, O8355, O8356, O8357, O8358, O8359, O8360, O8361, O8362, O8363, O8364, O8365, O8366, O8367, O8368, O8369, O8370, O8371, O8372, O8373, O8374, O8375, O8376, O8377, O8378, O8379, O8380, O8381, O8382, O8383, O8384, O8385, O8386, O8387, O8388, O8389, O8390, O8391, O8392, O8393, O8394, O8395, O8396, O8397, O8398, O8399, O8400, O8401, O8402, O8403, O8404, O8405, O8406, O8407, O8408, O8409, O8410, O8411, O8412, O8413, O8414, O8415, O8416, O8417, O8418, O8419, O8420, O8421, O8422, O8423, O8424, O8425, O8426, O8427, O8428, O8429, O8430, O8431, O8432, O8433, O8434, O8435, O8436, O8437, O8438, O8439, O8440, O8441, O8442, O8443, O8444, O8445, O8446, O8447, O8448, O8449, O8450, O8451, O8452, O8453, O8454, O8455, O8456, O8457, O8458, O8459, O8460, O8461, O8462, O8463, O8464, O8465, O8466, O8467, O8468, O8469, O8470, O8471, O8472, O8473, O8474, O8475, O8476, O8477, O8478, O8479, O8480, O8481, O8482, O8483, O8484, O8485, O8486, O8487, O8488, O8489, O8490, O8491, O8492, O8493, O8494, O8495, O8496, O8497, O8498, O8499, O8500, O8501, O8502, O8503, O8504, O8505, O8506, O8507, O8508, O8509, O8510, O8511, O8512, O8513, O8514, O8515, O8516, O8517, O8518, O8519, O8520, O8521, O8522, O8523, O8524, O8525, O8526, O8527, O8528, O8529, O8530, O8531, O8532, O8533, O8534, O8535, O8536, O8537, O8538, O8539, O8540, O8541, O8542, O8543, O8544, O8545, O8546, O8547, O8548, O8549, O8550, O8551, O8552, O8553, O8554, O8555, O8556, O8557, O8558, O8559, O8560, O8561, O8562, O8563, O8564, O8565, O8566, O8567, O8568, O8569, O8570, O8571, O8572, O8573, O8574, O8575, O8576, O8577, O8578, O8579, O8580, O8581, O8582, O8583, O8584, O8585, O8586, O8587, O8588, O8589, O8590, O8591, O8592, O8593, O8594, O8595, O8596, O8597, O8598, O8599, O8600, O8601, O8602, O8603, O8604, O8605, O8606, O8607, O8608, O8609, O8610, O8611, O8612, O8613, O8614, O8615, O8616, O8617, O8618, O8619, O8620, O8621, O8622, O8623, O8624, O8625, O8626, O8627, O8628, O8629, O8630, O8631, O8632, O8633, O8634, O8635, O8636, O8637, O8638, O8639, O8640, O8641, O8642, O8643, O8644, O8645, O8646, O8647, O8648, O8649, O8650, O8651, O8652, O8653, O8654, O8655, O8656, O8657, O8658, O8659, O8660, O8661, O8662, O8663, O8664, O8665, O8666, O8667, O8668, O8669, O8670, O8671, O8672, O8673, O8674, O8675, O8676, O8677, O8678, O8679, O8680, O8681, O8682, O8683, O8684, O8685, O8686, O8687, O8688, O8689, O8690, O8691, O8692, O8693, O8694, O8695, O8696, O8697, O8698, O8699, O8700, O8701, O8702, O8703, O8704, O8705, O8706, O8707, O8708, O8709, O8710, O8711, O8712, O8713, O8714, O8715, O8716, O8717, O8718, O8719, O8720, O8721, O8722, O8723, O8724, O8725, O8726, O8727, O8728, O8729, O8730, O8731, O8732, O8733, O8734, O8735, O8736, O8737, O8738, O8739, O8740, O8741, O8742, O8743, O8744, O8745, O8746, O8747, O8748, O8749, O8750, O8751, O8752, O8753, O8754, O8755, O8756, O8757, O8758, O8759, O8760, O8761, O8762, O8763, O8764, O8765, O8766, O8767, O8768, O8769, O8770, O8771, O8772, O8773, O8774, O8775, O8776, O8777, O8778, O8779, O8780, O8781, O8782, O8783, O8784, O8785, O8786, O8787, O8788, O8789, O8790, O8791, O8792, O8793, O8794, O8795, O8796, O8797, O8798, O8799, O8800, O8801, O8802, O8803, O8804, O8805, O8806, O8807, O8808, O8809, O8810, O8811, O8812, O8813, O8814, O8815, O8816, O8817, O8818, O8819, O8820, O8821, O8822, O8823, O8824, O8825, O8826, O8827, O8828, O8829, O8830, O8831, O8832, O8833, O8834, O8835, O8836, O8837, O8838, O8839, O8840, O8841, O8842, O8843, O8844, O8845, O8846, O8847, O8848, O8849, O8850, O8851, O8852, O8853, O8854, O8855, O8856, O8857, O8858, O8859, O8860, O8861, O8862, O8863, O8864, O8865, O8866, O8867, O8868, O8869, O8870, O8871, O8872, O8873, O8874, O8875, O8876, O8877, O8878, O8879, O8880, O8881, O8882, O8883, O8884, O8885, O8886, O8887, O8888, O8889, O8890, O8891, O8892, O8893, O8894, O8895, O8896, O8897, O8898, O8899, O8900, O8901, O8902, O8903, O8904, O8905, O8906, O8907, O8908, O8909, O8910, O8911, O8912, O8913, O8914, O8915, O8916, O8917, O8918, O8919, O8920, O8921, O8922, O8923, O8924, O8925, O8926, O8927, O8928, O8929, O8930, O8931, O8932, O8933, O8934, O8935, O8936, O8937, O8938, O8939, O8940, O8941, O8942, O8943, O8944, O8945, O8946, O8947, O8948, O8949, O8950, O8951, O8952, O8953, O8954, O8955, O8956, O8957, O8958, O8959, O8960, O8961, O8962, O8963, O8964, O8965, O8966, O8967, O8968, O8969, O8970, O8971, O8972, O8973, O8974, O8975, O8976, O8977, O8978, O8979, O8980, O8981, O8982, O8983, O8984, O8985, O8986, O8987, O8988, O8989, O8990, O8991, O8992, O8993, O8994, O8995, O8996, O8997, O8998, O8999, O9000, O9001, O9002, O9003, O9004, O9005, O9006, O9007, O9008, O9009, O9010, O9011, O9012, O9013, O9014, O9015, O9016, O9017, O9018, O9019, O9020, O9021, O9022, O9023, O9024, O9025, O9026, O9027, O9028, O9029, O9030, O9031, O9032, O9033, O9034, O9035, O9036, O9037, O9038, O9039, O9040, O9041, O9042, O9043, O9044, O9045, O9046, O9047, O9048, O9049, O9050, O9051, O9052, O9053, O9054, O9055, O9056, O9057, O9058, O9059, O9060, O9061, O9062, O9063, O9064, O9065, O9066, O9067, O9068, O9069, O9070, O9071, O9072, O9073, O9074, O9075, O9076, O9077, O9078, O9079, O9080, O9081, O9082, O9083, O9084, O9085, O9086, O9087, O9088, O9089, O9090, O9091, O9092, O9093, O9094, O9095, O9096, O9097, O9098, O9099, O9100, O9101, O9102, O9103, O9104, O9105, O9106, O9107, O9108, O9109, O9110, O9111, O9112, O9113, O9114, O9115, O9116, O9117, O9118, O9119, O9120, O9121, O9122, O9123, O9124, O9125, O9126, O9127, O9128, O9129, O9130, O9131, O9132, O9133, O9134, O9135, O9136, O9137, O9138, O9139, O9140, O9141, O9142, O9143, O9144, O9145, O9146, O9147, O9148, O9149, O9150, O9151, O9152, O9153, O9154, O9155, O9156, O9157, O9158, O9159, O9160, O9161, O9162, O9163, O9164, O9165, O9166, O9167, O9168, O9169, O9170, O9171, O9172, O9173, O9174, O9175, O9176, O9177, O9178, O9179, O9180, O9181, O9182, O9183, O9184, O9185, O9186, O9187, O9188, O9189, O9190, O9191, O9192, O9193, O9194, O9195, O9196, O9197, O9198, O9199, O9200, O9201, O9202, O9203, O9204, O9205, O9206, O9207, O9208, O9209, O9210, O9211, O9212, O9213, O9214, O9215, O9216, O9217, O9218, O9219, O9220, O9221, O9222, O9223, O9224, O9225, O9226, O9227, O9228, O9229, O9230, O9231, O9232, O9233, O9234, O9235, O9236, O9237, O9238, O9239, O9240, O9241, O9242, O9243, O9244, O9245, O9246, O9247, O9248, O9249, O9250, O9251, O9252, O9253, O9254, O9255, O9256, O9257, O9258, O9259, O9260, O9261, O9262, O9263, O9264, O9265, O9266, O9267, O9268, O9269, O9270, O9271, O9272, O9273, O9274, O9275, O9276, O9277, O9278, O9279, O9280, O9281, O9282, O9283, O9284, O9285, O9286, O9287, O9288, O9289, O9290, O9291, O9292, O9293, O9294, O9295, O9296, O9297, O9298, O9299, O9300, O9301, O9302, O9303, O9304, O9305, O9306, O9307, O9308, O9309, O9310, O9311, O9312, O9313, O9314, O9315, O9316, O9317, O9318, O9319, O9320, O9321, O9322, O9323, O9324, O9325, O9326, O9327, O9328, O9329, O9330, O9331, O9332, O9333, O9334, O9335, O9336, O9337, O9338, O9339, O9340, O9341, O9342, O9343, O9344, O9345, O9346, O9347, O9348, O9349, O9350, O9351, O9352, O9353, O9354, O9355, O9356, O9357, O9358, O9359, O9360, O9361, O9362, O9363, O9364, O9365, O9366, O9367, O9368, O9369, O9370, O9371, O9372, O9373, O9374, O9375, O9376, O9377, O9378, O9379, O9380, O9381, O9382, O9383, O9384, O9385, O9386, O9387, O9388, O9389, O9390, O9391, O9392, O9393, O9394, O9395, O9396, O9397, O9398, O9399, O9400, O9401, O9402, O9403, O9404, O9405, O9406, O9407, O9408, O9409, O9410, O9411, O9412, O9413, O9414, O9415, O9416, O9417, O9418, O9419, O9420, O9421, O9422, O9423, O9424, O9425, O9426, O9427, O9428, O9429, O9430, O9431, O9432, O9433, O9434, O9435, O9436, O9437, O9438, O9439, O9440, O9441, O9442, O9443, O9444, O9445, O9446, O9447, O9448, O9449, O9450, O9451, O9452, O9453, O9454, O9455, O9456, O9457, O9458, O9459, O9460, O9461, O9462, O9463, O9464, O9465, O9466, O9467, O9468, O9469, O9470, O9471, O9472, O9473, O9474, O9475, O9476, O9477, O9478, O9479, O9480, O9481, O9482, O9483, O9484, O9485, O9486, O9487, O9488, O9489, O9490, O9491, O9492, O9493, O9494, O9495, O9496, O9497, O9498, O9499, O9500, O9501, O9502, O9503, O9504, O9505, O9506, O9507, O9508, O9509, O9510, O9511, O9512, O9513, O9514, O9515, O9516, O9517, O9518, O9519, O9520, O9521, O9522, O9523, O9524, O9525, O9526, O9527, O9528, O9529, O9530, O9531, O9532, O9533, O9534, O9535, O9536, O9537, O9538, O9539, O9540, O9541, O9542, O9543, O9544, O9545, O9546, O9547, O9548, O9549, O9550, O9551, O9552, O9553, O9554, O9555, O9556, O9557, O9558, O9559, O9560, O9561, O9562, O9563, O9564, O9565, O9566, O9567, O9568, O9569, O9570, O9571, O9572, O9573, O9574, O9575, O9576, O9577, O9578, O9579, O9580, O9581, O9582, O9583, O9584, O9585, O9586, O9587, O9588, O9589, O9590, O9591, O9592, O9593, O9594, O9595, O9596, O9597, O9598, O9599, O9600, O9601, O9602, O9603, O9604, O9605, O9606, O9607, O9608, O9609, O9610, O9611, O9612, O9613, O9614, O9615, O9616, O9617, O9618, O9619, O9620, O9621, O9622, O9623, O9624, O9625, O9626, O9627, O9628, O9629, O9630, O9631, O9632, O9633, O9634, O9635, O9636, O9637, O9638, O9639, O9640, O9641, O9642, O9643, O9644, O9645, O9646, O9647, O9648, O9649, O9650, O9651, O9652, O9653, O9654, O9655, O9656, O9657, O9658, O9659, O9660, O9661, O9662, O9663, O9664, O9665, O9666, O9667, O9668, O9669, O9670, O9671, O9672, O9673, O9674, O9675, O9676, O9677, O9678, O9679, O9680, O9681, O9682, O9683, O9684, O9685, O9686, O9687, O9688, O9689, O9690, O9691, O9692, O9693, O9694, O9695, O9696, O9697, O9698, O9699, O9700, O9701, O9702, O9703, O9704, O9705, O9706, O9707, O9708, O9709, O9710, O9711, O9712, O9713, O9714, O9715, O9716, O9717, O9718, O9719, O9720, O9721, O9722, O9723, O9724, O9725, O9726, O9727, O9728, O9729, O9730, O9731, O9732, O9733, O9734, O9735, O9736, O9737, O9738, O9739, O9740, O9741, O9742, O9743, O9744, O9745, O9746, O9747, O9748, O9749, O9750, O9751, O9752, O9753, O9754, O9755, O9756, O9757, O9758, O9759, O9760, O9761, O9762, O9763, O9764, O9765, O9766, O9767, O9768, O9769, O9770, O9771, O9772, O9773, O9774, O9775, O9776, O9777, O9778, O9779, O9780, O9781, O9782, O9783, O9784, O9785, O9786, O9787, O9788, O9789, O9790, O9791, O9792, O9793, O9794, O9795, O9796, O9797, O9798, O9799, O9800, O9801, O9802, O9803, O9804, O9805, O9806, O9807, O9808, O9809, O9810, O9811, O9812, O9813, O9814, O9815, O9816, O9817, O9818, O9819, O9820, O9821, O9822, O9823, O9824, O9825, O9826, O9827, O9828, O9829, O9830, O9831, O9832, O9833, O9834, O9835, O9836, O9837, O9838, O9839, O9840, O9841, O9842, O9843, O9844, O9845, O9846, O9847, O9848, O9849, O9850, O9851, O9852, O9853, O9854, O9855, O9856, O9857, O9858, O9859, O9860, O9861, O9862, O9863, O9864, O9865, O9866, O9867, O9868, O9869, O9870, O9871, O9872, O9873, O9874, O9875, O9876, O9877, O9878, O9879, O9880, O9881, O9882, O9883, O9884, O9885, O9886, O9887, O9888, O9889, O9890, O9891, O9892, O9893, O9894, O9895, O9896, O9897, O9898, O9899, O9900, O9901, O9902, O9903, O9904, O9905, O9906, O9907, O9908, O9909, O9910, O9911, O9912, O9913, O9914, O9915, O9916, O9917, O9918, O9919, O9920, O9921, O9922, O9923, O9924, O9925, O9926, O9927, O9928, O9929, O9930, O9931, O9932, O9933, O9934, O9935, O9936, O9937, O9938, O9939, O9940, O9941, O9942, O9943, O9944, O9945, O9946, O9947, O9948, O9949, O9950, O9951, O9952, O9953, O9954, O9955, O9956, O9957, O9958, O9959, O9960, O9961, O9962, O9963, O9964, O9965, O9966, O9967, O9968, O9969, O9970, O9971, O9972, O9973, O9974, O9975, O9976, O9977, O9978, O9979, O9980, O9981, O9982, O9983, O9984, O9985, O9986, O9987, O9988, O9989, O9990, O9991, O9992, O9993, O9994, O9995, O9996, O9997, O9998, O9999, O10000, O10001, O10002, O10003, O10004, O10005, O10006, O10007, O10008, O10009, O10010, O10011, O10012, O10013, O10014, O10015, O10016, O10017, O10018, O10019, O10020, O10021, O10022, O10023, O10024, O10025, O10026, O10027, O10028, O10029, O10030, O10031, O10032, O10033, O10034, O10035, O10036, O10037, O10038, O10039, O10040, O10041, O10042, O10043, O10044, O10045, O10046, O10047, O10048, O10049, O10050, O10051, O10052, O10053, O10054, O10055, O10056, O10057, O10058, O10059, O10060, O10061, O10062, O10063, O10064, O10065, O10066, O10067, O10068, O10069, O10070, O10071, O10072, O10073, O10074, O10075, O10076, O10077, O10078, O10079, O10080, O10081, O10082, O10083, O10084, O10085, O10086, O10087, O10088, O10089, O10090, O10091, O10092, O10093, O10094, O10095, O10096, O10097, O10098, O10099, O10100, O10101, O10102, O10103, O10104, O10105, O10106, O10107, O10108, O10109, O10110, O10111, O10112, O10113, O10114, O10115, O10116, O10117, O10118, O10119, O10120, O10121, O10122, O10123, O10124, O10125, O10126, O10127, O10128, O10129, O10130, O10131, O10132, O10133, O10134, O10135, O10136, O10137, O10138, O10139, O10140, O10141, O10142, O10143, O10144, O10145, O10146, O10147, O10148, O10149, O10150, O10151, O10152, O10153, O10154, O10155, O10156, O10157, O10158, O10159, O10160, O10161, O10162, O10163, O10164, O10165, O10166, O10167, O10168, O10169, O10170, O10171, O10172, O10173, O10174, O10175, O10176, O10177, O10178, O10179, O10180, O10181, O10182, O10183, O10184, O10185, O10186, O10187, O10188, O10189, O10190, O10191, O10192, O10193, O10194, O10195, O10196, O10197, O10198, O10199, O10200, O10201, O10202, O10203, O10204, O10205, O10206, O10207, O10208, O10209, O10210, O10211, O10212, O10213, O10214, O10215, O10216, O10217, O10218, O10219, O10220, O10221, O10222, O10223, O10224, O10225, O10226, O10227, O10228, O10229, O10230, O10231, O10232, O10233, O10234, O10235, O10236, O10237, O10238, O10239, O10240, O10241, O10242, O10243, O10244, O10245, O10246, O10247, O10248, O10249, O10250, O10251, O10252, O10253, O10254, O10255, O10256, O10257, O10258, O10259, O10260, O10261, O10262, O10263, O10264, O10265, O10266, O10267, O10268, O10269, O10270, O10271, O10272, O10273, O10274, O10275, O10276, O10277, O10278, O10279, O10280, O10281, O10282, O10283, O10284, O10285, O10286, O10287, O10288, O10289, O10290, O10291, O10292, O10293, O10294, O10295, O10296, O10297, O10298, O10299, O10300, O10301, O10302, O10303, O10304, O10305, O10306, O10307, O10308, O10309, O10310, O10311, O10312, O10313, O10314, O10315, O10316, O10317, O10318, O10319, O10320, O10321, O10322, O10323, O10324, O10325, O10326, O10327, O10328, O10329, O10330, O10331, O10332, O10333, O10334, O10335, O10336, O10337, O10338, O10339, O10340, O10341, O10342, O10343, O10344, O10345, O10346, O10347, O10348, O10349, O10350, O10351, O10352, O10353, O10354, O10355, O10356, O10357, O10358, O10359, O10360, O10361, O10362, O10363, O10364, O10365, O10366, O10367, O10368, O10369, O10370, O10371, O10372, O10373, O10374, O10375, O10376, O10377, O10378, O10379, O10380, O10381, O10382, O10383, O10384, O10385, O10386, O10387, O10388, O10389, O10390, O10391, O10392, O10393, O10394, O10395, O10396, O10397, O10398, O10399, O10400, O10401, O10402, O10403, O10404, O10405, O10406, O10407, O10408, O10409, O10410, O10411, O10412, O10413, O10414, O10415, O10416, O10417, O10418, O10419, O10420, O10421, O10422, O10423, O10424, O10425, O10426, O10427, O10428, O10429, O10430, O10431, O10432, O10433, O10434, O10435, O10436, O10437, O10438, O10439, O10440, O10441, O10442, O10443, O10444, O10445, O10446, O10447, O10448, O10449, O10450, O10451, O10452, O10453, O10454, O10455, O10456, O10457, O10458, O10459, O10460, O10461, O10462, O10463, O10464, O10465, O10466, O10467, O10468, O10469, O10470, O10471, O10472, O10473, O10474, O10475, O10476, O10477, O10478, O10479, O10480, O10481, O10482, O10483, O10484, O10485, O10486, O10487, O10488, O10489, O10490, O10491, O10492, O10493, O10494, O10495, O10496, O10497, O10498, O10499, O10500, O10501, O10502, O10503, O10504, O10505, O10506, O10507, O10508, O10509, O10510, O10511, O10512, O10513, O10514, O10515, O10516, O10517, O10518, O10519, O10520, O10521, O10522, O10523, O10524, O10525, O10526, O10527, O10528, O10529, O10530, O10531, O10532, O10533, O10534, O10535, O10536, O10537, O10538, O10539, O10540, O10541, O10542, O10543, O10544, O10545, O10546, O10547, O10548, O10549, O10550, O10551, O10552, O10553, O10554, O10555, O10556, O10557, O10558, O10559, O10560, O10561, O10562, O10563, O10564, O10565, O10566, O10567, O10568, O10569, O10570, O10571, O10572, O10573, O10574, O10575, O10576, O10577, O10578, O10579, O10580, O10581, O10582, O10583, O10584, O10585, O10586, O10587, O10588, O10589, O10590, O10591, O10592, O10593, O10594, O10595, O10596, O10597, O10598, O10599, O10600, O10601, O10602, O10603, O10604, O10605, O10606, O10607, O10608, O10609, O10610, O10611, O10612, O10613, O10614, O10615, O10616, O10617, O10618, O10619, O10620, O10621, O10622, O10623, O10624, O10625, O10626, O10627, O10628, O10629, O10630, O10631, O10632, O10633, O10634, O10635, O10636, O10637, O10638, O10639, O10640, O10641, O10642, O10643, O10644, O10645, O10646, O10647, O10648, O10649, O10650, O10651, O10652, O10653, O10654, O10655, O10656, O10657, O10658, O10659, O10660, O10661, O10662, O10663, O10664, O10665, O10666, O10667, O10668, O10669, O10670, O10671, O10672, O10673, O10674, O10675, O10676, O10677, O10678, O10679, O10680, O10681, O10682, O10683, O10684, O10685, O10686, O10687, O10688, O10689, O10690, O10691, O10692, O10693, O10694, O10695, O10696, O10697, O10698, O10699, O10700, O10701, O10702, O10703, O10704, O10705, O10706, O10707, O10708, O10709, O10710, O10711, O10712, O10713, O10714, O10715, O10716, O10717, O10718, O10719, O10720, O10721, O10722, O10723, O10724, O10725, O10726, O10727, O10728, O10729, O10730, O10731, O10732, O10733, O10734, O10735, O10736, O10737, O10738, O10739, O10740, O10741, O10742, O10743, O10744, O10745, O10746, O10747, O10748, O10749, O10750, O10751, O10752, O10753, O10754, O10755, O10756, O10757, O10758, O10759, O10760, O10761, O10762, O10763, O10764, O10765, O10766, O10767, O10768, O10769, O10770, O10771, O10772, O10773, O10774, O10775, O10776, O10777, O10778, O10779, O10780, O10781, O10782, O10783, O10784, O10785, O10786, O10787, O10788, O10789, O10790, O10791, O10792, O10793, O10794, O10795, O10796, O10797, O10798, O10799, O10800, O10801, O10802, O10803, O10804, O10805, O10806, O10807, O10808, O10809, O10810, O10811, O10812, O10813, O10814, O10815, O10816, O10817, O10818, O10819, O10820, O10821, O10822, O10823, O10824, O10825, O10826, O10827, O10828, O10829, O10830, O10831, O10832, O10833, O10834, O10835, O10836, O10837, O10838, O10839, O10840, O10841, O10842, O10843, O10844, O10845, O10846, O10847, O10848, O10849, O10850, O10851, O10852, O10853, O10854, O10855, O10856, O10857, O10858, O10859, O10860, O10861, O10862, O10863, O10864, O10865, O10866, O10867, O10868, O10869, O10870, O10871, O10872, O10873, O10874, O10875, O10876, O10877, O10878, O10879, O10880, O10881, O10882, O10883, O10884, O10885, O10886, O10887, O10888, O10889, O10890, O10891, O10892, O10893, O10894, O10895, O10896, O10897, O10898, O10899, O10900, O10901, O10902, O10903, O10904, O10905, O10906, O10907, O10908, O10909, O10910, O10911, O10912, O10913, O10914, O10915, O10916, O10917, O10918, O10919, O10920, O10921, O10922, O10923, O10924, O10925, O10926, O10927, O10928, O10929, O10930, O10931, O10932, O10933, O10934, O10935, O10936, O10937, O10938, O10939, O10940, O10941, O10942, O10943, O10944, O10945, O10946, O10947, O10948, O10949, O10950, O10951, O10952, O10953, O10954, O10955, O10956, O10957, O10958, O10959, O10960, O10961, O10962, O10963, O10964, O10965, O10966, O10967, O10968, O10969, O10970, O10971, O10972, O10973, O10974, O10975, O10976, O10977, O10978, O10979, O10980, O10981, O10982, O10983, O10984, O10985, O10986, O10987, O10988, O10989, O10990, O10991, O10992, O10993, O10994, O10995, O10996, O10997, O10998, O10999, O11000, O11001, O11002, O11003, O11004, O11005, O11006, O11007, O11008, O11009, O11010, O11011, O11012, O11013, O11014, O11015, O11016, O11017, O11018, O11019, O11020, O11021, O11022, O11023, O11024, O11025, O11026, O11027, O11028, O11029, O11030, O11031, O11032, O11033, O11034, O11035, O11036, O11037, O11038, O11039, O11040, O11041, O11042, O11043, O11044, O11045, O11046, O11047, O11048, O11049, O11050, O11051, O11052, O11053, O11054, O11055, O11056, O11057, O11058, O11059, O11060, O11061, O11062, O11063, O11064, O11065, O11066, O11067, O11068, O11069, O11070, O11071, O11072, O11073, O11074, O11075, O11076, O11077, O11078, O11079, O11080, O11081, O11082, O11083, O11084, O11085, O11086, O11087, O11088, O11089, O11090, O11091, O11092, O11093, O11094, O11095, O11096, O11097, O11098, O11099, O11100, O11101, O11102, O11103, O11104, O11105, O11106, O11107, O11108, O11109, O11110, O11111, O11112, O11113, O11114, O11115, O11116, O11117, O11118, O11119, O11120, O11121, O11122, O11123, O11124, O11125, O11126, O11127, O11128, O11129, O11130, O11131, O11132, O11133, O11134, O11135, O11136, O11137, O11138, O11139, O11140, O11141, O11142, O11143, O11144, O11145, O11146, O11147, O11148, O11149, O11150, O11151, O11152, O11153, O11154, O11155, O11156, O11157, O11158, O11159, O11160, O11161, O11162, O11163, O11164, O11165, O11166, O11167, O11168, O11169, O11170, O11171, O11172, O11173, O11174, O11175, O11176, O11177, O11178, O11179, O11180, O11181, O11182, O11183, O11184, O11185, O11186, O11187, O11188, O11189, O11190, O11191, O11192, O11193, O11194, O11195, O11196, O11197, O11198, O11199, O11200, O11201, O11202, O11203, O11204, O11205, O11206, O11207, O11208, O11209, O11210, O11211, O11212, O11213, O11214, O11215, O11216, O11217, O11218, O11219, O11220, O11221, O11222, O11223, O11224, O11225, O11226, O11227, O11228, O11229, O11230, O11231, O11232, O11233, O11234, O11235, O11236, O11237, O11238, O11239, O11240, O11241, O11242, O11243, O11244, O11245, O11246, O11247, O11248, O11249, O11250, O11251, O11252, O11253, O11254, O11255, O11256, O11257, O11258, O11259, O11260, O11261, O11262, O11263, O11264, O11265, O11266, O11267, O11268, O11269, O11270, O11271, O11272, O11273, O11274, O11275, O11276, O11277, O11278, O11279, O11280, O11281, O11282, O11283, O11284, O11285, O11286, O11287, O11288, O11289, O11290, O11291, O11292, O11293, O11294, O11295, O11296, O11297, O11298, O11299, O11300, O11301, O11302, O11303, O11304, O11305, O11306, O11307, O11308, O11309, O11310, O11311, O11312, O11313, O11314, O11315, O11316, O11317, O11318, O11319, O11320, O11321, O11322, O11323, O11324, O11325, O11326, O11327, O11328, O11329, O11330, O11331, O11332, O11333, O11334, O11335, O11336, O11337, O11338, O11339, O11340, O11341, O11342, O11343, O11344, O11345, O11346, O11347, O11348, O11349, O11350, O11351, O11352, O11353, O11354, O11355, O11356, O11357, O11358, O11359, O11360, O11361, O11362, O11363, O11364, O11365, O11366, O11367, O11368, O11369, O11370, O11371, O11372, O11373, O11374, O11375, O11376, O11377, O11378, O11379, O11380, O11381, O11382, O11383, O11384, O11385, O11386, O11387, O11388, O11389, O11390, O11391, O11392, O11393, O11394, O11395, O11396, O11397, O11398, O11399, O11400, O11401, O11402, O11403, O11404, O11405, O11406, O11407, O11408, O11409, O11410, O11411, O11412, O11413, O11414, O11415, O11416, O11417, O11418, O11419, O11420, O11421, O11422, O11423, O11424, O11425, O11426, O11427, O11428, O11429, O11430, O11431, O11432, O11433, O11434, O11435, O11436, O11437, O11438, O11439, O11440, O11441, O11442, O11443, O11444, O11445, O11446, O11447, O11448, O11449, O11450, O11451, O11452, O11453, O11454, O11455, O11456, O11457, O11458, O11459, O11460, O11461, O11462, O11463, O11464, O11465, O11466, O11467, O11468, O11469, O11470, O11471, O11472, O11473, O11474, O11475, O11476, O11477, O11478, O11479, O11480, O11481, O11482, O11483, O11484, O11485, O11486, O11487, O11488, O11489, O11490, O11491, O11492, O11493, O11494, O11495, O11496, O11497, O11498, O11499, O11500, O11501, O11502, O11503, O11504, O11505, O11506, O11507, O11508, O11509, O11510, O11511, O11512, O11513, O11514, O11515, O11516, O11517, O11518, O11519, O11520, O11521, O11522, O11523, O11524, O11525, O11526, O11527, O11528, O11529, O11530, O11531, O11532, O11533, O11534, O11535, O11536, O11537, O11538, O11539, O11540, O11541, O11542, O11543, O11544, O11545, O11546, O11547, O11548, O11549, O11550, O11551, O11552, O11553, O11554, O11555, O11556, O11557, O11558, O11559, O11560, O11561, O11562, O11563, O11564, O11565, O11566, O11567, O11568, O11569, O11570, O11571, O11572, O11573, O11574, O11575, O11576, O11577, O11578, O11579, O11580, O11581, O11582, O11583, O11584, O11585, O11586, O11587, O11588, O11589, O11590, O11591, O11592, O11593, O11594, O11595, O11596, O11597, O11598, O11599, O11600, O11601, O11602, O11603, O11604, O11605, O11606, O11607, O11608, O11609, O11610, O11611, O11612, O11613, O11614, O11615, O11616, O11617, O11618, O11619, O11620, O11621, O11622, O11623, O11624, O11625, O11626, O11627, O11628, O11629, O11630, O11631, O11632, O11633, O11634, O11635, O11636, O11637, O11638, O11639, O11640, O11641, O11642, O11643, O11644, O11645, O11646, O11647, O11648, O11649, O11650, O11651, O11652, O11653, O11654, O11655, O11656, O11657, O11658, O11659, O11660, O11661, O11662, O11663, O11664, O11665, O11666, O11667, O11668, O11669, O11670, O11671, O11672, O11673, O11674, O11675, O11676, O11677, O11678, O11679, O11680, O11681, O11682, O11683, O11684, O11685, O11686, O11687, O11688, O11689, O11690, O11691, O11692, O11693, O11694, O11695, O11696, O11697, O11698, O11699, O11700, O11701, O11702, O11703, O11704, O11705, O11706, O11707, O11708, O11709, O11710, O11711, O11712, O11713, O11714, O11715, O11716, O11717, O11718, O11719, O11720, O11721, O11722, O11723, O11724, O11725, O11726, O11727, O11728, O11729, O11730, O11731, O11732, O11733, O11734, O11735, O11736, O11737, O11738, O11739, O11740, O11741, O11742, O11743, O11744, O11745, O11746, O11747, O11748, O11749, O11750, O11751, O11752, O11753, O11754, O11755, O11756, O11757, O11758, O11759, O11760, O11761, O11762, O11763, O11764, O11765, O11766, O11767, O11768, O11769, O11770, O11771, O11772, O11773, O11774, O11775, O11776, O11777, O11778, O11779, O11780, O11781, O11782, O11783, O11784, O11785, O11786, O11787, O11788, O11789, O11790, O11791, O11792, O11793, O11794, O11795, O11796, O11797, O11798, O11799, O11800, O11801, O11802, O11803, O11804, O11805, O11806, O11807, O11808, O11809, O11810, O11811, O11812, O11813, O11814, O11815, O11816, O11817, O11818, O11819, O11820, O11821, O11822, O11823, O11824, O11825, O11826, O11827, O11828, O11829, O11830, O11831, O11832, O11833, O11834, O11835, O11836, O11837, O11838, O11839, O11840, O11841, O11842, O11843, O11844, O11845, O11846, O11847, O11848, O11849, O11850, O11851, O11852, O11853, O11854, O11855, O11856, O11857, O11858, O11859, O11860, O11861, O11862, O11863, O11864, O11865, O11866, O11867, O11868, O11869, O11870, O11871, O11872, O11873, O11874, O11875, O11876, O11877, O11878, O11879, O11880, O11881, O11882, O11883, O11884, O11885, O11886, O11887, O11888, O11889, O11890, O11891, O11892, O11893, O11894, O11895, O11896, O11897, O11898, O11899, O11900, O11901, O11902, O11903, O11904, O11905, O11906, O11907, O11908, O11909, O11910, O11911, O11912, O11913, O11914, O11915, O11916, O11917, O11918, O11919, O11920, O11921, O11922, O11923, O11924, O11925, O11926, O11927, O11928, O11929, O11930, O11931, O11932, O11933, O11934, O11935, O11936, O11937, O11938, O11939, O11940, O11941, O11942, O11943, O11944, O11945, O11946, O11947, O11948, O11949, O11950, O11951, O11952, O11953, O11954, O11955, O11956, O11957, O11958, O11959, O11960, O11961, O11962, O11963, O11964, O11965, O11966, O11967, O11968, O11969, O11970, O11971, O11972, O11973, O11974, O11975, O11976, O11977, O11978, O11979, O11980, O11981, O11982, O11983, O11984, O11985, O11986, O11987, O11988, O11989, O11990, O11991, O11992, O11993, O11994, O11995, O11996, O11997, O11998, O11999, O12000, O12001, O12002, O12003, O12004, O12005, O12006, O12007, O12008, O12009, O12010, O12011, O12012, O12013, O12014, O12015, O12016, O12017, O12018, O12019, O12020, O12021, O12022, O12023, O12024, O12025, O12026, O12027, O12028, O12029, O12030, O12031, O12032, O12033, O12034, O12035, O12036, O12037, O12038, O12039, O12040, O12041, O12042, O12043, O12044, O12045, O12046, O12047, O12048, O12049, O12050, O12051, O12052, O12053, O12054, O12055, O12056, O12057, O12058, O12059, O12060, O12061, O12062, O12063, O12064, O12065, O12066, O12067, O12068, O12069, O12070, O12071, O12072, O12073, O12074, O12075, O12076, O12077, O12078, O12079, O12080, O12081, O12082, O12083, O12084, O12085, O12086, O12087, O12088, O12089, O12090, O12091, O12092, O12093, O12094, O12095, O12096, O12097, O12098, O12099, O12100, O12101, O12102, O12103, O12104, O12105, O12106, O12107, O12108, O12109, O12110, O12111, O12112, O12113, O12114, O12115, O12116, O12117, O12118, O12119, O12120, O12121, O12122, O12123, O12124, O12125, O12126, O12127, O12128, O12129, O12130, O12131, O12132, O12133, O12134, O12135, O12136, O12137, O12138, O12139, O12140, O12141, O12142, O12143, O12144, O12145, O12146, O12147, O12148, O12149, O12150, O12151, O12152, O12153, O12154, O12155, O12156, O12157, O12158, O12159, O12160, O12161, O12162, O12163, O12164, O12165, O12166, O12167, O12168, O12169, O12170, O12171, O12172, O12173, O12174, O12175, O12176, O12177, O12178, O12179, O12180, O12181, O12182, O12183, O12184, O12185, O12186, O12187, O12188, O12189, O12190, O12191, O12192, O12193, O12194, O12195, O12196, O12197, O12198, O12199, O12200, O12201, O12202, O12203, O12204, O12205, O12206, O12207, O12208, O12209, O12210, O12211, O12212, O12213, O12214, O12215, O12216, O12217, O12218, O12219, O12220, O12221, O12222, O12223, O12224, O12225, O12226, O12227, O12228, O12229, O12230, O12231, O12232, O12233, O12234, O12235, O12236, O12237, O12238, O12239, O12240, O12241, O12242, O12243, O12244, O12245, O12246, O12247, O12248, O12249, O12250, O12251, O12252, O12253, O12254, O12255, O12256, O12257, O12258, O12259, O12260, O12261, O12262, O12263, O12264, O12265, O12266, O12267, O12268, O12269, O12270, O12271, O12272, O12273, O12274, O12275, O12276, O12277, O12278, O12279, O12280, O12281, O12282, O12283, O12284, O12285, O12286, O12287, O12288, O12289, O12290, O12291, O12292, O12293, O12294, O12295, O12296, O12297, O12298, O12299, O12300, O12301, O12302, O12303, O12304, O12305, O12306, O12307, O12308, O12309, O12310, O12311, O12312, O12313, O12314, O12315, O12316, O12317, O12318, O12319, O12320, O12321, O12322, O12323, O12324, O12325, O12326, O12327, O12328, O12329, O12330, O12331, O12332, O12333, O12334, O12335, O12336, O12337, O12338, O12339, O12340, O12341, O12342, O12343, O12344, O12345, O12346, O12347, O12348, O12349, O12350, O12351, O12352, O12353, O12354, O12355, O12356, O12357, O12358, O12359, O12360, O12361, O12362, O12363, O12364, O12365, O12366, O12367, O12368, O12369, O12370, O12371, O12372, O12373, O12374, O12375, O12376, O12377, O12378, O12379, O12380, O12381, O12382, O12383, O12384, O12385, O12386, O12387, O12388, O12389, O12390, O12391, O12392, O12393, O12394, O12395, O12396, O12397, O12398, O12399, O12400, O12401, O12402, O12403, O12404, O12405, O12406, O12407, O12408, O12409, O12410, O12411, O12412, O12413, O12414, O12415, O12416, O12417, O12418, O12419, O12420, O12421, O12422, O12423, O12424, O12425, O12426, O12427, O12428, O12429, O12430, O12431, O12432, O12433, O12434, O12435, O12436, O12437, O12438, O12439, O12440, O12441, O12442, O12443, O12444, O12445, O12446, O12447, O12448, O12449, O12450, O12451, O12452, O12453, O12454, O12455, O12456, O12457, O12458, O12459, O12460, O12461, O12462, O12463, O12464, O12465, O12466, O12467, O12468, O12469, O12470, O12471, O12472, O12473, O12474, O12475, O12476, O12477, O12478, O12479, O12480, O12481, O12482, O12483, O12484, O12485, O12486, O12487, O12488, O12489, O12490, O12491, O12492, O12493, O12494, O12495, O12496, O12497, O12498, O12499, O12500, O12501, O12502, O12503, O12504, O12505, O12506, O12507, O12508, O12509, O12510, O12511, O12512, O12513, O12514, O12515, O12516, O12517, O12518, O12519, O12520, O12521, O12522, O12523, O12524, O12525, O12526, O12527, O12528, O12529, O12530, O12531, O12532, O12533, O12534, O12535, O12536, O12537, O12538, O12539, O12540, O12541, O12542, O12543, O12544, O12545, O12546, O12547, O12548, O12549, O12550, O12551, O12552, O12553, O12554, O12555, O12556, O12557, O12558, O12559, O12560, O12561, O12562, O12563, O12564, O12565, O12566, O12567, O12568, O12569, O12570, O12571, O12572, O12573, O12574, O12575, O12576, O12577, O12578, O12579, O12580, O12581, O12582, O12583, O12584, O12585, O12586, O12587, O12588, O12589, O12590, O12591, O12592, O12593, O12594, O12595, O12596, O12597, O12598, O12599, O12600, O12601, O12602, O12603, O12604, O12605, O12606, O12607, O12608, O12609, O12610, O12611, O12612, O12613, O12614, O12615, O12616, O12617, O12618, O12619, O12620, O12621, O12622, O12623, O12624, O12625, O12626, O12627, O12628, O12629, O12630, O12631, O12632, O12633, O12634, O12635, O12636, O12637, O12638, O12639, O12640, O12641, O12642, O12643, O12644, O12645, O12646, O12647, O12648, O12649, O12650, O12651, O12652, O12653, O12654, O12655, O12656, O12657, O12658, O12659, O12660, O12661, O12662, O12663, O12664, O12665, O12666, O12667, O12668, O12669, O12670, O12671, O12672, O12673, O12674, O12675, O12676, O12677, O12678, O12679, O12680, O12681, O12682, O12683, O12684, O12685, O12686, O12687, O12688, O12689, O12690, O12691, O12692, O12693, O12694, O12695, O12696, O12697, O12698, O12699, O12700, O12701, O12702, O12703, O12704, O12705, O12706, O12707, O12708, O12709, O12710, O12711, O12712, O12713, O12714, O12715, O12716, O12717, O12718, O12719, O12720, O12721, O12722, O12723, O12724, O12725, O12726, O12727, O12728, O12729, O12730, O12731, O12732, O12733, O12734, O12735, O12736, O12737, O12738, O12739, O12740, O12741, O12742, O12743, O12744, O12745, O12746, O12747, O12748, O12749, O12750, O12751, O12752, O12753, O12754, O12755, O12756, O12757, O12758, O12759, O12760, O12761, O12762, O12763, O12764, O12765, O12766, O12767, O12768, O12769, O12770, O12771, O12772, O12773, O12774, O12775, O12776, O12777, O12778, O12779, O12780, O12781, O12782, O12783, O12784, O12785, O12786, O12787, O12788, O12789, O12790, O12791, O12792, O12793, O12794, O12795, O12796, O12797, O12798, O12799, O12800, O12801, O12802, O12803, O12804, O12805, O12806, O12807, O12808, O12809, O12810, O12811, O12812, O12813, O12814, O12815, O12816, O12817, O12818, O12819, O12820, O12821, O12822, O12823, O12824, O12825, O12826, O12827, O12828, O12829, O12830, O12831, O12832, O12833, O12834, O12835, O12836, O12837, O12838, O12839, O12840, O12841, O12842, O12843, O12844, O12845, O12846, O12847, O12848, O12849, O12850, O12851, O12852, O12853, O12854, O12855, O12856, O12857, O12858, O12859, O12860, O12861, O12862, O12863, O12864, O12865, O12866, O12867, O12868, O12869, O12870, O12871, O12872, O12873, O12874, O12875, O12876, O12877, O12878, O12879, O12880, O12881, O12882, O12883, O12884, O12885, O12886, O12887, O12888, O12889, O12890, O12891, O12892, O12893, O12894, O12895, O12896, O12897, O12898, O12899, O12900, O12901, O12902, O12903, O12904, O12905, O12906, O12907, O12908, O12909, O12910, O12911, O12912, O12913, O12914, O12915, O12916, O12917, O12918, O12919, O12920, O12921, O12922, O12923, O12924, O12925, O12926, O12927, O12928, O12929, O12930, O12931, O12932, O12933, O12934, O12935, O12936, O12937, O12938, O12939, O12940, O12941, O12942, O12943, O12944, O12945, O12946, O12947, O12948, O12949, O12950, O12951, O12952, O12953, O12954, O12955, O12956, O12957, O12958, O12959, O12960, O12961, O12962, O12963, O12964, O12965, O12966, O12967, O12968, O12969, O12970, O12971, O12972, O12973, O12974, O12975, O12976, O12977, O12978, O12979, O12980, O12981, O12982, O12983, O12984, O12985, O12986, O12987, O12988, O12989, O12990, O12991, O12992, O12993, O12994, O12995, O12996, O12997, O12998, O12999, O13000, O13001, O13002, O13003, O13004, O13005, O13006, O13007, O13008, O13009, O13010, O13011, O13012, O13013, O13014, O13015, O13016, O13017, O13018, O13019, O13020, O13021, O13022, O13023, O13024, O13025, O13026, O13027, O13028, O13029, O13030, O13031, O13032, O13033, O13034, O13035, O13036, O13037, O13038, O13039, O13040, O13041, O13042, O13043, O13044, O13045, O13046, O13047, O13048, O13049, O13050, O13051, O13052, O13053, O13054, O13055, O13056, O13057, O13058, O13059, O13060, O13061, O13062, O13063, O13064, O13065, O13066, O13067, O13068, O13069, O13070, O13071, O13072, O13073, O13074, O13075, O13076, O13077, O13078, O13079, O13080, O13081, O13082, O13083, O13084, O13085, O13086, O13087, O13088, O13089, O13090, O13091, O13092, O13093, O13094, O13095, O13096, O13097, O13098, O13099, O13100, O13101, O13102, O13103, O13104, O13105, O13106, O13107, O13108, O13109, O13110, O13111, O13112, O13113, O13114, O13115, O13116, O13117, O13118, O13119, O13120, O13121, O13122, O13123, O13124, O13125, O13126, O13127, O13128, O13129, O13130, O13131, O13132, O13133, O13134, O13135, O13136, O13137, O13138, O13139, O13140, O13141, O13142, O13143, O13144, O13145, O13146, O13147, O13148, O13149, O13150, O13151, O13152, O13153, O13154, O13155, O13156, O13157, O13158, O13159, O13160, O13161, O13162, O13163, O13164, O13165, O13166, O13167, O13168, O13169, O13170, O13171, O13172, O13173, O13174, O13175, O13176, O13177, O13178, O13179, O13180, O13181, O13182, O13183, O13184, O13185, O13186, O13187, O13188, O13189, O13190, O13191, O13192, O13193, O13194, O13195, O13196, O13197, O13198, O13199, O13200, O13201, O13202, O13203, O13204, O13205, O13206, O13207, O13208, O13209, O13210, O13211, O13212, O13213, O13214, O13215, O13216, O13217, O13218, O13219, O13220, O13221, O13222, O13223, O13224, O13225, O13226, O13227, O13228, O13229, O13230, O13231, O13232, O13233, O13234, O13235, O13236, O13237, O13238, O13239, O13240, O13241, O13242, O13243, O13244, O13245, O13246, O13247, O13248, O13249, O13250, O13251, O13252, O13253, O13254, O13255, O13256, O13257, O13258, O13259, O13260, O13261, O13262, O13263, O13264, O13265, O13266, O13267, O13268, O13269, O13270, O13271, O13272, O13273, O13274, O13275, O13276, O13277, O13278, O13279, O13280, O13281, O13282, O13283, O13284, O13285, O13286, O13287, O13288, O13289, O13290, O13291, O13292, O13293, O13294, O13295, O13296, O13297, O13298, O13299, O13300, O13301, O13302, O13303, O13304, O13305, O13306, O13307, O13308, O13309, O13310, O13311, O13312, O13313, O13314, O13315, O13316, O13317, O13318, O13319, O13320, O13321, O13322, O13323, O13324, O13325, O13326, O13327, O13328, O13329, O13330, O13331, O13332, O13333, O13334, O13335, O13336, O13337, O13338, O13339, O13340, O13341, O13342, O13343, O13344, O13345, O13346, O13347, O13348, O13349, O13350, O13351, O13352, O13353, O13354, O13355, O13356, O13357, O13358, O13359, O13360, O13361, O13362, O13363, O13364, O13365, O13366, O13367, O13368, O13369, O13370, O13371, O13372, O13373, O13374, O13375, O13376, O13377, O13378, O13379, O13380, O13381, O13382, O13383, O13384, O13385, O13386, O13387, O13388, O13389, O13390, O13391, O13392, O13393, O13394, O13395, O13396, O13397, O13398, O13399, O13400, O13401, O13402, O13403, O13404, O13405, O13406, O13407, O13408, O13409, O13410, O13411, O13412, O13413, O13414, O13415, O13416, O13417, O13418, O13419, O13420, O13421, O13422, O13423, O13424, O13425, O13426, O13427, O13428, O13429, O13430, O13431, O13432, O13433, O13434, O13435, O13436, O13437, O13438, O13439, O13440, O13441, O13442, O13443, O13444, O13445, O13446, O13447, O13448, O13449, O13450, O13451, O13452, O13453, O13454, O13455, O13456, O13457, O13458, O13459, O13460, O13461, O13462, O13463, O13464, O13465, O13466, O13467, O13468, O13469, O13470, O13471, O13472, O13473, O13474, O13475, O13476, O13477, O13478, O13479, O13480, O13481, O13482, O13483, O13484, O13485, O13486, O13487, O13488, O13489, O13490, O13491, O13492, O13493, O13494, O13495, O13496, O13497, O13498, O13499, O13500, O13501, O13502, O13503, O13504, O13505, O13506, O13507, O13508, O13509, O13510, O13511, O13512, O13513, O13514, O13515, O13516, O13517, O13518, O13519, O13520, O13521, O13522, O13523, O13524, O13525, O13526, O13527, O13528, O13529, O13530, O13531, O13532, O13533, O13534, O13535, O13536, O13537, O13538, O13539, O13540, O13541, O13542, O13543, O13544, O13545, O13546, O13547, O13548, O13549, O13550, O13551, O13552, O13553, O13554, O13555, O13556, O13557, O13558, O13559, O13560, O13561, O13562, O13563, O13564, O13565, O13566, O13567, O13568, O13569, O13570, O13571, O13572, O13573, O13574, O13575, O13576, O13577, O13578, O13579, O13580, O13581, O13582, O13583, O13584, O13585, O13586, O13587, O13588, O13589, O13590, O13591, O13592, O13593, O13594, O13595, O13596, O13597, O13598, O13599, O13600, O13601, O13602, O13603, O13604, O13605, O13606, O13607, O13608, O13609, O13610, O13611, O13612, O13613, O13614, O13615, O13616, O13617, O13618, O13619, O13620, O13621, O13622, O13623, O13624, O13625, O13626, O13627, O13628, O13629, O13630, O13631, O13632, O13633, O13634, O13635, O13636, O13637, O13638, O13639, O13640, O13641, O13642, O13643, O13644, O13645, O13646, O13647, O13648, O13649, O13650, O13651, O13652, O13653, O13654, O13655, O13656, O13657, O13658, O13659, O13660, O13661, O13662, O13663, O13664, O13665, O13666, O13667, O13668, O13669, O13670, O13671, O13672, O13673, O13674, O13675, O13676, O13677, O13678, O13679, O13680, O13681, O13682, O13683, O13684, O13685, O13686, O13687, O13688, O13689, O13690, O13691, O13692, O13693, O13694, O13695, O13696, O13697, O13698, O13699, O13700, O13701, O13702, O13703, O13704, O13705, O13706, O13707, O13708, O13709, O13710, O13711, O13712, O13713, O13714, O13715, O13716, O13717, O13718, O13719, O13720, O13721, O13722, O13723, O13724, O13725, O13726, O13727, O13728, O13729, O13730, O13731, O13732, O13733, O13734, O13735, O13736, O13737, O13738, O13739, O13740, O13741, O13742, O13743, O13744, O13745, O13746, O13747, O13748, O13749, O13750, O13751, O13752, O13753, O13754, O13755, O13756, O13757, O13758, O13759, O13760, O13761, O13762, O13763, O13764, O13765, O13766, O13767, O13768, O13769, O13770, O13771, O13772, O13773, O13774, O13775, O13776, O13777, O13778, O13779, O13780, O13781, O13782, O13783, O13784, O13785, O13786, O13787, O13788, O13789, O13790, O13791, O13792, O13793, O13794, O13795, O13796, O13797, O13798, O13799, O13800, O13801, O13802, O13803, O13804, O13805, O13806, O13807, O13808, O13809, O13810, O13811, O13812, O13813, O13814, O13815, O13816, O13817, O13818, O13819, O13820, O13821, O13822, O13823, O13824, O13825, O13826, O13827, O13828, O13829, O13830, O13831, O13832, O13833, O13834, O13835, O13836, O13837, O13838, O13839, O13840, O13841, O13842, O13843, O13844, O13845, O13846, O13847, O13848, O13849, O13850, O13851, O13852, O13853, O13854, O13855, O13856, O13857, O13858, O13859, O13860, O13861, O13862, O13863, O13864, O13865, O13866, O13867, O13868, O13869, O13870, O13871, O13872, O13873, O13874, O13875, O13876, O13877, O13878, O13879, O13880, O13881, O13882, O13883, O13884, O13885, O13886, O13887, O13888, O13889, O13890, O13891, O13892, O13893, O13894, O13895, O13896, O13897, O13898, O13899, O13900, O13901, O13902, O13903, O13904, O13905, O13906, O13907, O13908, O13909, O13910, O13911, O13912, O13913, O13914, O13915, O13916, O13917, O13918, O13919, O13920, O13921, O13922, O13923, O13924, O13925, O13926, O13927, O13928, O13929, O13930, O13931, O13932, O13933, O13934, O13935, O13936, O13937, O13938, O13939, O13940, O13941, O13942, O13943, O13944, O13945, O13946, O13947, O13948, O13949, O13950, O13951, O13952, O13953, O13954, O13955, O13956, O13957, O13958, O13959, O13960, O13961, O13962, O13963, O13964, O13965, O13966, O13967, O13968, O13969, O13970, O13971, O13972, O13973, O13974, O13975, O13976, O13977, O13978, O13979, O13980, O13981, O13982, O13983, O13984, O13985, O13986, O13987, O13988, O13989, O13990, O13991, O13992, O13993, O13994, O13995, O13996, O13997, O13998, O13999, O14000, O14001, O14002, O14003, O14004, O14005, O14006, O14007, O14008, O14009, O14010, O14011, O14012, O14013, O14014, O14015, O14016, O14017, O14018, O14019, O14020, O14021, O14022, O14023, O14024, O14025, O14026, O14027, O14028, O14029, O14030, O14031, O14032, O14033, O14034, O14035, O14036, O14037, O14038, O14039, O14040, O14041, O14042, O14043, O14044, O14045, O14046, O14047, O14048, O14049, O14050, O14051, O14052, O14053, O14054, O14055, O14056, O14057, O14058, O14059, O14060, O14061, O14062, O14063, O14064, O14065, O14066, O14067, O14068, O14069, O14070, O14071, O14072, O14073, O14074, O14075, O14076, O14077, O14078, O14079, O14080, O14081, O14082, O14083, O14084, O14085, O14086, O14087, O14088, O14089, O14090, O14091, O14092, O14093, O14094, O14095, O14096, O14097, O14098, O14099, O14100, O14101, O14102, O14103, O14104, O14105, O14106, O14107, O14108, O14109, O14110, O14111, O14112, O14113, O14114, O14115, O14116, O14117, O14118, O14119, O14120, O14121, O14122, O14123, O14124, O14125, O14126, O14127, O14128, O14129, O14130, O14131, O14132, O14133, O14134, O14135, O14136, O14137, O14138, O14139, O14140, O14141, O14142, O14143, O14144, O14145, O14146, O14147, O14148, O14149, O14150, O14151, O14152, O14153, O14154, O14155, O14156, O14157, O14158, O14159, O14160, O14161, O14162, O14163, O14164, O14165, O14166, O14167, O14168, O14169, O14170, O14171, O14172, O14173, O14174, O14175, O14176, O14177, O14178, O14179, O14180, O14181, O14182, O14183, O14184, O14185, O14186, O14187, O14188, O14189, O14190, O14191, O14192, O14193, O14194, O14195, O14196, O14197, O14198, O14199, O14200, O14201, O14202, O14203, O14204, O14205, O14206, O14207, O14208, O14209, O14210, O14211, O14212, O14213, O14214, O14215, O14216, O14217, O14218, O14219, O14220, O14221, O14222, O14223, O14224, O14225, O14226, O14227, O14228, O14229, O14230, O14231, O14232, O14233, O14234, O14235, O14236, O14237, O14238, O14239, O14240, O14241, O14242, O14243, O14244, O14245, O14246, O14247, O14248, O14249, O14250, O14251, O14252, O14253, O14254, O14255, O14256, O14257, O14258, O14259, O14260, O14261, O14262, O14263, O14264, O14265, O14266, O14267, O14268, O14269, O14270, O14271, O14272, O14273, O14274, O14275, O14276, O14277, O14278, O14279, O14280, O14281, O14282, O14283, O14284, O14285, O14286, O14287, O14288, O14289, O14290, O14291, O14292, O14293, O14294, O14295, O14296, O14297, O14298, O14299, O14300, O14301, O14302, O14303, O14304, O14305, O14306, O14307, O14308, O14309, O14310, O14311, O14312, O14313, O14314, O14315, O14316, O14317, O14318, O14319, O14320, O14321, O14322, O14323, O14324, O14325, O14326, O14327, O14328, O14329, O14330, O14331, O14332, O14333, O14334, O14335, O14336, O14337, O14338, O14339, O14340, O14341, O14342, O14343, O14344, O14345, O14346, O14347, O14348, O14349, O14350, O14351, O14352, O14353, O14354, O14355, O14356, O14357, O14358, O14359, O14360, O14361, O14362, O14363, O14364, O14365, O14366, O14367, O14368, O14369, O14370, O14371, O14372, O14373, O14374, O14375, O14376, O14377, O14378, O14379, O14380, O14381, O14382, O14383, O14384, O14385, O14386, O14387, O14388, O14389, O14390, O14391, O14392, O14393, O14394, O14395, O14396, O14397, O14398, O14399, O14400, O14401, O14402, O14403, O14404, O14405, O14406, O14407, O14408, O14409, O14410, O14411, O14412, O14413, O14414, O14415, O14416, O14417, O14418, O14419, O14420, O14421, O14422, O14423, O14424, O14425, O14426, O14427, O14428, O14429, O14430, O14431, O14432, O14433, O14434, O14435, O14436, O14437, O14438, O14439, O14440, O14441, O14442, O14443, O14444, O14445, O14446, O14447, O14448, O14449, O14450, O14451, O14452, O14453, O14454, O14455, O14456, O14457, O14458, O14459, O14460, O14461, O14462, O14463, O14464, O14465, O14466, O14467, O14468, O14469, O14470, O14471, O14472, O14473, O14474, O14475, O14476, O14477, O14478, O14479, O14480, O14481, O14482, O14483, O14484, O14485, O14486, O14487, O14488, O14489, O14490, O14491, O14492, O14493, O14494, O14495, O14496, O14497, O14498, O14499, O14500, O14501, O14502, O14503, O14504, O14505, O14506, O14507, O14508, O14509, O14510, O14511, O14512, O14513, O14514, O14515, O14516, O14517, O14518, O14519, O14520, O14521, O14522, O14523, O14524, O14525, O14526, O14527, O14528, O14529, O14530, O14531, O14532, O14533, O14534, O14535, O14536, O14537, O14538, O14539, O14540, O14541, O14542, O14543, O14544, O14545, O14546, O14547, O14548, O14549, O14550, O14551, O14552, O14553, O14554, O14555, O14556, O14557, O14558, O14559, O14560, O14561, O14562, O14563, O14564, O14565, O14566, O14567, O14568, O14569, O14570, O14571, O14572, O14573, O14574, O14575, O14576, O14577, O14578, O14579, O14580, O14581, O14582, O14583, O14584, O14585, O14586, O14587, O14588, O14589, O14590, O14591, O14592, O14593, O14594, O14595, O14596, O14597, O14598, O14599, O14600, O14601, O14602, O14603, O14604, O14605, O14606, O14607, O14608, O14609, O14610, O14611, O14612, O14613, O14614, O14615, O14616, O14617, O14618, O14619, O14620, O14621, O14622, O14623, O14624, O14625, O14626, O14627, O14628, O14629, O14630, O14631, O14632, O14633, O14634, O14635, O14636, O14637, O14638, O14639, O14640, O14641, O14642, O14643, O14644, O14645, O14646, O14647, O14648, O14649, O14650, O14651, O14652, O14653, O14654, O14655, O14656, O14657, O14658, O14659, O14660, O14661, O14662, O14663, O14664, O14665, O14666, O14667, O14668, O14669, O14670, O14671, O14672, O14673, O14674, O14675, O14676, O14677, O14678, O14679, O14680, O14681, O14682, O14683, O14684, O14685, O14686, O14687, O14688, O14689, O14690, O14691, O14692, O14693, O14694, O14695, O14696, O14697, O14698, O14699, O14700, O14701, O14702, O14703, O14704, O14705, O14706, O14707, O14708, O14709, O14710, O14711, O14712, O14713, O14714, O14715, O14716, O14717, O14718, O14719, O14720, O14721, O14722, O14723, O14724, O14725, O14726, O14727, O14728, O14729, O14730, O14731, O14732, O14733, O14734, O14735, O14736, O14737, O14738, O14739, O14740, O14741, O14742, O14743, O14744, O14745, O14746, O14747, O14748, O14749, O14750, O14751, O14752, O14753, O14754, O14755, O14756, O14757, O14758, O14759, O14760, O14761, O14762, O14763, O14764, O14765, O14766, O14767, O14768, O14769, O14770, O14771, O14772, O14773, O14774, O14775, O14776, O14777, O14778, O14779, O14780, O14781, O14782, O14783, O14784, O14785, O14786, O14787, O14788, O14789, O14790, O14791, O14792, O14793, O14794, O14795, O14796, O14797, O14798, O14799, O14800, O14801, O14802, O14803, O14804, O14805, O14806, O14807, O14808, O14809, O14810, O14811, O14812, O14813, O14814, O14815, O14816, O14817, O14818, O14819, O14820, O14821, O14822, O14823, O14824, O14825, O14826, O14827, O14828, O14829, O14830, O14831, O14832, O14833, O14834, O14835, O14836, O14837, O14838, O14839, O14840, O14841, O14842, O14843, O14844, O14845, O14846, O14847, O14848, O14849, O14850, O14851, O14852, O14853, O14854, O14855, O14856, O14857, O14858, O14859, O14860, O14861, O14862, O14863, O14864, O14865, O14866, O14867, O14868, O14869, O14870, O14871, O14872, O14873, O14874, O14875, O14876, O14877, O14878, O14879, O14880, O14881, O14882, O14883, O14884, O14885, O14886, O14887, O14888, O14889, O14890, O14891, O14892, O14893, O14894, O14895, O14896, O14897, O14898, O14899, O14900, O14901, O14902, O14903, O14904, O14905, O14906, O14907, O14908, O14909, O14910, O14911, O14912, O14913, O14914, O14915, O14916, O14917, O14918, O14919, O14920, O14921, O14922, O14923, O14924, O14925, O14926, O14927, O14928, O14929, O14930, O14931, O14932, O14933, O14934, O14935, O14936, O14937, O14938, O14939, O14940, O14941, O14942, O14943, O14944, O14945, O14946, O14947, O14948, O14949, O14950, O14951, O14952, O14953, O14954, O14955, O14956, O14957, O14958, O14959, O14960, O14961, O14962, O14963, O14964, O14965, O14966, O14967, O14968, O14969, O14970, O14971, O14972, O14973, O14974, O14975, O14976, O14977, O14978, O14979, O14980, O14981, O14982, O14983, O14984, O14985, O14986, O14987, O14988, O14989, O14990, O14991, O14992, O14993, O14994, O14995, O14996, O14997, O14998, O14999, O15000, O15001, O15002, O15003, O15004, O15005, O15006, O15007, O15008, O15009, O15010, O15011, O15012, O15013, O15014, O15015, O15016, O15017, O15018, O15019, O15020, O15021, O15022, O15023, O15024, O15025, O15026, O15027, O15028, O15029, O15030, O15031, O15032, O15033, O15034, O15035, O15036, O15037, O15038, O15039, O15040, O15041, O15042, O15043, O15044, O15045, O15046, O15047, O15048, O15049, O15050, O15051, O15052, O15053, O15054, O15055, O15056, O15057, O15058, O15059, O15060, O15061, O15062, O15063, O15064, O15065, O15066, O15067, O15068, O15069, O15070, O15071, O15072, O15073, O15074, O15075, O15076, O15077, O15078, O15079, O15080, O15081, O15082, O15083, O15084, O15085, O15086, O15087, O15088, O15089, O15090, O15091, O15092, O15093, O15094, O15095, O15096, O15097, O15098, O15099, O15100, O15101, O15102, O15103, O15104, O15105, O15106, O15107, O15108, O15109, O15110, O15111, O15112, O15113, O15114, O15115, O15116, O15117, O15118, O15119, O15120, O15121, O15122, O15123, O15124, O15125, O15126, O15127, O15128, O15129, O15130, O15131, O15132, O15133, O15134, O15135, O15136, O15137, O15138, O15139, O15140, O15141, O15142, O15143, O15144, O15145, O15146, O15147, O15148, O15149, O15150, O15151, O15152, O15153, O15154, O15155, O15156, O15157, O15158, O15159, O15160, O15161, O15162, O15163, O15164, O15165, O15166, O15167, O15168, O15169, O15170, O15171, O15172, O15173, O15174, O15175, O15176, O15177, O15178, O15179, O15180, O15181, O15182, O15183, O15184, O15185, O15186, O15187, O15188, O15189, O15190, O15191, O15192, O15193, O15194, O15195, O15196, O15197, O15198, O15199, O15200, O15201, O15202, O15203, O15204, O15205, O15206, O15207, O15208, O15209, O15210, O15211, O15212, O15213, O15214, O15215, O15216, O15217, O15218, O15219, O15220, O15221, O15222, O15223, O15224, O15225, O15226, O15227, O15228, O15229, O15230, O15231, O15232, O15233, O15234, O15235, O15236, O15237, O15238, O15239, O15240, O15241, O15242, O15243, O15244, O15245, O15246, O15247, O15248, O15249, O15250, O15251, O15252, O15253, O15254, O15255, O15256, O15257, O15258, O15259, O15260, O15261, O15262, O15263, O15264, O15265, O15266, O15267, O15268, O15269, O15270, O15271, O15272, O15273, O15274, O15275, O15276, O15277, O15278, O15279, O15280, O15281, O15282, O15283, O15284, O15285, O15286, O15287, O15288, O15289, O15290, O15291, O15292, O15293, O15294, O15295, O15296, O15297, O15298, O15299, O15300, O15301, O15302, O15303, O15304, O15305, O15306, O15307, O15308, O15309, O15310, O15311, O15312, O15313, O15314, O15315, O15316, O15317, O15318, O15319, O15320, O15321, O15322, O15323, O15324, O15325, O15326, O15327, O15328, O15329, O15330, O15331, O15332, O15333, O15334, O15335, O15336, O15337, O15338, O15339, O15340, O15341, O15342, O15343, O15344, O15345, O15346, O15347, O15348, O15349, O15350, O15351, O15352, O15353, O15354, O15355, O15356, O15357, O15358, O15359, O15360, O15361, O15362, O15363, O15364, O15365, O15366, O15367, O15368, O15369, O15370, O15371, O15372, O15373, O15374, O15375, O15376, O15377, O15378, O15379, O15380, O15381, O15382, O15383, O15384, O15385, O15386, O15387, O15388, O15389, O15390, O15391, O15392, O15393, O15394, O15395, O15396, O15397, O15398, O15399, O15400, O15401, O15402, O15403, O15404, O15405, O15406, O15407, O15408, O15409, O15410, O15411, O15412, O15413, O15414, O15415, O15416, O15417, O15418, O15419, O15420, O15421, O15422, O15423, O15424, O15425, O15426, O15427, O15428, O15429, O15430, O15431, O15432, O15433, O15434, O15435, O15436, O15437, O15438, O15439, O15440, O15441, O15442, O15443, O15444, O15445, O15446, O15447, O15448, O15449, O15450, O15451, O15452, O15453, O15454, O15455, O15456, O15457, O15458, O15459, O15460, O15461, O15462, O15463, O15464, O15465, O15466, O15467, O15468, O15469, O15470, O15471, O15472, O15473, O15474, O15475, O15476, O15477, O15478, O15479, O15480, O15481, O15482, O15483, O15484, O15485, O15486, O15487, O15488, O15489, O15490, O15491, O15492, O15493, O15494, O15495, O15496, O15497, O15498, O15499, O15500, O15501, O15502, O15503, O15504, O15505, O15506, O15507, O15508, O15509, O15510, O15511, O15512, O15513, O15514, O15515, O15516, O15517, O15518, O15519, O15520, O15521, O15522, O15523, O15524, O15525, O15526, O15527, O15528, O15529, O15530, O15531, O15532, O15533, O15534, O15535, O15536, O15537, O15538, O15539, O15540, O15541, O15542, O15543, O15544, O15545, O15546, O15547, O15548, O15549, O15550, O15551, O15552, O15553, O15554, O15555, O15556, O15557, O15558, O15559, O15560, O15561, O15562, O15563, O15564, O15565, O15566, O15567, O15568, O15569, O15570, O15571, O15572, O15573, O15574, O15575, O15576, O15577, O15578, O15579, O15580, O15581, O15582, O15583, O15584, O15585, O15586, O15587, O15588, O15589, O15590, O15591, O15592, O15593, O15594, O15595, O15596, O15597, O15598, O15599, O15600, O15601, O15602, O15603, O15604, O15605, O15606, O15607, O15608, O15609, O15610, O15611, O15612, O15613, O15614, O15615, O15616, O15617, O15618, O15619, O15620, O15621, O15622, O15623, O15624, O15625, O15626, O15627, O15628, O15629, O15630, O15631, O15632, O15633, O15634, O15635, O15636, O15637, O15638, O15639, O15640, O15641, O15642, O15643, O15644, O15645, O15646, O15647, O15648, O15649, O15650, O15651, O15652, O15653, O15654, O15655, O15656, O15657, O15658, O15659, O15660, O15661, O15662, O15663, O15664, O15665, O15666, O15667, O15668, O15669, O15670, O15671, O15672, O15673, O15674, O15675, O15676, O15677, O15678, O15679, O15680, O15681, O15682, O15683, O15684, O15685, O15686, O15687, O15688, O15689, O15690, O15691, O15692, O15693, O15694, O15695, O15696, O15697, O15698, O15699, O15700, O15701, O15702, O15703, O15704, O15705, O15706, O15707, O15708, O15709, O15710, O15711, O15712, O15713, O15714, O15715, O15716, O15717, O15718, O15719, O15720, O15721, O15722, O15723, O15724, O15725, O15726, O15727, O15728, O15729, O15730, O15731, O15732, O15733, O15734, O15735, O15736, O15737, O15738, O15739, O15740, O15741, O15742, O15743, O15744, O15745, O15746, O15747, O15748, O15749, O15750, O15751, O15752, O15753, O15754, O15755, O15756, O15757, O15758, O15759, O15760, O15761, O15762, O15763, O15764, O15765, O15766, O15767, O15768, O15769, O15770, O15771, O15772, O15773, O15774, O15775, O15776, O15777, O15778, O15779, O15780, O15781, O15782, O15783, O15784, O15785, O15786, O15787, O15788, O15789, O15790, O15791, O15792, O15793, O15794, O15795, O15796, O15797, O15798, O15799, O15800, O15801, O15802, O15803, O15804, O15805, O15806, O15807, O15808, O15809, O15810, O15811, O15812, O15813, O15814, O15815, O15816, O15817, O15818, O15819, O15820, O15821, O15822, O15823, O15824, O15825, O15826, O15827, O15828, O15829, O15830, O15831, O15832, O15833, O15834, O15835, O15836, O15837, O15838, O15839, O15840, O15841, O15842, O15843, O15844, O15845, O15846, O15847, O15848, O15849, O15850, O15851, O15852, O15853, O15854, O15855, O15856, O15857, O15858, O15859, O15860, O15861, O15862, O15863, O15864, O15865, O15866, O15867, O15868, O15869, O15870, O15871, O15872, O15873, O15874, O15875, O15876, O15877, O15878, O15879, O15880, O15881, O15882, O15883, O15884, O15885, O15886, O15887, O15888, O15889, O15890, O15891, O15892, O15893, O15894, O15895, O15896, O15897, O15898, O15899, O15900, O15901, O15902, O15903, O15904, O15905, O15906, O15907, O15908, O15909, O15910, O15911, O15912, O15913, O15914, O15915, O15916, O15917, O15918, O15919, O15920, O15921, O15922, O15923, O15924, O15925, O15926, O15927, O15928, O15929, O15930, O15931, O15932, O15933, O15934, O15935, O15936, O15937, O15938, O15939, O15940, O15941, O15942, O15943, O15944, O15945, O15946, O15947, O15948, O15949, O15950, O15951, O15952, O15953, O15954, O15955, O15956, O15957, O15958, O15959, O15960, O15961, O15962, O15963, O15964, O15965, O15966, O15967, O15968, O15969, O15970, O15971, O15972, O15973, O15974, O15975, O15976, O15977, O15978, O15979, O15980, O15981, O15982, O15983, O15984, O15985, O15986, O15987, O15988, O15989, O15990, O15991, O15992, O15993, O15994, O15995, O15996, O15997, O15998, O15999, O16000, O16001, O16002, O16003, O16004, O16005, O16006, O16007, O16008, O16009, O16010, O16011, O16012, O16013, O16014, O16015, O16016, O16017, O16018, O16019, O16020, O16021, O16022, O16023, O16024, O16025, O16026, O16027, O16028, O16029, O16030, O16031, O16032, O16033, O16034, O16035, O16036, O16037, O16038, O16039, O16040, O16041, O16042, O16043, O16044, O16045, O16046, O16047, O16048, O16049, O16050, O16051, O16052, O16053, O16054, O16055, O16056, O16057, O16058, O16059, O16060, O16061, O16062, O16063, O16064, O16065, O16066, O16067, O16068, O16069, O16070, O16071, O16072, O16073, O16074, O16075, O16076, O16077, O16078, O16079, O16080, O16081, O16082, O16083, O16084, O16085, O16086, O16087, O16088, O16089, O16090, O16091, O16092, O16093, O16094, O16095, O16096, O16097, O16098, O16099, O16100, O16101, O16102, O16103, O16104, O16105, O16106, O16107, O16108, O16109, O16110, O16111, O16112, O16113, O16114, O16115, O16116, O16117, O16118, O16119, O16120, O16121, O16122, O16123, O16124, O16125, O16126, O16127, O16128, O16129, O16130, O16131, O16132, O16133, O16134, O16135, O16136, O16137, O16138, O16139, O16140, O16141, O16142, O16143, O16144, O16145, O16146, O16147, O16148, O16149, O16150, O16151, O16152, O16153, O16154, O16155, O16156, O16157, O16158, O16159, O16160, O16161, O16162, O16163, O16164, O16165, O16166, O16167, O16168, O16169, O16170, O16171, O16172, O16173, O16174, O16175, O16176, O16177, O16178, O16179, O16180, O16181, O16182, O16183, O16184, O16185, O16186, O16187, O16188, O16189, O16190, O16191, O16192, O16193, O16194, O16195, O16196, O16197, O16198, O16199, O16200, O16201, O16202, O16203, O16204, O16205, O16206, O16207, O16208, O16209, O16210, O16211, O16212, O16213, O16214, O16215, O16216, O16217, O16218, O16219, O16220, O16221, O16222, O16223, O16224, O16225, O16226, O16227, O16228, O16229, O16230, O16231, O16232, O16233, O16234, O16235, O16236, O16237, O16238, O16239, O16240, O16241, O16242, O16243, O16244, O16245, O16246, O16247, O16248, O16249, O16250, O16251, O16252, O16253, O16254, O16255, O16256, O16257, O16258, O16259, O16260, O16261, O16262, O16263, O16264, O16265, O16266, O16267, O16268, O16269, O16270, O16271, O16272, O16273, O16274, O16275, O16276, O16277, O16278, O16279, O16280, O16281, O16282, O16283, O16284, O16285, O16286, O16287, O16288, O16289, O16290, O16291, O16292, O16293, O16294, O16295, O16296, O16297, O16298, O16299, O16300, O16301, O16302, O16303, O16304, O16305, O16306, O16307, O16308, O16309, O16310, O16311, O16312, O16313, O16314, O16315, O16316, O16317, O16318, O16319, O16320, O16321, O16322, O16323, O16324, O16325, O16326, O16327, O16328, O16329, O16330, O16331, O16332, O16333, O16334, O16335, O16336, O16337, O16338, O16339, O16340, O16341, O16342, O16343, O16344, O16345, O16346, O16347, O16348, O16349, O16350, O16351, O16352, O16353, O16354, O16355, O16356, O16357, O16358, O16359, O16360, O16361, O16362, O16363, O16364, O16365, O16366, O16367, O16368, O16369, O16370, O16371, O16372, O16373, O16374, O16375, O16376, O16377, O16378, O16379, O16380, O16381, O16382, O16383, O16384, O16385, O16386, O16387, O16388, O16389, O16390, O16391, O16392, O16393, O16394, O16395, O16396, O16397, O16398, O16399, O16400, O16401, O16402, O16403, O16404, O16405, O16406, O16407, O16408, O16409, O16410, O16411, O16412, O16413, O16414, O16415, O16416, O16417, O16418, O16419, O16420, O16421, O16422, O16423, O16424, O16425, O16426, O16427, O16428, O16429, O16430, O16431, O16432, O16433, O16434, O16435, O16436, O16437, O16438, O16439, O16440, O16441, O16442, O16443, O16444, O16445, O16446, O16447, O16448, O16449, O16450, O16451, O16452, O16453, O16454, O16455, O16456, O16457, O16458, O16459, O16460, O16461, O16462, O16463, O16464, O16465, O16466, O16467, O16468, O16469, O16470, O16471, O16472, O16473, O16474, O16475, O16476, O16477, O16478, O16479, O16480, O16481, O16482, O16483, O16484, O16485, O16486, O16487, O16488, O16489, O16490, O16491, O16492, O16493, O16494, O16495, O16496, O16497, O16498, O16499, O16500, O16501, O16502, O16503, O16504, O16505, O16506, O16507, O16508, O16509, O16510, O16511, O16512, O16513, O16514, O16515, O16516, O16517, O16518, O16519, O16520, O16521, O16522, O16523, O16524, O16525, O16526, O16527, O16528, O16529, O16530, O16531, O16532, O16533, O16534, O16535, O16536, O16537, O16538, O16539, O16540, O16541, O16542, O16543, O16544, O16545, O16546, O16547, O16548, O16549, O16550, O16551, O16552, O16553, O16554, O16555, O16556, O16557, O16558, O16559, O16560, O16561, O16562, O16563, O16564, O16565, O16566, O16567, O16568, O16569, O16570, O16571, O16572, O16573, O16574, O16575, O16576, O16577, O16578, O16579, O16580, O16581, O16582, O16583, O16584, O16585, O16586, O16587, O16588, O16589, O16590, O16591, O16592, O16593, O16594, O16595, O16596, O16597, O16598, O16599, O16600, O16601, O16602, O16603, O16604, O16605, O16606, O16607, O16608, O16609, O16610, O16611, O16612, O16613, O16614, O16615, O16616, O16617, O16618, O16619, O16620, O16621, O16622, O16623, O16624, O16625, O16626, O16627, O16628, O16629, O16630, O16631, O16632, O16633, O16634, O16635, O16636, O16637, O16638, O16639, O16640, O16641, O16642, O16643, O16644, O16645, O16646, O16647, O16648, O16649, O16650, O16651, O16652, O16653, O16654, O16655, O16656, O16657, O16658, O16659, O16660, O16661, O16662, O16663, O16664, O16665, O16666, O16667, O16668, O16669, O16670, O16671, O16672, O16673, O16674, O16675, O16676, O16677, O16678, O16679, O16680, O16681, O16682, O16683, O16684, O16685, O16686, O16687, O16688, O16689, O16690, O16691, O16692, O16693, O16694, O16695, O16696, O16697, O16698, O16699, O16700, O16701, O16702, O16703, O16704, O16705, O16706, O16707, O16708, O16709, O16710, O16711, O16712, O16713, O16714, O16715, O16716, O16717, O16718, O16719, O16720, O16721, O16722, O16723, O16724, O16725, O16726, O16727, O16728, O16729, O16730, O16731, O16732, O16733, O16734, O16735, O16736, O16737, O16738, O16739, O16740, O16741, O16742, O16743, O16744, O16745, O16746, O16747, O16748, O16749, O16750, O16751, O16752, O16753, O16754, O16755, O16756, O16757, O16758, O16759, O16760, O16761, O16762, O16763, O16764, O16765, O16766, O16767, O16768, O16769, O16770, O16771, O16772, O16773, O16774, O16775, O16776, O16777, O16778, O16779, O16780, O16781, O16782, O16783, O16784, O16785, O16786, O16787, O16788, O16789, O16790, O16791, O16792, O16793, O16794, O16795, O16796, O16797, O16798, O16799, O16800, O16801, O16802, O16803, O16804, O16805, O16806, O16807, O16808, O16809, O16810, O16811, O16812, O16813, O16814, O16815, O16816, O16817, O16818, O16819, O16820, O16821, O16822, O16823, O16824, O16825, O16826, O16827, O16828, O16829, O16830, O16831, O16832, O16833, O16834, O16835, O16836, O16837, O16838, O16839, O16840, O16841, O16842, O16843, O16844, O16845, O16846, O16847, O16848, O16849, O16850, O16851, O16852, O16853, O16854, O16855, O16856, O16857, O16858, O16859, O16860, O16861, O16862, O16863, O16864, O16865, O16866, O16867, O16868, O16869, O16870, O16871, O16872, O16873, O16874, O16875, O16876, O16877, O16878, O16879, O16880, O16881, O16882, O16883, O16884, O16885, O16886, O16887, O16888, O16889, O16890, O16891, O16892, O16893, O16894, O16895, O16896, O16897, O16898, O16899, O16900, O16901, O16902, O16903, O16904, O16905, O16906, O16907, O16908, O16909, O16910, O16911, O16912, O16913, O16914, O16915, O16916, O16917, O16918, O16919, O16920, O16921, O16922, O16923, O16924, O16925, O16926, O16927, O16928, O16929, O16930, O16931, O16932, O16933, O16934, O16935, O16936, O16937, O16938, O16939, O16940, O16941, O16942, O16943, O16944, O16945, O16946, O16947, O16948, O16949, O16950, O16951, O16952, O16953, O16954, O16955, O16956, O16957, O16958, O16959, O16960, O16961, O16962, O16963, O16964, O16965, O16966, O16967, O16968, O16969, O16970, O16971, O16972, O16973, O16974, O16975, O16976, O16977, O16978, O16979, O16980, O16981, O16982, O16983, O16984, O16985, O16986, O16987, O16988, O16989, O16990, O16991, O16992, O16993, O16994, O16995, O16996, O16997, O16998, O16999, O17000, O17001, O17002, O17003, O17004, O17005, O17006, O17007, O17008, O17009, O17010, O17011, O17012, O17013, O17014, O17015, O17016, O17017, O17018, O17019, O17020, O17021, O17022, O17023, O17024, O17025, O17026, O17027, O17028, O17029, O17030, O17031, O17032, O17033, O17034, O17035, O17036, O17037, O17038, O17039, O17040, O17041, O17042, O17043, O17044, O17045, O17046, O17047, O17048, O17049, O17050, O17051, O17052, O17053, O17054, O17055, O17056, O17057, O17058, O17059, O17060, O17061, O17062, O17063, O17064, O17065, O17066, O17067, O17068, O17069, O17070, O17071, O17072, O17073, O17074, O17075, O17076, O17077, O17078, O17079, O17080, O17081, O17082, O17083, O17084, O17085, O17086, O17087, O17088, O17089, O17090, O17091, O17092, O17093, O17094, O17095, O17096, O17097, O17098, O17099, O17100, O17101, O17102, O17103, O17104, O17105, O17106, O17107, O17108, O17109, O17110, O17111, O17112, O17113, O17114, O17115, O17116, O17117, O17118, O17119, O17120, O17121, O17122, O17123, O17124, O17125, O17126, O17127, O17128, O17129, O17130, O17131, O17132, O17133, O17134, O17135, O17136, O17137, O17138, O17139, O17140, O17141, O17142, O17143, O17144, O17145, O17146, O17147, O17148, O17149, O17150, O17151, O17152, O17153, O17154, O17155, O17156, O17157, O17158, O17159, O17160, O17161, O17162, O17163, O17164, O17165, O17166, O17167, O17168, O17169, O17170, O17171, O17172, O17173, O17174, O17175, O17176, O17177, O17178, O17179, O17180, O17181, O17182, O17183, O17184, O17185, O17186, O17187, O17188, O17189, O17190, O17191, O17192, O17193, O17194, O17195, O17196, O17197, O17198, O17199, O17200, O17201, O17202, O17203, O17204, O17205, O17206, O17207, O17208, O17209, O17210, O17211, O17212, O17213, O17214, O17215, O17216, O17217, O17218, O17219, O17220, O17221, O17222, O17223, O17224, O17225, O17226, O17227, O17228, O17229, O17230, O17231, O17232, O17233, O17234, O17235, O17236, O17237, O17238, O17239, O17240, O17241, O17242, O17243, O17244, O17245, O17246, O17247, O17248, O17249, O17250, O17251, O17252, O17253, O17254, O17255, O17256, O17257, O17258, O17259, O17260, O17261, O17262, O17263, O17264, O17265, O17266, O17267, O17268, O17269, O17270, O17271, O17272, O17273, O17274, O17275, O17276, O17277, O17278, O17279, O17280, O17281, O17282, O17283, O17284, O17285, O17286, O17287, O17288, O17289, O17290, O17291, O17292, O17293, O17294, O17295, O17296, O17297, O17298, O17299, O17300, O17301, O17302, O17303, O17304, O17305, O17306, O17307, O17308, O17309, O17310, O17311, O17312, O17313, O17314, O17315, O17316, O17317, O17318, O17319, O17320, O17321, O17322, O17323, O17324, O17325, O17326, O17327, O17328, O17329, O17330, O17331, O17332, O17333, O17334, O17335, O17336, O17337, O17338, O17339, O17340, O17341, O17342, O17343, O17344, O17345, O17346, O17347, O17348, O17349, O17350, O17351, O17352, O17353, O17354, O17355, O17356, O17357, O17358, O17359, O17360, O17361, O17362, O17363, O17364, O17365, O17366, O17367, O17368, O17369, O17370, O17371, O17372, O17373, O17374, O17375, O17376, O17377, O17378, O17379, O17380, O17381, O17382, O17383, O17384, O17385, O17386, O17387, O17388, O17389, O17390, O17391, O17392, O17393, O17394, O17395, O17396, O17397, O17398, O17399, O17400, O17401, O17402, O17403, O17404, O17405, O17406, O17407, O17408, O17409, O17410, O17411, O17412, O17413, O17414, O17415, O17416, O17417, O17418, O17419, O17420, O17421, O17422, O17423, O17424, O17425, O17426, O17427, O17428, O17429, O17430, O17431, O17432, O17433, O17434, O17435, O17436, O17437, O17438, O17439, O17440, O17441, O17442, O17443, O17444, O17445, O17446, O17447, O17448, O17449, O17450, O17451, O17452, O17453, O17454, O17455, O17456, O17457, O17458, O17459, O17460, O17461, O17462, O17463, O17464, O17465, O17466, O17467, O17468, O17469, O17470, O17471, O17472, O17473, O17474, O17475, O17476, O17477, O17478, O17479, O17480, O17481, O17482, O17483, O17484, O17485, O17486, O17487, O17488, O17489, O17490, O17491, O17492, O17493, O17494, O17495, O17496, O17497, O17498, O17499, O17500, O17501, O17502, O17503, O17504, O17505, O17506, O17507, O17508, O17509, O17510, O17511, O17512, O17513, O17514, O17515, O17516, O17517, O17518, O17519, O17520, O17521, O17522, O17523, O17524, O17525, O17526, O17527, O17528, O17529, O17530, O17531, O17532, O17533, O17534, O17535, O17536, O17537, O17538, O17539, O17540, O17541, O17542, O17543, O17544, O17545, O17546, O17547, O17548, O17549, O17550, O17551, O17552, O17553, O17554, O17555, O17556, O17557, O17558, O17559, O17560, O17561, O17562, O17563, O17564, O17565, O17566, O17567, O17568, O17569, O17570, O17571, O17572, O17573, O17574, O17575, O17576, O17577, O17578, O17579, O17580, O17581, O17582, O17583, O17584, O17585, O17586, O17587, O17588, O17589, O17590, O17591, O17592, O17593, O17594, O17595, O17596, O17597, O17598, O17599, O17600, O17601, O17602, O17603, O17604, O17605, O17606, O17607, O17608, O17609, O17610, O17611, O17612, O17613, O17614, O17615, O17616, O17617, O17618, O17619, O17620, O17621, O17622, O17623, O17624, O17625, O17626, O17627, O17628, O17629, O17630, O17631, O17632, O17633, O17634, O17635, O17636, O17637, O17638, O17639, O17640, O17641, O17642, O17643, O17644, O17645, O17646, O17647, O17648, O17649, O17650, O17651, O17652, O17653, O17654, O17655, O17656, O17657, O17658, O17659, O17660, O17661, O17662, O17663, O17664, O17665, O17666, O17667, O17668, O17669, O17670, O17671, O17672, O17673, O17674, O17675, O17676, O17677, O17678, O17679, O17680, O17681, O17682, O17683, O17684, O17685, O17686, O17687, O17688, O17689, O17690, O17691, O17692, O17693, O17694, O17695, O17696, O17697, O17698, O17699, O17700, O17701, O17702, O17703, O17704, O17705, O17706, O17707, O17708, O17709, O17710, O17711, O17712, O17713, O17714, O17715, O17716, O17717, O17718, O17719, O17720, O17721, O17722, O17723, O17724, O17725, O17726, O17727, O17728, O17729, O17730, O17731, O17732, O17733, O17734, O17735, O17736, O17737, O17738, O17739, O17740, O17741, O17742, O17743, O17744, O17745, O17746, O17747, O17748, O17749, O17750, O17751, O17752, O17753, O17754, O17755, O17756, O17757, O17758, O17759, O17760, O17761, O17762, O17763, O17764, O17765, O17766, O17767, O17768, O17769, O17770, O17771, O17772, O17773, O17774, O17775, O17776, O17777, O17778, O17779, O17780, O17781, O17782, O17783, O17784, O17785, O17786, O17787, O17788, O17789, O17790, O17791, O17792, O17793, O17794, O17795, O17796, O17797, O17798, O17799, O17800, O17801, O17802, O17803, O17804, O17805, O17806, O17807, O17808, O17809, O17810, O17811, O17812, O17813, O17814, O17815, O17816, O17817, O17818, O17819, O17820, O17821, O17822, O17823, O17824, O17825, O17826, O17827, O17828, O17829, O17830, O17831, O17832, O17833, O17834, O17835, O17836, O17837, O17838, O17839, O17840, O17841, O17842, O17843, O17844, O17845, O17846, O17847, O17848, O17849, O17850, O17851, O17852, O17853, O17854, O17855, O17856, O17857, O17858, O17859, O17860, O17861, O17862, O17863, O17864, O17865, O17866, O17867, O17868, O17869, O17870, O17871, O17872, O17873, O17874, O17875, O17876, O17877, O17878, O17879, O17880, O17881, O17882, O17883, O17884, O17885, O17886, O17887, O17888, O17889, O17890, O17891, O17892, O17893, O17894, O17895, O17896, O17897, O17898, O17899, O17900, O17901, O17902, O17903, O17904, O17905, O17906, O17907, O17908, O17909, O17910, O17911, O17912, O17913, O17914, O17915, O17916, O17917, O17918, O17919, O17920, O17921, O17922, O17923, O17924, O17925, O17926, O17927, O17928, O17929, O17930, O17931, O17932, O17933, O17934, O17935, O17936, O17937, O17938, O17939, O17940, O17941, O17942, O17943, O17944, O17945, O17946, O17947, O17948, O17949, O17950, O17951, O17952, O17953, O17954, O17955, O17956, O17957, O17958, O17959, O17960, O17961, O17962, O17963, O17964, O17965, O17966, O17967, O17968, O17969, O17970, O17971, O17972, O17973, O17974, O17975, O17976, O17977, O17978, O17979, O17980, O17981, O17982, O17983, O17984, O17985, O17986, O17987, O17988, O17989, O17990, O17991, O17992, O17993, O17994, O17995, O17996, O17997, O17998, O17999, O18000, O18001, O18002, O18003, O18004, O18005, O18006, O18007, O18008, O18009, O18010, O18011, O18012, O18013, O18014, O18015, O18016, O18017, O18018, O18019, O18020, O18021, O18022, O18023, O18024, O18025, O18026, O18027, O18028, O18029, O18030, O18031, O18032, O18033, O18034, O18035, O18036, O18037, O18038, O18039, O18040, O18041, O18042, O18043, O18044, O18045, O18046, O18047, O18048, O18049, O18050, O18051, O18052, O18053, O18054, O18055, O18056, O18057, O18058, O18059, O18060, O18061, O18062, O18063, O18064, O18065, O18066, O18067, O18068, O18069, O18070, O18071, O18072, O18073, O18074, O18075, O18076, O18077, O18078, O18079, O18080, O18081, O18082, O18083, O18084, O18085, O18086, O18087, O18088, O18089, O18090, O18091, O18092, O18093, O18094, O18095, O18096, O18097, O18098, O18099, O18100, O18101, O18102, O18103, O18104, O18105, O18106, O18107, O18108, O18109, O18110, O18111, O18112, O18113, O18114, O18115, O18116, O18117, O18118, O18119, O18120, O18121, O18122, O18123, O18124, O18125, O18126, O18127, O18128, O18129, O18130, O18131, O18132, O18133, O18134, O18135, O18136, O18137, O18138, O18139, O18140, O18141, O18142, O18143, O18144, O18145, O18146, O18147, O18148, O18149, O18150, O18151, O18152, O18153, O18154, O18155, O18156, O18157, O18158, O18159, O18160, O18161, O18162, O18163, O18164, O18165, O18166, O18167, O18168, O18169, O18170, O18171, O18172, O18173, O18174, O18175, O18176, O18177, O18178, O18179, O18180, O18181, O18182, O18183, O18184, O18185, O18186, O18187, O18188, O18189, O18190, O18191, O18192, O18193, O18194, O18195, O18196, O18197, O18198, O18199, O18200, O18201, O18202, O18203, O18204, O18205, O18206, O18207, O18208, O18209, O18210, O18211, O18212, O18213, O18214, O18215, O18216, O18217, O18218, O18219, O18220, O18221, O18222, O18223, O18224, O18225, O18226, O18227, O18228, O18229, O18230, O18231, O18232, O18233, O18234, O18235, O18236, O18237, O18238, O18239, O18240, O18241, O18242, O18243, O18244, O18245, O18246, O18247, O18248, O18249, O18250, O18251, O18252, O18253, O18254, O18255, O18256, O18257, O18258, O18259, O18260, O18261, O18262, O18263, O18264, O18265, O18266, O18267, O18268, O18269, O18270, O18271, O18272, O18273, O18274, O18275, O18276, O18277, O18278, O18279, O18280, O18281, O18282, O18283, O18284, O18285, O18286, O18287, O18288, O18289, O18290, O18291, O18292, O18293, O18294, O18295, O18296, O18297, O18298, O18299, O18300, O18301, O18302, O18303, O18304, O18305, O18306, O18307, O18308, O18309, O18310, O18311, O18312, O18313, O18314, O18315, O18316, O18317, O18318, O18319, O18320, O18321, O18322, O18323, O18324, O18325, O18326, O18327, O18328, O18329, O18330, O18331, O18332, O18333, O18334, O18335, O18336, O18337, O18338, O18339, O18340, O18341, O18342, O18343, O18344, O18345, O18346, O18347, O18348, O18349, O18350, O18351, O18352, O18353, O18354, O18355, O18356, O18357, O18358, O18359, O18360, O18361, O18362, O18363, O18364, O18365, O18366, O18367, O18368, O18369, O18370, O18371, O18372, O18373, O18374, O18375, O18376, O18377, O18378, O18379, O18380, O18381, O18382, O18383, O18384, O18385, O18386, O18387, O18388, O18389, O18390, O18391, O18392, O18393, O18394, O18395, O18396, O18397, O18398, O18399, O18400, O18401, O18402, O18403, O18404, O18405, O18406, O18407, O18408, O18409, O18410, O18411, O18412, O18413, O18414, O18415, O18416, O18417, O18418, O18419, O18420, O18421, O18422, O18423, O18424, O18425, O18426, O18427, O18428, O18429, O18430, O18431, O18432, O18433, O18434, O18435, O18436, O18437, O18438, O18439, O18440, O18441, O18442, O18443, O18444, O18445, O18446, O18447, O18448, O18449, O18450, O18451, O18452, O18453, O18454, O18455, O18456, O18457, O18458, O18459, O18460, O18461, O18462, O18463, O18464, O18465, O18466, O18467, O18468, O18469, O18470, O18471, O18472, O18473, O18474, O18475, O18476, O18477, O18478, O18479, O18480, O18481, O18482, O18483, O18484, O18485, O18486, O18487, O18488, O18489, O18490, O18491, O18492, O18493, O18494, O18495, O18496, O18497, O18498, O18499, O18500, O18501, O18502, O18503, O18504, O18505, O18506, O18507, O18508, O18509, O18510, O18511, O18512, O18513, O18514, O18515, O18516, O18517, O18518, O18519, O18520, O18521, O18522, O18523, O18524, O18525, O18526, O18527, O18528, O18529, O18530, O18531, O18532, O18533, O18534, O18535, O18536, O18537, O18538, O18539, O18540, O18541, O18542, O18543, O18544, O18545, O18546, O18547, O18548, O18549, O18550, O18551, O18552, O18553, O18554, O18555, O18556, O18557, O18558, O18559, O18560, O18561, O18562, O18563, O18564, O18565, O18566, O18567, O18568, O18569, O18570, O18571, O18572, O18573, O18574, O18575, O18576, O18577, O18578, O18579, O18580, O18581, O18582, O18583, O18584, O18585, O18586, O18587, O18588, O18589, O18590, O18591, O18592, O18593, O18594, O18595, O18596, O18597, O18598, O18599, O18600, O18601, O18602, O18603, O18604, O18605, O18606, O18607, O18608, O18609, O18610, O18611, O18612, O18613, O18614, O18615, O18616, O18617, O18618, O18619, O18620, O18621, O18622, O18623, O18624, O18625, O18626, O18627, O18628, O18629, O18630, O18631, O18632, O18633, O18634, O18635, O18636, O18637, O18638, O18639, O18640, O18641, O18642, O18643, O18644, O18645, O18646, O18647, O18648, O18649, O18650, O18651, O18652, O18653, O18654, O18655, O18656, O18657, O18658, O18659, O18660, O18661, O18662, O18663, O18664, O18665, O18666, O18667, O18668, O18669, O18670, O18671, O18672, O18673, O18674, O18675, O18676, O18677, O18678, O18679, O18680, O18681, O18682, O18683, O18684, O18685, O18686, O18687, O18688, O18689, O18690, O18691, O18692, O18693, O18694, O18695, O18696, O18697, O18698, O18699, O18700, O18701, O18702, O18703, O18704, O18705, O18706, O18707, O18708, O18709, O18710, O18711, O18712, O18713, O18714, O18715, O18716, O18717, O18718, O18719, O18720, O18721, O18722, O18723, O18724, O18725, O18726, O18727, O18728, O18729, O18730, O18731, O18732, O18733, O18734, O18735, O18736, O18737, O18738, O18739, O18740, O18741, O18742, O18743, O18744, O18745, O18746, O18747, O18748, O18749, O18750, O18751, O18752, O18753, O18754, O18755, O18756, O18757, O18758, O18759, O18760, O18761, O18762, O18763, O18764, O18765, O18766, O18767, O18768, O18769, O18770, O18771, O18772, O18773, O18774, O18775, O18776, O18777, O18778, O18779, O18780, O18781, O18782, O18783, O18784, O18785, O18786, O18787, O18788, O18789, O18790, O18791, O18792, O18793, O18794, O18795, O18796, O18797, O18798, O18799, O18800, O18801, O18802, O18803, O18804, O18805, O18806, O18807, O18808, O18809, O18810, O18811, O18812, O18813, O18814, O18815, O18816, O18817, O18818, O18819, O18820, O18821, O18822, O18823, O18824, O18825, O18826, O18827, O18828, O18829, O18830, O18831, O18832, O18833, O18834, O18835, O18836, O18837, O18838, O18839, O18840, O18841, O18842, O18843, O18844, O18845, O18846, O18847, O18848, O18849, O18850, O18851, O18852, O18853, O18854, O18855, O18856, O18857, O18858, O18859, O18860, O18861, O18862, O18863, O18864, O18865, O18866, O18867, O18868, O18869, O18870, O18871, O18872, O18873, O18874, O18875, O18876, O18877, O18878, O18879, O18880, O18881, O18882, O18883, O18884, O18885, O18886, O18887, O18888, O18889, O18890, O18891, O18892, O18893, O18894, O18895, O18896, O18897, O18898, O18899, O18900, O18901, O18902, O18903, O18904, O18905, O18906, O18907, O18908, O18909, O18910, O18911, O18912, O18913, O18914, O18915, O18916, O18917, O18918, O18919, O18920, O18921, O18922, O18923, O18924, O18925, O18926, O18927, O18928, O18929, O18930, O18931, O18932, O18933, O18934, O18935, O18936, O18937, O18938, O18939, O18940, O18941, O18942, O18943, O18944, O18945, O18946, O18947, O18948, O18949, O18950, O18951, O18952, O18953, O18954, O18955, O18956, O18957, O18958, O18959, O18960, O18961, O18962, O18963, O18964, O18965, O18966, O18967, O18968, O18969, O18970, O18971, O18972, O18973, O18974, O18975, O18976, O18977, O18978, O18979, O18980, O18981, O18982, O18983, O18984, O18985, O18986, O18987, O18988, O18989, O18990, O18991, O18992, O18993, O18994, O18995, O18996, O18997, O18998, O18999, O19000, O19001, O19002, O19003, O19004, O19005, O19006, O19007, O19008, O19009, O19010, O19011, O19012, O19013, O19014, O19015, O19016, O19017, O19018, O19019, O19020, O19021, O19022, O19023, O19024, O19025, O19026, O19027, O19028, O19029, O19030, O19031, O19032, O19033, O19034, O19035, O19036, O19037, O19038, O19039, O19040, O19041, O19042, O19043, O19044, O19045, O19046, O19047, O19048, O19049, O19050, O19051, O19052, O19053, O19054, O19055, O19056, O19057, O19058, O19059, O19060, O19061, O19062, O19063, O19064, O19065, O19066, O19067, O19068, O19069, O19070, O19071, O19072, O19073, O19074, O19075, O19076, O19077, O19078, O19079, O19080, O19081, O19082, O19083, O19084, O19085, O19086, O19087, O19088, O19089, O19090, O19091, O19092, O19093, O19094, O19095, O19096, O19097, O19098, O19099, O19100, O19101, O19102, O19103, O19104, O19105, O19106, O19107, O19108, O19109, O19110, O19111, O19112, O19113, O19114, O19115, O19116, O19117, O19118, O19119, O19120, O19121, O19122, O19123, O19124, O19125, O19126, O19127, O19128, O19129, O19130, O19131, O19132, O19133, O19134, O19135, O19136, O19137, O19138, O19139, O19140, O19141, O19142, O19143, O19144, O19145, O19146, O19147, O19148, O19149, O19150, O19151, O19152, O19153, O19154, O19155, O19156, O19157, O19158, O19159, O19160, O19161, O19162, O19163, O19164, O19165, O19166, O19167, O19168, O19169, O19170, O19171, O19172, O19173, O19174, O19175, O19176, O19177, O19178, O19179, O19180, O19181, O19182, O19183, O19184, O19185, O19186, O19187, O19188, O19189, O19190, O19191, O19192, O19193, O19194, O19195, O19196, O19197, O19198, O19199, O19200, O19201, O19202, O19203, O19204, O19205, O19206, O19207, O19208, O19209, O19210, O19211, O19212, O19213, O19214, O19215, O19216, O19217, O19218, O19219, O19220, O19221, O19222, O19223, O19224, O19225, O19226, O19227, O19228, O19229, O19230, O19231, O19232, O19233, O19234, O19235, O19236, O19237, O19238, O19239, O19240, O19241, O19242, O19243, O19244, O19245, O19246, O19247, O19248, O19249, O19250, O19251, O19252, O19253, O19254, O19255, O19256, O19257, O19258, O19259, O19260, O19261, O19262, O19263, O19264, O19265, O19266, O19267, O19268, O19269, O19270, O19271, O19272, O19273, O19274, O19275, O19276, O19277, O19278, O19279, O19280, O19281, O19282, O19283, O19284, O19285, O19286, O19287, O19288, O19289, O19290, O19291, O19292, O19293, O19294, O19295, O19296, O19297, O19298, O19299, O19300, O19301, O19302, O19303, O19304, O19305, O19306, O19307, O19308, O19309, O19310, O19311, O19312, O19313, O19314, O19315, O19316, O19317, O19318, O19319, O19320, O19321, O19322, O19323, O19324, O19325, O19326, O19327, O19328, O19329, O19330, O19331, O19332, O19333, O19334, O19335, O19336, O19337, O19338, O19339, O19340, O19341, O19342, O19343, O19344, O19345, O19346, O19347, O19348, O19349, O19350, O19351, O19352, O19353, O19354, O19355, O19356, O19357, O19358, O19359, O19360, O19361, O19362, O19363, O19364, O19365, O19366, O19367, O19368, O19369, O19370, O19371, O19372, O19373, O19374, O19375, O19376, O19377, O19378, O19379, O19380, O19381, O19382, O19383, O19384, O19385, O19386, O19387, O19388, O19389, O19390, O19391, O19392, O19393, O19394, O19395, O19396, O19397, O19398, O19399, O19400, O19401, O19402, O19403, O19404, O19405, O19406, O19407, O19408, O19409, O19410, O19411, O19412, O19413, O19414, O19415, O19416, O19417, O19418, O19419, O19420, O19421, O19422, O19423, O19424, O19425, O19426, O19427, O19428, O19429, O19430, O19431, O19432, O19433, O19434, O19435, O19436, O19437, O19438, O19439, O19440, O19441, O19442, O19443, O19444, O19445, O19446, O19447, O19448, O19449, O19450, O19451, O19452, O19453, O19454, O19455, O19456, O19457, O19458, O19459, O19460, O19461, O19462, O19463, O19464, O19465, O19466, O19467, O19468, O19469, O19470, O19471, O19472, O19473, O19474, O19475, O19476, O19477, O19478, O19479, O19480, O19481, O19482, O19483, O19484, O19485, O19486, O19487, O19488, O19489, O19490, O19491, O19492, O19493, O19494, O19495, O19496, O19497, O19498, O19499, O19500, O19501, O19502, O19503, O19504, O19505, O19506, O19507, O19508, O19509, O19510, O19511, O19512, O19513, O19514, O19515, O19516, O19517, O19518, O19519, O19520, O19521, O19522, O19523, O19524, O19525, O19526, O19527, O19528, O19529, O19530, O19531, O19532, O19533, O19534, O19535, O19536, O19537, O19538, O19539, O19540, O19541, O19542, O19543, O19544, O19545, O19546, O19547, O19548, O19549, O19550, O19551, O19552, O19553, O19554, O19555, O19556, O19557, O19558, O19559, O19560, O19561, O19562, O19563, O19564, O19565, O19566, O19567, O19568, O19569, O19570, O19571, O19572, O19573, O19574, O19575, O19576, O19577, O19578, O19579, O19580, O19581, O19582, O19583, O19584, O19585, O19586, O19587, O19588, O19589, O19590, O19591, O19592, O19593, O19594, O19595, O19596, O19597, O19598, O19599, O19600, O19601, O19602, O19603, O19604, O19605, O19606, O19607, O19608, O19609, O19610, O19611, O19612, O19613, O19614, O19615, O19616, O19617, O19618, O19619, O19620, O19621, O19622, O19623, O19624, O19625, O19626, O19627, O19628, O19629, O19630, O19631, O19632, O19633, O19634, O19635, O19636, O19637, O19638, O19639, O19640, O19641, O19642, O19643, O19644, O19645, O19646, O19647, O19648, O19649, O19650, O19651, O19652, O19653, O19654, O19655, O19656, O19657, O19658, O19659, O19660, O19661, O19662, O19663, O19664, O19665, O19666, O19667, O19668, O19669, O19670, O19671, O19672, O19673, O19674, O19675, O19676, O19677, O19678, O19679, O19680, O19681, O19682, O19683, O19684, O19685, O19686, O19687, O19688, O19689, O19690, O19691, O19692, O19693, O19694, O19695, O19696, O19697, O19698, O19699, O19700, O19701, O19702, O19703, O19704, O19705, O19706, O19707, O19708, O19709, O19710, O19711, O19712, O19713, O19714, O19715, O19716, O19717, O19718, O19719, O19720, O19721, O19722, O19723, O19724, O19725, O19726, O19727, O19728, O19729, O19730, O19731, O19732, O19733, O19734, O19735, O19736, O19737, O19738, O19739, O19740, O19741, O19742, O19743, O19744, O19745, O19746, O19747, O19748, O19749, O19750, O19751, O19752, O19753, O19754, O19755, O19756, O19757, O19758, O19759, O19760, O19761, O19762;
  wire W12294, W38549, W21249, W12301, W12299, W12296, W12295, W21253, W12292, W29509, W12289, W12288, W29506, W12325, W38530, W12321, W21243, W38533, W29517, W29503, W38537, W12314, W38540, W12310, W12309, W12308, W21266, W21264, W12263, W12262, W12261, W12260, W38599, W38600, W38595, W12253, W29496, W21269, W29495, W38609, W12274, W29500, W38574, W38579, W12277, W38580, W38585, W29499, W38591, W21262, W12266, W38471, W29537, W12378, W21229, W12376, W12375, W12373, W12372, W12371, W38474, W38477, W12366, W12391, W12398, W38444, W21220, W12394, W29543, W12390, W29541, W29540, W29539, W12384, W12335, W12343, W12341, W12340, W12339, W12338, W12345, W12334, W29525, W12332, W12329, W38524, W12354, W12364, W21234, W38493, W12356, W29490, W38504, W38508, W12350, W21236, W12348, W38511, W12148, W12147, W12146, W12144, W12143, W12141, W12140, W38714, W12138, W12137, W38722, W21310, W12165, W29469, W21297, W21298, W12157, W29466, W21303, W12101, W12109, W12108, W12105, W38745, W29452, W38739, W29451, W29450, W12096, W38757, W12092, W29444, W38729, W12126, W12125, W12123, W29455, W12168, W12116, W12115, W12114, W12113, W38738, W12218, W21278, W29485, W38644, W29484, W12220, W38634, W12217, W12215, W12214, W12213, W38650, W12210, W38627, W38614, W12243, W12238, W38623, W21276, W12234, W12232, W12231, W29487, W38678, W12187, W12186, W12182, W21290, W12190, W12178, W38688, W12172, W12171, W12208, W38663, W38664, W12201, W12400, W38669, W21283, W12196, W21284, W38674, W21286, W21149, W12615, W12614, W21145, W38218, W12610, W29616, W29620, W12604, W38225, W21150, W12598, W38205, W12631, W21141, W12629, W12628, W12626, W29622, W12621, W12618, W38251, W38252, W21158, W38258, W38260, W21159, W12566, W21160, W38265, W38267, W12559, W12587, W38231, W12594, W29612, W12591, W12589, W38199, W29611, W38240, W12584, W38241, W12578, W38135, W38123, W12692, W12687, W38132, W12695, W38139, W12683, W38152, W29641, W12704, W12711, W12710, W21117, W38110, W12706, W12705, W12675, W12703, W12701, W21118, W12699, W29647, W12653, W38177, W38180, W12649, W12647, W29626, W12640, W29624, W38197, W12674, W12673, W38157, W29640, W12666, W38270, W12662, W38170, W21129, W12658, W12655, W12448, W38382, W12455, W29561, W12452, W21203, W12446, W12445, W38398, W12442, W12440, W38360, W38361, W12473, W12472, W12469, W12438, W38369, W12465, W21196, W38374, W38375, W12410, W12419, W12418, W12417, W12415, W21216, W12413, W21214, W12408, W21218, W12403, W12436, W12435, W29553, W12431, W12429, W29567, W29550, W21211, W12425, W21212, W29548, W12421, W12529, W29596, W29594, W38300, W12531, W12530, W21174, W38305, W38308, W12525, W38310, W21175, W21164, W12555, W38272, W38275, W12547, W29601, W12545, W29600, W12541, W12486, W12495, W12494, W29574, W12492, W12490, W12488, W29577, W12481, W21191, W29569, W38329, W12517, W12516, W12514, W38321, W38323, W12500, W38337, W38338, W29308, W11675, W11678, W39184, W11666, W39186, W11663, W11662, W39188, W39161, W11697, W21464, W11694, W11693, W11692, W29315, W11660, W11683, W11681, W11680, W11641, W11640, W11638, W11635, W29298, W29297, W39215, W11628, W39220, W39197, W11656, W29302, W21477, W11653, W11651, W39157, W11649, W11647, W11646, W11645, W11644, W29299, W11758, W21444, W11754, W39103, W21445, W21441, W39107, W39108, W11745, W11744, W21434, W11776, W11771, W11770, W11769, W21438, W29340, W11709, W21456, W39142, W29322, W39146, W11710, W11707, W11706, W21462, W11701, W11699, W11730, W21448, W39120, W11736, W21449, W29332, W29331, W39127, W39133, W11722, W11513, W11521, W11520, W39323, W11517, W29250, W39322, W21525, W11508, W21529, W39346, W11530, W39301, W21517, W11535, W29257, W11533, W11532, W39310, W39313, W39314, W39319, W11524, W11474, W11482, W29241, W11478, W11477, W11476, W39369, W39376, W11471, W21539, W11468, W11467, W21530, W21531, W11500, W11498, W29243, W11493, W39298, W11491, W11488, W21536, W21501, W11601, W21498, W11594, W11590, W39261, W39263, W29272, W11584, W11582, W39234, W11620, W39225, W29289, W11616, W21491, W11609, W29282, W11552, W39286, W11559, W29264, W11555, W11553, W11563, W39292, W11550, W39294, W29263, W29262, W11544, W11543, W11579, W39271, W11576, W11574, W29269, W39078, W11571, W11570, W39279, W11568, W11567, W39281, W21508, W38890, W38881, W21369, W11983, W29405, W11980, W21373, W11976, W38892, W38897, W11969, W38899, W29399, W11966, W11996, W38857, W21360, W21362, W11999, W11998, W29416, W38870, W38876, W38877, W11939, W11947, W11937, W21389, W11931, W11930, W38949, W29396, W38904, W38906, W21379, W29394, W21381, W11954, W38916, W38917, W29391, W11949, W21385, W12058, W38787, W12065, W21334, W12060, W12067, W12057, W38794, W12053, W29434, W12051, W38771, W38767, W12084, W12083, W12081, W12080, W12079, W21337, W21329, W12073, W21331, W12069, W12018, W38839, W12022, W29423, W12019, W21353, W21354, W29421, W12013, W21357, W38852, W12010, W12009, W21338, W12047, W21342, W21343, W12040, W38818, W21345, W21391, W12036, W21347, W38828, W11825, W11833, W11832, W11831, W11830, W11829, W11828, W11827, W39039, W39045, W11819, W11818, W11817, W21419, W39031, W39022, W21413, W39026, W11846, W21414, W11840, W11839, W21416, W11837, W39036, W39070, W11795, W11789, W21428, W21425, W11784, W11783, W11782, W21430, W39074, W21431, W11805, W21421, W11812, W21422, W11810, W11809, W11808, W39053, W29362, W11804, W29355, W11801, W11800, W11799, W11797, W11908, W21399, W11905, W38980, W29376, W11898, W38987, W11895, W11894, W38989, W11891, W11927, W29387, W29385, W11924, W29384, W11921, W38956, W38961, W21396, W38965, W11913, W11862, W11871, W11870, W11867, W21405, W11864, W11863, W29370, W39012, W11857, W11888, W11887, W11884, W38999, W11882, W39000, W11879, W11878, W11876, W39002, W11874, W11873, W20849, W37278, W13552, W13550, W37279, W20848, W13547, W13546, W37287, W20851, W37293, W13537, W37294, W13572, W13570, W13569, W13568, W13567, W13564, W13562, W13559, W13558, W37274, W13556, W13507, W13515, W13514, W20857, W13512, W13511, W13510, W20860, W29908, W13501, W37338, W37307, W13533, W37301, W37304, W13573, W37308, W37309, W20855, W13519, W29913, W37215, W13627, W13626, W13625, W13624, W37214, W13622, W37208, W13620, W20831, W29938, W13616, W29936, W37224, W13648, W13646, W13645, W37186, W37191, W13639, W20825, W20826, W37198, W29941, W37255, W13593, W13591, W37249, W37252, W37245, W20841, W13581, W37258, W37259, W29929, W37261, W29928, W13611, W13609, W13608, W13607, W13605, W37233, W13496, W29870, W13396, W37445, W20890, W20891, W29871, W13389, W37456, W13385, W37457, W37462, W13380, W13407, W13416, W37426, W13414, W13411, W37432, W37435, W13378, W13406, W13404, W29876, W37441, W13401, W13400, W13356, W29859, W29858, W13353, W13352, W20906, W20908, W13347, W13343, W29847, W13366, W29867, W13373, W13372, W13370, W37472, W29879, W13364, W13363, W13360, W37479, W37368, W13472, W29894, W37372, W13468, W29892, W37367, W13462, W13461, W37383, W13456, W37351, W13495, W13493, W13491, W13490, W13486, W37387, W37354, W13481, W29896, W37418, W13432, W37414, W13429, W20880, W13426, W29881, W37423, W13420, W13419, W37396, W20875, W13450, W13449, W13448, W13649, W37401, W13439, W13438, W13437, W36972, W13868, W13867, W30024, W13864, W13861, W20746, W36974, W13856, W36977, W30025, W13884, W36938, W13882, W20743, W13879, W13851, W36955, W20744, W13874, W20745, W20761, W13826, W13824, W13823, W20759, W13819, W37006, W13816, W30005, W30003, W13811, W20766, W37001, W13850, W30019, W13845, W36990, W13842, W36936, W37002, W13831, W13830, W13829, W13828, W13940, W36880, W13938, W13936, W36881, W13941, W13931, W30039, W36890, W13926, W13925, W13924, W36863, W13954, W13953, W36862, W36892, W30041, W13896, W30030, W13901, W13900, W13899, W36926, W13895, W13894, W13893, W13891, W30035, W13919, W36897, W13917, W13806, W36908, W20737, W36911, W36912, W20738, W13906, W37135, W13708, W37130, W13704, W20803, W13702, W37134, W37126, W13699, W13698, W20805, W37139, W13693, W13692, W13691, W29955, W13717, W13726, W13725, W37115, W13723, W29961, W13718, W20801, W37122, W13714, W20802, W37124, W13711, W37175, W13669, W13665, W13664, W20818, W20820, W13653, W20821, W37149, W13687, W37144, W37145, W37147, W13683, W37148, W13681, W37111, W20808, W20812, W29952, W13672, W13786, W37043, W20774, W13782, W37046, W37049, W13779, W37042, W13776, W29989, W13772, W20780, W37059, W13769, W29998, W20769, W13803, W13801, W13800, W13799, W37035, W13795, W13793, W13792, W37041, W13789, W13746, W29976, W13742, W13740, W13747, W13735, W20794, W13733, W13732, W29965, W37103, W20796, W13756, W29982, W37068, W13762, W20784, W37072, W13757, W37510, W13753, W13751, W29977, W12919, W29719, W21040, W12926, W37899, W12924, W12920, W37895, W12917, W29715, W21043, W29714, W21045, W12911, W12947, W12946, W29723, W12943, W12941, W29711, W12933, W12931, W37951, W29705, W12888, W12883, W12890, W21058, W21059, W12875, W12872, W37962, W37929, W37914, W29710, W37923, W37926, W12901, W21034, W37932, W12895, W21051, W37941, W37942, W12994, W13002, W29740, W29739, W37837, W29738, W21022, W12993, W12991, W21024, W12986, W29743, W21012, W13017, W37823, W13015, W13014, W37825, W13009, W13008, W13006, W21017, W12957, W12965, W21032, W12963, W12961, W12960, W12958, W29728, W12956, W12955, W12954, W12953, W12951, W12950, W12975, W12981, W12980, W12979, W29732, W12977, W29731, W12870, W12974, W37859, W12972, W29729, W12967, W38055, W38051, W29661, W12770, W38054, W12767, W12774, W38056, W12763, W38062, W12759, W12757, W38032, W21089, W29668, W29667, W29660, W29664, W21095, W38049, W12776, W29662, W21110, W21111, W38094, W12726, W12723, W21114, W12719, W12718, W12714, W12754, W38072, W38074, W38076, W21104, W12793, W21106, W12739, W21107, W12841, W29688, W12849, W12848, W12846, W12844, W21069, W12840, W37987, W12838, W37990, W12835, W12832, W29692, W12869, W21062, W12866, W12865, W29695, W29694, W12861, W12830, W12859, W12858, W12856, W12855, W29691, W37975, W12803, W21084, W12808, W12807, W12806, W12804, W21083, W12802, W21086, W38024, W38025, W12796, W12820, W12828, W21076, W29682, W21079, W21080, W13022, W29678, W38010, W38012, W29676, W12814, W12813, W13229, W13237, W13236, W37597, W29812, W13233, W20947, W13230, W37595, W20949, W13224, W13223, W37612, W37615, W13255, W20941, W20942, W20943, W29807, W13246, W37592, W13244, W13199, W13197, W37626, W13190, W13189, W13188, W13187, W37642, W20954, W20952, W13216, W37618, W13213, W13211, W20953, W37579, W13207, W13206, W20955, W13204, W37625, W13202, W13306, W13316, W13315, W20927, W29833, W13307, W13304, W37545, W13300, W13299, W20919, W13334, W13333, W20917, W20918, W37517, W13326, W13294, W20920, W13322, W13318, W37566, W29822, W13270, W13269, W13268, W13267, W37564, W13265, W13264, W13263, W37572, W37573, W37557, W37554, W13291, W13287, W13286, W13285, W13182, W13283, W13280, W13277, W13072, W37767, W13082, W37771, W29763, W20998, W13065, W29761, W37778, W29771, W29777, W13101, W37736, W13099, W13098, W13096, W29772, W13062, W13091, W13088, W37752, W13083, W37796, W13043, W37797, W37801, W13035, W13031, W13029, W13027, W29752, W13024, W13061, W21001, W37785, W37787, W13047, W13046, W13152, W20965, W13157, W13155, W20968, W37681, W13150, W37682, W37685, W13144, W13179, W37649, W37650, W13174, W13141, W29800, W37658, W20963, W20984, W37710, W37718, W13114, W37709, W29780, W29779, W13108, W29778, W29790, W37692, W37695, W13136, W13135, W13134, W13131, W29789, W20976, W13127, W13123, W9802, W9810, W9809, W9808, W28729, W9803, W22051, W9797, W9796, W41079, W28733, W41072, W9822, W41114, W9818, W9817, W9814, W9813, W41134, W9770, W9769, W22057, W9762, W41149, W41154, W9757, W41117, W9789, W9788, W41125, W9781, W9779, W9778, W9777, W9776, W9885, W41026, W28750, W9881, W9880, W9878, W22034, W9886, W28747, W41038, W9873, W41040, W22036, W22037, W9868, W9901, W41012, W9899, W28753, W9896, W22038, W9893, W9891, W41022, W9887, W9838, W41054, W9846, W41056, W9843, W9842, W9841, W9840, W41053, W9837, W28735, W41064, W22047, W9830, W9856, W9866, W9865, W9863, W9862, W9860, W22040, W9855, W9854, W22042, W9852, W9643, W41266, W28677, W9645, W22095, W9653, W9640, W9638, W9635, W22087, W9672, W9670, W9667, W28680, W9633, W9661, W9660, W41258, W41261, W9656, W9654, W28664, W9611, W9609, W9608, W28665, W28669, W22112, W9592, W9586, W9624, W41280, W22097, W41287, W41288, W41290, W9621, W22100, W41293, W41294, W9615, W9719, W22072, W9725, W9724, W41203, W41192, W9718, W22077, W41207, W41209, W9714, W9712, W28692, W22064, W9755, W9754, W9753, W9746, W9745, W41216, W22069, W9732, W28687, W9691, W28689, W9689, W9688, W9687, W22084, W9685, W41235, W28686, W9680, W9679, W9678, W9675, W22081, W9708, W9706, W9705, W41219, W28691, W9701, W9904, W9698, W9696, W9695, W22082, W40771, W10112, W28823, W10110, W21959, W10107, W10106, W10115, W28821, W10103, W10102, W40781, W21961, W40757, W21952, W10130, W10129, W28825, W10125, W10122, W10121, W10119, W10068, W10075, W28816, W10073, W40813, W10070, W40815, W40816, W10064, W10061, W10059, W21964, W28820, W10094, W40792, W10089, W10088, W10085, W40798, W10083, W10081, W10192, W10190, W21932, W40688, W10186, W40693, W40695, W40684, W10174, W28852, W10215, W21922, W10213, W40669, W10208, W10202, W10200, W40681, W40683, W10194, W21942, W28834, W21946, W10147, W10145, W10142, W40747, W28832, W10139, W28831, W40752, W10135, W28829, W21941, W40714, W28840, W40716, W40721, W10165, W28838, W10162, W10161, W10160, W10156, W9955, W28774, W40950, W9959, W9957, W9953, W40957, W22013, W9948, W9947, W28780, W28785, W28783, W40923, W9977, W9946, W22005, W9974, W9972, W9971, W22007, W9969, W9967, W22022, W9923, W40996, W9921, W9920, W40999, W40990, W9913, W9912, W41003, W28757, W41005, W41006, W9906, W9944, W9941, W28765, W9938, W40982, W9930, W10032, W10040, W28802, W40854, W21984, W21986, W40867, W10024, W40833, W28808, W21974, W21975, W10052, W21976, W28799, W21978, W21979, W28804, W10044, W21981, W10003, W21994, W28793, W9999, W28791, W9997, W21997, W9993, W28786, W9990, W9988, W9987, W40913, W40886, W10021, W40876, W10019, W28798, W10015, W9585, W40888, W21991, W10008, W10006, W41749, W9167, W9164, W41747, W9162, W9161, W9158, W28499, W9156, W22266, W9154, W41751, W9151, W9150, W22267, W28500, W41735, W9181, W28503, W9178, W9177, W9175, W9174, W9173, W9172, W22262, W9170, W9169, W9126, W9124, W9121, W41791, W9118, W9128, W41800, W28483, W41804, W9112, W22280, W9108, W9138, W9147, W28492, W22272, W9186, W9137, W41772, W28490, W9237, W28520, W22240, W41681, W9240, W41683, W9247, W9236, W41686, W22241, W9232, W9230, W9255, W41665, W28527, W9257, W22234, W9228, W9254, W28523, W41673, W9250, W9248, W9208, W28515, W9205, W41714, W9210, W9198, W41722, W22254, W22255, W22257, W28517, W41694, W9226, W9224, W9223, W41700, W41807, W22245, W22246, W9215, W9214, W22312, W41906, W9012, W41911, W9001, W9000, W28444, W28442, W9021, W41883, W9023, W9022, W41920, W9020, W9019, W9015, W9013, W22325, W8966, W8962, W8961, W28425, W8957, W8956, W8955, W22331, W8950, W8949, W41926, W9032, W8978, W8977, W41938, W41942, W41835, W9087, W28477, W28476, W28474, W9083, W9082, W28473, W9088, W28471, W9074, W9072, W28470, W9106, W9103, W22283, W9099, W9096, W9095, W41820, W9091, W41823, W28457, W9050, W41864, W41869, W9051, W9039, W9038, W9037, W9034, W9059, W9065, W9062, W9061, W22230, W28468, W9057, W28467, W9053, W9052, W9486, W9485, W28619, W28618, W9477, W9476, W22161, W41462, W9469, W9468, W9499, W22141, W28631, W28630, W9506, W22145, W9502, W22148, W22164, W22149, W28627, W41432, W28623, W41434, W41488, W9443, W9442, W41486, W28599, W9433, W9432, W9431, W28601, W9464, W22166, W28602, W9511, W9453, W9452, W22170, W9450, W41483, W9448, W22121, W9565, W28651, W9560, W9568, W41371, W28649, W22125, W41375, W9554, W28648, W9551, W22117, W9581, W22118, W22128, W9573, W9521, W9530, W9528, W28638, W9523, W9531, W22138, W22139, W22140, W22130, W41383, W28645, W9545, W9544, W9543, W9428, W9538, W9536, W9535, W41391, W9316, W41612, W41613, W9322, W9320, W9319, W9315, W9314, W9312, W9310, W9334, W9340, W28557, W22205, W28556, W9332, W28534, W9284, W9279, W9278, W41653, W41645, W9272, W9271, W28532, W9268, W22229, W28542, W28546, W22217, W9299, W9298, W9296, W22202, W41637, W9293, W9292, W9289, W9406, W41531, W9402, W41532, W28591, W9397, W9396, W41539, W41514, W9427, W9425, W41506, W9423, W9420, W9390, W28595, W9413, W22178, W28569, W41561, W41568, W9363, W9361, W28565, W9352, W22201, W9378, W41545, W41548, W9384, W28584, W9381, W9380, W9379, W10216, W9376, W9374, W29129, W11068, W21663, W39800, W11064, W11062, W11061, W11069, W21665, W11057, W11056, W29126, W11053, W39812, W11051, W11077, W11085, W11083, W11082, W39791, W21661, W11076, W11074, W11072, W11070, W11024, W11018, W39849, W21672, W11048, W21669, W11045, W11044, W39816, W21670, W29124, W11038, W11035, W11034, W21642, W11141, W11139, W39723, W29154, W21639, W29152, W21641, W11143, W11132, W29150, W11129, W11128, W11160, W11157, W11156, W11153, W11150, W11149, W39709, W39772, W21653, W11101, W11099, W39775, W11097, W11105, W21655, W39779, W29133, W11088, W11123, W21647, W11119, W11118, W29143, W11112, W21650, W39768, W29140, W39771, W11106, W39952, W29094, W10911, W10909, W21707, W10916, W10904, W10903, W39962, W39965, W10899, W29092, W10897, W10924, W39922, W39925, W10932, W10930, W10929, W39968, W10922, W29096, W39945, W21728, W10875, W39992, W29078, W10868, W10865, W29072, W10861, W40007, W29070, W29069, W21711, W21712, W10892, W21713, W10937, W39980, W10879, W39990, W10877, W39877, W10989, W10986, W10984, W10991, W10981, W21687, W10979, W10978, W10976, W10975, W39887, W11008, W11006, W39864, W11002, W10999, W10996, W21685, W10992, W21695, W10955, W10950, W10945, W10942, W10939, W29104, W10964, W39889, W21690, W10967, W10966, W10965, W11161, W21691, W10958, W10957, W11368, W11364, W39502, W39507, W11359, W11357, W11356, W11355, W11354, W21572, W11350, W11378, W21561, W11386, W21562, W39480, W21563, W11382, W21564, W11380, W29205, W21566, W39485, W11372, W39489, W29209, W21581, W11330, W21578, W29202, W39541, W11325, W11331, W29198, W11319, W29196, W11316, W21585, W39556, W11348, W39516, W21574, W11342, W39527, W39530, W11333, W39408, W11439, W29227, W11433, W39420, W11431, W11430, W39424, W11453, W11463, W11461, W11460, W11458, W39394, W11450, W11447, W21556, W11405, W39454, W39456, W29218, W39450, W39466, W29217, W21558, W11393, W21559, W29220, W11423, W11421, W29222, W29221, W11414, W11412, W11411, W11410, W39669, W21618, W11216, W21621, W39667, W39671, W39674, W11203, W11201, W21616, W11233, W39641, W11231, W11230, W39644, W11227, W11199, W39646, W11223, W11222, W11221, W11220, W39652, W21631, W11180, W11179, W11178, W11177, W11175, W11181, W11170, W11169, W11168, W11166, W39699, W11163, W11162, W11190, W11197, W21625, W39681, W11194, W39684, W11191, W29170, W29166, W11188, W39688, W21629, W11182, W11284, W21594, W21595, W21596, W11287, W11286, W11285, W39575, W29186, W39589, W39590, W29185, W29184, W11278, W11277, W11276, W11311, W29194, W39561, W21588, W39564, W29189, W11298, W29188, W21593, W21613, W11243, W11236, W21602, W11272, W39599, W11270, W11269, W39600, W11267, W40016, W29180, W11259, W40451, W40460, W10437, W10424, W10422, W21863, W28922, W10419, W21865, W10445, W10453, W10452, W10451, W10447, W10417, W10444, W10442, W28913, W40500, W28908, W28906, W28902, W10415, W28918, W40477, W10410, W10454, W28914, W10403, W10402, W10401, W10400, W40486, W10505, W10515, W40368, W21841, W40372, W10508, W40378, W21839, W10503, W21846, W21848, W21829, W21831, W28962, W10531, W40348, W10526, W10524, W21857, W10470, W10469, W10468, W40421, W28936, W10459, W10458, W10457, W10491, W10490, W40396, W40400, W10375, W10482, W21852, W10480, W40408, W10269, W40601, W10275, W10270, W40614, W10265, W21909, W10263, W28871, W40587, W10294, W10293, W28868, W10287, W10286, W10285, W10283, W10225, W10237, W40640, W10232, W10224, W10223, W10222, W40654, W40655, W21921, W10217, W10259, W10258, W10257, W10256, W10254, W10253, W10244, W10243, W10241, W10355, W10354, W10353, W40537, W21892, W40542, W10346, W10344, W10343, W10339, W10338, W10374, W10372, W10370, W10369, W21888, W10367, W10366, W10337, W10364, W21889, W10362, W10360, W10315, W40568, W40569, W21901, W10308, W10316, W40575, W10305, W40582, W10299, W40558, W10336, W10335, W10334, W10333, W10331, W10330, W10328, W40339, W10324, W10323, W10321, W28882, W10319, W21900, W10317, W10746, W10754, W40108, W10755, W40124, W10739, W10738, W40133, W10735, W40134, W10769, W10768, W21759, W40100, W10762, W10761, W10760, W29041, W40107, W29024, W40154, W10713, W10711, W10709, W10708, W10705, W29023, W10702, W10700, W40171, W10697, W10731, W40142, W10726, W29047, W29029, W10719, W10717, W10716, W10822, W10833, W10832, W40038, W29063, W10824, W10834, W40049, W10820, W10819, W10817, W10816, W40052, W21742, W10843, W21732, W10849, W40025, W29067, W40056, W10840, W21736, W10836, W10835, W10791, W21749, W21750, W10786, W10784, W40076, W10782, W10781, W21751, W21753, W40089, W21756, W10811, W29058, W40066, W40067, W10696, W40071, W10797, W21746, W40281, W10596, W40275, W40276, W10591, W21808, W21809, W28983, W10584, W10578, W10577, W40263, W10612, W10610, W21803, W28986, W28985, W21806, W40296, W40264, W21807, W10600, W10599, W10555, W40323, W21825, W40327, W10550, W28967, W40335, W21828, W10544, W10543, W40338, W10540, W10565, W21818, W40304, W10567, W28973, W10615, W28972, W10562, W40317, W10560, W28971, W21823, W10664, W10673, W40200, W10674, W40211, W10661, W10659, W40212, W10657, W40215, W21782, W29018, W10690, W21779, W29015, W21781, W10654, W40192, W29011, W10675, W10623, W28994, W10630, W10629, W10627, W10624, W10634, W10621, W28990, W10618, W10617, W10616, W10652, W10649, W21792, W40222, W28999, W10641, W10638, W40234, W40238, W19579, W33541, W19574, W19575, W19577, W31260, W33553, W19571, W17336, W31255, W33560, W33563, W33570, W19570, W17367, W17366, W17365, W17364, W31265, W33532, W19569, W33572, W17358, W17357, W17356, W33536, W33538, W17352, W19594, W33591, W17303, W31243, W33604, W17297, W17295, W33607, W17292, W33608, W19596, W19584, W17326, W17324, W33576, W17322, W33578, W31266, W33581, W33583, W31249, W31248, W17312, W31246, W17310, W33477, W17423, W17422, W33473, W17419, W17417, W33470, W19550, W19551, W33483, W17410, W17409, W31279, W31286, W17442, W19543, W17440, W31287, W19545, W17435, W31277, W17432, W31283, W33469, W17429, W17427, W17378, W33505, W19561, W17385, W17384, W19563, W33515, W17380, W19564, W33519, W33521, W17373, W17372, W33524, W19556, W31275, W33492, W17400, W17399, W17398, W17395, W19558, W17393, W17392, W33500, W33721, W17184, W17183, W17182, W17180, W31194, W17187, W19637, W17176, W19638, W17174, W17173, W17172, W33724, W17198, W17208, W17207, W19627, W31205, W17200, W17169, W17197, W17196, W31197, W17192, W17190, W17189, W33715, W19652, W33748, W19650, W33756, W33760, W19651, W17142, W19647, W19653, W33766, W33769, W19655, W33773, W31191, W17168, W19639, W17166, W17164, W19642, W33734, W17209, W17159, W31186, W33743, W17154, W17153, W31233, W17263, W17262, W33643, W19606, W31227, W17256, W33651, W33653, W31241, W17283, W17282, W17281, W19600, W19611, W17269, W17218, W17226, W33681, W19622, W17221, W33691, W17219, W17227, W33694, W17213, W17212, W33698, W19624, W17236, W31219, W17245, W17240, W33667, W19616, W17443, W17235, W19618, W17230, W33679, W19620, W17657, W33216, W33218, W33221, W17662, W33224, W17659, W33226, W19463, W19464, W33231, W19465, W19466, W33201, W33184, W33188, W17682, W31372, W19461, W33212, W33213, W33275, W31354, W17624, W17622, W17620, W17619, W31350, W17617, W31349, W19482, W17612, W17611, W17610, W17609, W33278, W19486, W17604, W17647, W17645, W17642, W33252, W31361, W19471, W17637, W17687, W19472, W17634, W17632, W33263, W19475, W33265, W17735, W33126, W19438, W19439, W17740, W17739, W33132, W17734, W17731, W17729, W31388, W19443, W33140, W17752, W17757, W19434, W17755, W19435, W17725, W31394, W17750, W17749, W33121, W17747, W17746, W31392, W33175, W17707, W17706, W17703, W33169, W19454, W31378, W19449, W17696, W17695, W33182, W33146, W33148, W17720, W33149, W17717, W31342, W17715, W33153, W31385, W19448, W33157, W17490, W31307, W33403, W33405, W33406, W31303, W19528, W33397, W17489, W33413, W17486, W17485, W33419, W19518, W17520, W17519, W33371, W31300, W33377, W31314, W33384, W33387, W17453, W33444, W31293, W17459, W19538, W17455, W17452, W33455, W31288, W17446, W19542, W17471, W19532, W19533, W17476, W33429, W33367, W17470, W33435, W19534, W33437, W33439, W19498, W17582, W17581, W31335, W33306, W33307, W17577, W19497, W33309, W17573, W19499, W31334, W17570, W33316, W17565, W17564, W33295, W33287, W19490, W33289, W33290, W17596, W33292, W17593, W33325, W33296, W17590, W17585, W33355, W19509, W17540, W33346, W33347, W31322, W33354, W17542, W17530, W17528, W19515, W17552, W17560, W33327, W17558, W31327, W33332, W33333, W19506, W17549, W17548, W17547, W17546, W16708, W34177, W16709, W34187, W34190, W34191, W16702, W16701, W34192, W16739, W19793, W34166, W16729, W16722, W16666, W19817, W16671, W16670, W16668, W19813, W16665, W19819, W19820, W16661, W34232, W16658, W16695, W34206, W16687, W31010, W16682, W16681, W34217, W16678, W16787, W19775, W19776, W19777, W19779, W16790, W34109, W16788, W16784, W34111, W16782, W34114, W16779, W34082, W31067, W34084, W16809, W19769, W31066, W31059, W16805, W31064, W16803, W31062, W19774, W34097, W34133, W16758, W16757, W16756, W16754, W34135, W16760, W16749, W31049, W34142, W34143, W16745, W16743, W34117, W31057, W16773, W16657, W16768, W16767, W34127, W19783, W16762, W16544, W16553, W34336, W34337, W34340, W34342, W30965, W16554, W16543, W30963, W34346, W16539, W16537, W34349, W19857, W30971, W19855, W16569, W34324, W34328, W16563, W16535, W16559, W16557, W16556, W34335, W34378, W34367, W16510, W16509, W16507, W30953, W19874, W16514, W16499, W16498, W19878, W16524, W16533, W16531, W34354, W30961, W30960, W19866, W19852, W16521, W16519, W34363, W16517, W34265, W16636, W16634, W19830, W34258, W19831, W16630, W34262, W19833, W31005, W16624, W16623, W16622, W34268, W34272, W19836, W34239, W16655, W16654, W34236, W16652, W34237, W16648, W16615, W16646, W19824, W19825, W19826, W16582, W16593, W16590, W16589, W30978, W19847, W16583, W16581, W34311, W30973, W16614, W30995, W34275, W19838, W16607, W16816, W19839, W16602, W17027, W33888, W17025, W17024, W17023, W33890, W33893, W17017, W19697, W33900, W33902, W17010, W19699, W33869, W17043, W19686, W17040, W17039, W19688, W17035, W19690, W33880, W19691, W31146, W16980, W19706, W16984, W16983, W16982, W16990, W16977, W16976, W16975, W16973, W16972, W16998, W31139, W33908, W19702, W17001, W16999, W19684, W16997, W31130, W19705, W16992, W17098, W19662, W17108, W19663, W17103, W19660, W17096, W33810, W33775, W17128, W17126, W31181, W33780, W33785, W33787, W33788, W33790, W17114, W31160, W17066, W33846, W17063, W33848, W17060, W17068, W33856, W33857, W17052, W33859, W17049, W33862, W19673, W33832, W33835, W33836, W19675, W17076, W33841, W17072, W17071, W16863, W19743, W16871, W31086, W16868, W34033, W16862, W19749, W19750, W34041, W16857, W16882, W16890, W16888, W31093, W34013, W16885, W16884, W16854, W31090, W16879, W16878, W16877, W16831, W16830, W19760, W31072, W16837, W16824, W19763, W16819, W34079, W16853, W34050, W16848, W16847, W16846, W16844, W16843, W16842, W31081, W19756, W31080, W19718, W16947, W16946, W19717, W16944, W33959, W16941, W31112, W16938, W16937, W19720, W16934, W31116, W16969, W31125, W31124, W16961, W33945, W19722, W16958, W19715, W16955, W31114, W33952, W19733, W31105, W33988, W16909, W16908, W33997, W16899, W16897, W16895, W34008, W16931, W16927, W19724, W16923, W31395, W16919, W16918, W19726, W18598, W18609, W32228, W19130, W32234, W32238, W32240, W18610, W19135, W19136, W19137, W32214, W32215, W18622, W18587, W18618, W32224, W18615, W18614, W31710, W18612, W32227, W18568, W18566, W32268, W19145, W18563, W18562, W18561, W18569, W19148, W32276, W32278, W32279, W19149, W18552, W19140, W18586, W32253, W18583, W19139, W18580, W18579, W32259, W32260, W31698, W31695, W32162, W18683, W18682, W18679, W32160, W31728, W18685, W31727, W32165, W32168, W18670, W18668, W18701, W18666, W18693, W18692, W18690, W18688, W32151, W32201, W32194, W32199, W19116, W18636, W32204, W31715, W32206, W32210, W18630, W32180, W18665, W18663, W31725, W19114, W18660, W18659, W32179, W18551, W32182, W18654, W18653, W32183, W19115, W32186, W32396, W19194, W18446, W31643, W18444, W18443, W32395, W18441, W19197, W19199, W32419, W18470, W32369, W18466, W32377, W19185, W31656, W32382, W18459, W19189, W18454, W31622, W18407, W18406, W31624, W32450, W18403, W18402, W18401, W18400, W32454, W19216, W18396, W32459, W19219, W32464, W18389, W32429, W32421, W31634, W19204, W18424, W18423, W18422, W32428, W32366, W32430, W31628, W19210, W19212, W32444, W32445, W31682, W18532, W31687, W31686, W32303, W18526, W31683, W18521, W32309, W19163, W18516, W18547, W32288, W18540, W31689, W18538, W18537, W32295, W18534, W18493, W32338, W32340, W32345, W32348, W18481, W18478, W19179, W19181, W32313, W32315, W32316, W32317, W19164, W19165, W32321, W18505, W31680, W18500, W31676, W32333, W18913, W31923, W18922, W18921, W18919, W18917, W31929, W31932, W19044, W18908, W31939, W18905, W31941, W18933, W31906, W31908, W18940, W18938, W18935, W18934, W18903, W31913, W19038, W31915, W18926, W19052, W31965, W19050, W31972, W18878, W31964, W18873, W18867, W18866, W31985, W31953, W18901, W31797, W31948, W18897, W31951, W19034, W18892, W18891, W18889, W18887, W31962, W18991, W18997, W31843, W18995, W31847, W18992, W19000, W18990, W31848, W18985, W19023, W19025, W31824, W19016, W19018, W19014, W31830, W31831, W19010, W18981, W31835, W19006, W31836, W19020, W18953, W18961, W18960, W31884, W18955, W31892, W31896, W19030, W18948, W19032, W18971, W18977, W31863, W31864, W18974, W18973, W31873, W31874, W18966, W31813, W31877, W31812, W18751, W18761, W32089, W18758, W32090, W32094, W32095, W18762, W18750, W18747, W19092, W19093, W18743, W18742, W18771, W18781, W18779, W19081, W32074, W19082, W31746, W19083, W32078, W32081, W32083, W31753, W32085, W19101, W32120, W18719, W18718, W19100, W32122, W18715, W32123, W18722, W32125, W32129, W19103, W32132, W18706, W19104, W18730, W18739, W31743, W31735, W18735, W32111, W18733, W32112, W19099, W18728, W32115, W18726, W32116, W32118, W18723, W19065, W32011, W32013, W18843, W18828, W18826, W31771, W32032, W32033, W18853, W18861, W18860, W31989, W18858, W18857, W32034, W31783, W31998, W18848, W18845, W19061, W18790, W18799, W18797, W18796, W32055, W19077, W18792, W18791, W32051, W18789, W18788, W32064, W19078, W18783, W18810, W18818, W18813, W32041, W32043, W18808, W18807, W18806, W18805, W32047, W32892, W17983, W17981, W17979, W17978, W17977, W17975, W19360, W32893, W19361, W17970, W17968, W31463, W17966, W31461, W17993, W18003, W19348, W19349, W17999, W31472, W17994, W17963, W17991, W17990, W32879, W19355, W32929, W17942, W17940, W32922, W32927, W32915, W19373, W17929, W32939, W17925, W17924, W17962, W17961, W32901, W17958, W17957, W17956, W19368, W32867, W17951, W17947, W32910, W32911, W17944, W18060, W18054, W32817, W19335, W32830, W18045, W18041, W18071, W18078, W32790, W32791, W19324, W18040, W31500, W18068, W32860, W31475, W18019, W19342, W18017, W32858, W18023, W19344, W19345, W19346, W19347, W32866, W31479, W18038, W18036, W31480, W32839, W18032, W19378, W18030, W31478, W18027, W32846, W19340, W18024, W17809, W17820, W17816, W33061, W17812, W17811, W33066, W17822, W17808, W33068, W33069, W17802, W33042, W17842, W31424, W19409, W17839, W17838, W33039, W19411, W33041, W17800, W33048, W17828, W17827, W33051, W17825, W17772, W17779, W17778, W19426, W19427, W33097, W33087, W17771, W33104, W17767, W19431, W33110, W17762, W17790, W33073, W17797, W17795, W31404, W33029, W17789, W17788, W33083, W31401, W17785, W31400, W17783, W17893, W17902, W19384, W17899, W17898, W17896, W31444, W17894, W32967, W19387, W31443, W32980, W19390, W17885, W19381, W31449, W17918, W32948, W19380, W32955, W17910, W32960, W17907, W17906, W32962, W19402, W17864, W17860, W33006, W17858, W31431, W17851, W33022, W19405, W33026, W31426, W17874, W31440, W17880, W31439, W17876, W17875, W19394, W32993, W19396, W18281, W32562, W19253, W31568, W18283, W18292, W32572, W32573, W19258, W19259, W32578, W32580, W32581, W18273, W32543, W18306, W32546, W31581, W18302, W31580, W18272, W19250, W18296, W18295, W32560, W18247, W18246, W18245, W31554, W19266, W18252, W32615, W18237, W18236, W31550, W32619, W32582, W32583, W32593, W18264, W18263, W19244, W32597, W32598, W18256, W32493, W32483, W18368, W31608, W18364, W18359, W18358, W18356, W32497, W19229, W18353, W32500, W18386, W32467, W32469, W32470, W18382, W31614, W32501, W18378, W31612, W18375, W18374, W18373, W19224, W32481, W18322, W18330, W31599, W18328, W32525, W18325, W32526, W32527, W32528, W31597, W18316, W18315, W32537, W32504, W18348, W32505, W19231, W32507, W19232, W32511, W19234, W18339, W19236, W18335, W18334, W19304, W31517, W19302, W32723, W18129, W32724, W18123, W32728, W18119, W18144, W18152, W18150, W18149, W32705, W19297, W18143, W18141, W19298, W19299, W31518, W19312, W18098, W18097, W19314, W19316, W32775, W19311, W32778, W18088, W19318, W31505, W32782, W18109, W32733, W31512, W32745, W32751, W18111, W32760, W32763, W18103, W18102, W32766, W19284, W18209, W18206, W31533, W19282, W32642, W18200, W32658, W32659, W31531, W32661, W32662, W32624, W32625, W18228, W18227, W18225, W19272, W32629, W32664, W19274, W18219, W18218, W19275, W32636, W19276, W18163, W18171, W18170, W18168, W31522, W18166, W18165, W32686, W18159, W32698, W18157, W19295, W18155, W19287, W18189, W18188, W18186, W32670, W32673, W32674, W16494, W18180, W18176, W18175, W32685, W20437, W20434, W14814, W14813, W35995, W20435, W35999, W20436, W30355, W14804, W14803, W14831, W30360, W14829, W20430, W14826, W14825, W35981, W30358, W35989, W30356, W14771, W14779, W14777, W20447, W20448, W14773, W20449, W20450, W14763, W20454, W36022, W14797, W20440, W20441, W30353, W14791, W36021, W14833, W30350, W14785, W30349, W14781, W30384, W30388, W14890, W35908, W35909, W14884, W14881, W14880, W30382, W14877, W14912, W14911, W14910, W35879, W14908, W35880, W35881, W20397, W35920, W35889, W30392, W20400, W14897, W14844, W14852, W35954, W14846, W14845, W20423, W30364, W30363, W14836, W14835, W30379, W20410, W14873, W14872, W20412, W14869, W14760, W14866, W35932, W35934, W30373, W20418, W14650, W14658, W30297, W36162, W14655, W14653, W30296, W36165, W14659, W14649, W20500, W14646, W36168, W20501, W36147, W14674, W14671, W36171, W14666, W14665, W14664, W20496, W14660, W14609, W36202, W14615, W14614, W36206, W14612, W14611, W30275, W14608, W30274, W14605, W30271, W20516, W14601, W36178, W14634, W36188, W36146, W30282, W30281, W30276, W14621, W36198, W36199, W20473, W30333, W36071, W14732, W14727, W36084, W14725, W30321, W36089, W20475, W36095, W14750, W14759, W20457, W14754, W14753, W30339, W14715, W14749, W14747, W14746, W30335, W36063, W14687, W30315, W30307, W14690, W30306, W14697, W14686, W36131, W20489, W30305, W20476, W36103, W20478, W20479, W30319, W14707, W14913, W30317, W14704, W36111, W20316, W35671, W15133, W15130, W15128, W30471, W15126, W15122, W35685, W20319, W15146, W15155, W30477, W20308, W35659, W15149, W35662, W20320, W15143, W15142, W15141, W15086, W15095, W15093, W35707, W15091, W15088, W20329, W15097, W15085, W35714, W15082, W20331, W15079, W15078, W15106, W35691, W15115, W15113, W15109, W35697, W15107, W15105, W20325, W15102, W15101, W15098, W35591, W15214, W15211, W20290, W15207, W15216, W15204, W15202, W15199, W20283, W15239, W20277, W35573, W15232, W15231, W15230, W20285, W35584, W15221, W20287, W15219, W30502, W35640, W15175, W15174, W35634, W35636, W30484, W15169, W15168, W15165, W20304, W15162, W15160, W15185, W15189, W15188, W30491, W15186, W30490, W30488, W15182, W15180, W35630, W20372, W20368, W35813, W14970, W14967, W30419, W20374, W20375, W20377, W35829, W14956, W14986, W14992, W20361, W35799, W35800, W14985, W30426, W14981, W14980, W14979, W35807, W20386, W35854, W14932, W14929, W14928, W14927, W35850, W14925, W35871, W14915, W20396, W20381, W14946, W14945, W14999, W30409, W30407, W35845, W35846, W14938, W30406, W30441, W35741, W15053, W15052, W15051, W15048, W15056, W20340, W15044, W20342, W15041, W35749, W20343, W35731, W20333, W15072, W15070, W35728, W15068, W15037, W35732, W30444, W15062, W15060, W15057, W20355, W15017, W15015, W35773, W35774, W35779, W15018, W35782, W15007, W15006, W15005, W15003, W15002, W15001, W15028, W15036, W20346, W30437, W35758, W30436, W20351, W15023, W35768, W14172, W30133, W14181, W36642, W36645, W36647, W20649, W20654, W30125, W20656, W30124, W20658, W36661, W14192, W14199, W36628, W14195, W36631, W14193, W20660, W36633, W14189, W36635, W36690, W20667, W14138, W14136, W14135, W14143, W14133, W14131, W36697, W20669, W14126, W36702, W20662, W36670, W14157, W36673, W36675, W14153, W36679, W36680, W30114, W14145, W36558, W36561, W20621, W14257, W14268, W14253, W30160, W14251, W30159, W36576, W20615, W14286, W20613, W14283, W14282, W36543, W14279, W30155, W14275, W30173, W14272, W14271, W14214, W36605, W14221, W36608, W20639, W20640, W14217, W14215, W36602, W14213, W14212, W20641, W14205, W14204, W20633, W36582, W30152, W14243, W14242, W30150, W36589, W14124, W14235, W36592, W36595, W36599, W14006, W14012, W14011, W36807, W20716, W36810, W14015, W36814, W14004, W30053, W14000, W20720, W13997, W36791, W14032, W14031, W14030, W30063, W14028, W14027, W14026, W30050, W36796, W20712, W14020, W14019, W20714, W13968, W13976, W13974, W30046, W13972, W36848, W36841, W13967, W13966, W13965, W36849, W36850, W13986, W13995, W13994, W36825, W20722, W13989, W13988, W30065, W13984, W13982, W13981, W13979, W20678, W30103, W14101, W14100, W14096, W14095, W14104, W36735, W36736, W36737, W36738, W14087, W30094, W14113, W36704, W14122, W30109, W14083, W14112, W14111, W36716, W20677, W14106, W36721, W20704, W14050, W14049, W20702, W14047, W36778, W20703, W36774, W14043, W20705, W30068, W14036, W36754, W14077, W14076, W14073, W14072, W14071, W14287, W36758, W36760, W14065, W14058, W14055, W14494, W14502, W14500, W14498, W20548, W14489, W14487, W36325, W14513, W14524, W14523, W14520, W14516, W30249, W14512, W14511, W14509, W14508, W36344, W20552, W30238, W36347, W14462, W36351, W14457, W36355, W20556, W36361, W14450, W14448, W36335, W14483, W36328, W14480, W36332, W20535, W36340, W36341, W14471, W14470, W14469, W30239, W14574, W20519, W14581, W14579, W14576, W14575, W36239, W20521, W14571, W36241, W20522, W14567, W14566, W14591, W14599, W14598, W36215, W36220, W36222, W36229, W36233, W36274, W14544, W36266, W14542, W30263, W20530, W20531, W14538, W14537, W36278, W36279, W30262, W36282, W14530, W36284, W30259, W36254, W14564, W14563, W14562, W36249, W14558, W14557, W36365, W14553, W36260, W14548, W36263, W36484, W14346, W36485, W30194, W36487, W36488, W14336, W36504, W36505, W14330, W14329, W14328, W36506, W14363, W14362, W36467, W36469, W14326, W20593, W20594, W30199, W14353, W14352, W14350, W30178, W14307, W14305, W14304, W36518, W20610, W14308, W36533, W14293, W14292, W36535, W36537, W14317, W14325, W14324, W14323, W14321, W14320, W14319, W36509, W14314, W14313, W36514, W14309, W30215, W14426, W30221, W14421, W14420, W36397, W14427, W14414, W14413, W20575, W20577, W20578, W36412, W14437, W30231, W30230, W36372, W14441, W20562, W20563, W36381, W14433, W14432, W14430, W30224, W14380, W36451, W20587, W36435, W14376, W30203, W14372, W14371, W14403, W14402, W36417, W14399, W15241, W30210, W36428, W20583, W16078, W16076, W16075, W16079, W34757, W16067, W16066, W34761, W34762, W16059, W16089, W16096, W34726, W34729, W34764, W16088, W16086, W30814, W16083, W30790, W20021, W16032, W20024, W16028, W16027, W34786, W16021, W16019, W16017, W16056, W16055, W16052, W34770, W16098, W16045, W30794, W16043, W34779, W34782, W16038, W16146, W16157, W16155, W16153, W16152, W19991, W16158, W30825, W34676, W19994, W16140, W34678, W34679, W16167, W16174, W16173, W16170, W16137, W16166, W16164, W16162, W16161, W34662, W16159, W16116, W20001, W16111, W34707, W16119, W34713, W16106, W34714, W16104, W30817, W16102, W34717, W16099, W30824, W16136, W34683, W34684, W34687, W19995, W34693, W16124, W19998, W19999, W34916, W34917, W15916, W15914, W15919, W20060, W15903, W30747, W20064, W20055, W15936, W15934, W34899, W15932, W30755, W15900, W15927, W34909, W34912, W15923, W20057, W15868, W20073, W15875, W20075, W15872, W20077, W34958, W34949, W34960, W15866, W15865, W15858, W15890, W34936, W15895, W15892, W34895, W34944, W15887, W15885, W15884, W20070, W34837, W30779, W15993, W15992, W34833, W30775, W34838, W34843, W20038, W15977, W34809, W16013, W16012, W30782, W34811, W34812, W16008, W16004, W16002, W20031, W30780, W15999, W30766, W34874, W34875, W15954, W34876, W30767, W34887, W15943, W20051, W30760, W15938, W15967, W15974, W34852, W15970, W30770, W34857, W15966, W34859, W20043, W34863, W15961, W30768, W34867, W16380, W16390, W16388, W16385, W16383, W19917, W19918, W16375, W30899, W34487, W16370, W34459, W16410, W16408, W16405, W16403, W34458, W34488, W16399, W34461, W16394, W30916, W19913, W16342, W16351, W34506, W16347, W16346, W34507, W16344, W16352, W16341, W34511, W19931, W16337, W19932, W16335, W16367, W16366, W19924, W16364, W19926, W30895, W16411, W19928, W16357, W16354, W16464, W16474, W34402, W16472, W19887, W16466, W16465, W16475, W16460, W19893, W16457, W16456, W16455, W30937, W30945, W34388, W16491, W16487, W30946, W16483, W16482, W19884, W19886, W34443, W30930, W19901, W34439, W34441, W16424, W16434, W16422, W16420, W34448, W34449, W16415, W16413, W30922, W16451, W16450, W34419, W16446, W16444, W16441, W34426, W16438, W16437, W34430, W16435, W16235, W16233, W34611, W19963, W16238, W19965, W16225, W16222, W34620, W16220, W34598, W34591, W34592, W16254, W16252, W16249, W16248, W30856, W30860, W16243, W16242, W34600, W16240, W16239, W16188, W16199, W16197, W16195, W19979, W19980, W30843, W16189, W16187, W34648, W16185, W16182, W16181, W16209, W16217, W30855, W34623, W34624, W19969, W30854, W16210, W30852, W16207, W19972, W16203, W19975, W30885, W34537, W16314, W16312, W16310, W16308, W16316, W16305, W16304, W16303, W16302, W16301, W34531, W30892, W16329, W34530, W16297, W34533, W16318, W30886, W34580, W34572, W16272, W34573, W34574, W19953, W30868, W19955, W30867, W34589, W16258, W34561, W30883, W16295, W34552, W34559, W16284, W30877, W34565, W30869, W35344, W15448, W15447, W15446, W15444, W15443, W15442, W30583, W30582, W15438, W15437, W15474, W20203, W15472, W35331, W15467, W35333, W15436, W15463, W15462, W30591, W15459, W15458, W20208, W20226, W35369, W20220, W35371, W35381, W30576, W15407, W15418, W15404, W15403, W15402, W20227, W35400, W15426, W30581, W20216, W35360, W15431, W20218, W15427, W30579, W35367, W30610, W20192, W35283, W35285, W15523, W15522, W15532, W35293, W15515, W15514, W15541, W30618, W35264, W15547, W30615, W35267, W20186, W35270, W15511, W30613, W15535, W30611, W30598, W15492, W35308, W15489, W30596, W15486, W15494, W15480, W15477, W15476, W35300, W35295, W30600, W15506, W35298, W35301, W15499, W15498, W15496, W15300, W15298, W15294, W35503, W20258, W35510, W35515, W15310, W15318, W15316, W35482, W15313, W15312, W15311, W15281, W15308, W35486, W15306, W15302, W30525, W30528, W20268, W35547, W20269, W35551, W20266, W15250, W15247, W35556, W35530, W15280, W20262, W35522, W15274, W35526, W35528, W35475, W15268, W35429, W35421, W35422, W15375, W15374, W35426, W15371, W15370, W15379, W35431, W20234, W35433, W15364, W15363, W15362, W15360, W15396, W15395, W15388, W35415, W15383, W20231, W35417, W35420, W15336, W15332, W20245, W15330, W35459, W15327, W15326, W15324, W15322, W20249, W15320, W35440, W15355, W15354, W15353, W30556, W30555, W20241, W35456, W35457, W15340, W30685, W35065, W15757, W35069, W15753, W35070, W15760, W20116, W35076, W30679, W15742, W15770, W30697, W15776, W20108, W35050, W35053, W20109, W20112, W15764, W15763, W15711, W15723, W35096, W35098, W20128, W15709, W15707, W20130, W15704, W15703, W15740, W35089, W35090, W15779, W15731, W15730, W35092, W15727, W34992, W15838, W15836, W30728, W15834, W15831, W15827, W15825, W15824, W30725, W15855, W20082, W34974, W15849, W15821, W15846, W30729, W15842, W15841, W15791, W30716, W30713, W15798, W35028, W15795, W15794, W35030, W15802, W15790, W30705, W15785, W20102, W30701, W35011, W15818, W20088, W15815, W15813, W15811, W35012, W30718, W20093, W15596, W30635, W35209, W15601, W20169, W15599, W15598, W35206, W35214, W30633, W35222, W15590, W15589, W15588, W15614, W35196, W15618, W35201, W15613, W35203, W15610, W15607, W15606, W35251, W35238, W35242, W30627, W35249, W35236, W30622, W15556, W35259, W20174, W15586, W30632, W15584, W20172, W15582, W15581, W30630, W15579, W15624, W35230, W20175, W35235, W15573, W30662, W15682, W15680, W35135, W30663, W15675, W20138, W35140, W35141, W35143, W30661, W35145, W20143, W15666, W35125, W35117, W15699, W15698, W20133, W20135, W15687, W15686, W35131, W35132, W35173, W15643, W35175, W35182, W15635, W20160, W35189, W15627, W15625, W15664, W35149, W15659, W15657, W35156, W15653, W20149, W3342, W3338, W47631, W3333, W3332, W3329, W3328, W3353, W3360, W26508, W47613, W24234, W3351, W26506, W3349, W3348, W3347, W3346, W3304, W3302, W3301, W3300, W3296, W26487, W3290, W3289, W3287, W3285, W24254, W3315, W26499, W3323, W3319, W3318, W3317, W24244, W3310, W3308, W24216, W26534, W3425, W3423, W3422, W3421, W3418, W3416, W3427, W3414, W47557, W47559, W47560, W3409, W3407, W47529, W26538, W3441, W3435, W3434, W3432, W3431, W3430, W3429, W3373, W3383, W3379, W24227, W3374, W3372, W24229, W3368, W3393, W26527, W3397, W3391, W3389, W3387, W26457, W3185, W3184, W3183, W26455, W24288, W3180, W24289, W24290, W3175, W26454, W24292, W3170, W3169, W24284, W26461, W47763, W3197, W3190, W47775, W3138, W3147, W24302, W3145, W3144, W3143, W3139, W3135, W3134, W3133, W26438, W3131, W3167, W26451, W26450, W47815, W3159, W3158, W3204, W47822, W3152, W24300, W3150, W3256, W3263, W3251, W3249, W3248, W3247, W3246, W24256, W3278, W24257, W26480, W3271, W3270, W3268, W3267, W3266, W24262, W3213, W24276, W24277, W3219, W3218, W3217, W24279, W3210, W24281, W47751, W26468, W26467, W3237, W3236, W3231, W3228, W3227, W3226, W3225, W3223, W3647, W3654, W3653, W3652, W3651, W26596, W26597, W3646, W3644, W3643, W3640, W3639, W3671, W24142, W3638, W3663, W3661, W3660, W3659, W47319, W3617, W3616, W3615, W24154, W3610, W3608, W26592, W3605, W47372, W24158, W47338, W3635, W3634, W3633, W3632, W3630, W24141, W24150, W3625, W3623, W3621, W47239, W3731, W24119, W24120, W24116, W3727, W3725, W3724, W26618, W3721, W24123, W24124, W26629, W3756, W3752, W24114, W3743, W3742, W3741, W3696, W26609, W47278, W24132, W47285, W3688, W26610, W3686, W3684, W47299, W3708, W3717, W3716, W3715, W3712, W24126, W3710, W3709, W3707, W47266, W3704, W26611, W3700, W3492, W26558, W24193, W24194, W3496, W24196, W3493, W24191, W3491, W3490, W3488, W24197, W3486, W3485, W24198, W26563, W3515, W3513, W3483, W24186, W24187, W3505, W24190, W3463, W24205, W3459, W47516, W3456, W3450, W26542, W3448, W3472, W3481, W26556, W3476, W26555, W24182, W26545, W3466, W3465, W3581, W3578, W3576, W3575, W3574, W26579, W3582, W3569, W3568, W26575, W3565, W24172, W47386, W3600, W26588, W26585, W3596, W3592, W3558, W3589, W3588, W26583, W3585, W24180, W26568, W3536, W3532, W3530, W3525, W47448, W3522, W3521, W3556, W24175, W3552, W24176, W3550, W3549, W3547, W3546, W3544, W3541, W2712, W2721, W2720, W2718, W2717, W26300, W2715, W2714, W26299, W24444, W2710, W48274, W2705, W26298, W24440, W24441, W2735, W24442, W2732, W2702, W48254, W48256, W2724, W2674, W2682, W2681, W2679, W2678, W2677, W26289, W2671, W26287, W2691, W2701, W26295, W48283, W2694, W2693, W24439, W2690, W2688, W24453, W24454, W2798, W2794, W24415, W2786, W26325, W2816, W26332, W2813, W48160, W2810, W48165, W2804, W2803, W2800, W24435, W2758, W2757, W2754, W2752, W2751, W2750, W2749, W26310, W24437, W2745, W2741, W2777, W24423, W24424, W2771, W2665, W2765, W26312, W26311, W2762, W2761, W26252, W2570, W2568, W26250, W2563, W24490, W2557, W2556, W2555, W2590, W26261, W24481, W24491, W2581, W26255, W26254, W26233, W2530, W2529, W2527, W24503, W24505, W2522, W2521, W48459, W2517, W24507, W26238, W2553, W2551, W2550, W26244, W24495, W2546, W2543, W26236, W2647, W2646, W2645, W2644, W26283, W2642, W26282, W2636, W24468, W48325, W26286, W2661, W24460, W26284, W2657, W48350, W2655, W2654, W2652, W2651, W2609, W2608, W2607, W26265, W2605, W2604, W2603, W2610, W2600, W26262, W2594, W2592, W2627, W2626, W2624, W2621, W26267, W3025, W24337, W3031, W26407, W3029, W3028, W3027, W3026, W24336, W3022, W3020, W47952, W26409, W3047, W24333, W24334, W3043, W47957, W3040, W3039, W26408, W3036, W3035, W2985, W26399, W26398, W26397, W2986, W24345, W2984, W2983, W2981, W2980, W24350, W3014, W3013, W26404, W3011, W3009, W3007, W24342, W24331, W3004, W3003, W3000, W2999, W2997, W3102, W26431, W3108, W3107, W3106, W3104, W24315, W24316, W47877, W3097, W26425, W26436, W24306, W3125, W3124, W3123, W3122, W24308, W3119, W3118, W3114, W3060, W3072, W3069, W3066, W3059, W26411, W3057, W3056, W3054, W3053, W3081, W47892, W3086, W3080, W3079, W26422, W3076, W3075, W2866, W2874, W26355, W2870, W2868, W2876, W2864, W26351, W24396, W2857, W2884, W2894, W48074, W24385, W2888, W24397, W48087, W26358, W2880, W24391, W2878, W48145, W26342, W24407, W2832, W26337, W2829, W24409, W26343, W2825, W48147, W48148, W2821, W2820, W2847, W2855, W24398, W2853, W26350, W2851, W24400, W2848, W26364, W2845, W2844, W2843, W2842, W2841, W2839, W26384, W2950, W2949, W2955, W2943, W2941, W2939, W2938, W2935, W2966, W2976, W2974, W26393, W26390, W2934, W2964, W2961, W2960, W24362, W2903, W2913, W2912, W24378, W2910, W2908, W48063, W26365, W2901, W2898, W24383, W2928, W2927, W2925, W24374, W26369, W47214, W2920, W24376, W24377, W4590, W4588, W4585, W23836, W4583, W26878, W23834, W4580, W4579, W23838, W4577, W4575, W4599, W4608, W4607, W4605, W4604, W4603, W4602, W4569, W26882, W46432, W23833, W4541, W26870, W46473, W4547, W4544, W4542, W4551, W46486, W4533, W23849, W4565, W4563, W4609, W4555, W4554, W4552, W4659, W4667, W23802, W4665, W26911, W26909, W4661, W4669, W26906, W26904, W4652, W23810, W4688, W4685, W4680, W46360, W46361, W4676, W4675, W4674, W4672, W4671, W23800, W4618, W4628, W4626, W4624, W26894, W4622, W4621, W46415, W4616, W26891, W23826, W46422, W4610, W23812, W26902, W4645, W4644, W23814, W4642, W23815, W4640, W4637, W4635, W4632, W23821, W46587, W4428, W4423, W4432, W46595, W4414, W4413, W4412, W4410, W4441, W4452, W26835, W23880, W4448, W4443, W4442, W4409, W4439, W23885, W46573, W4433, W4382, W4390, W26819, W23899, W4386, W4384, W4383, W4391, W4381, W4379, W4377, W23895, W46605, W46606, W4403, W23897, W4453, W46615, W4394, W4392, W4502, W46511, W4509, W26861, W26860, W4506, W4505, W4503, W26859, W4497, W26853, W4494, W4520, W4527, W23853, W4522, W26852, W26862, W4517, W4515, W4514, W4513, W4471, W4470, W4469, W23873, W26838, W4466, W4464, W4472, W4461, W4458, W23876, W23877, W4454, W4481, W4492, W26848, W46533, W26847, W4484, W4482, W4479, W4475, W4473, W46100, W23720, W23721, W46094, W4897, W26999, W23718, W4892, W46102, W23723, W4889, W46107, W23724, W4911, W27012, W4919, W27010, W46074, W4910, W27005, W27004, W46082, W23717, W4904, W4859, W26994, W26993, W4863, W23732, W4858, W23733, W26992, W4852, W4876, W4883, W23726, W4880, W4877, W46059, W4874, W4873, W4871, W4870, W23729, W45993, W4982, W27036, W4980, W23685, W4977, W27037, W23687, W27034, W23689, W45967, W5001, W45971, W4998, W27047, W4995, W4990, W4989, W4988, W4987, W45980, W4930, W4940, W27020, W4937, W4934, W4933, W27016, W23707, W23700, W4929, W4928, W46052, W4926, W27014, W27023, W23696, W4955, W23697, W23735, W4949, W46037, W4946, W4736, W4744, W4742, W4738, W23779, W4732, W4728, W26944, W4762, W4759, W26947, W23783, W4752, W4746, W4697, W4703, W4700, W4699, W4698, W4707, W46345, W4716, W4720, W4765, W26930, W4713, W26929, W46329, W26977, W4825, W23746, W4819, W26971, W26970, W4810, W4809, W4807, W4846, W23738, W4841, W4806, W4838, W4835, W4834, W4832, W26980, W4773, W4784, W23762, W46242, W4786, W26952, W4771, W4770, W46227, W46210, W46212, W23756, W46219, W26964, W4794, W4792, W46229, W4788, W24052, W3965, W47007, W3960, W24051, W26686, W3957, W24053, W3954, W3951, W3949, W3948, W26693, W26691, W3981, W3977, W46999, W24045, W26687, W3969, W3968, W3920, W3928, W3927, W3926, W3924, W26675, W24061, W24063, W3917, W3914, W3912, W24058, W3946, W3945, W3939, W24038, W3937, W3936, W3934, W3930, W4044, W4042, W46928, W24020, W46931, W24016, W4035, W4034, W4031, W26716, W4057, W4065, W24008, W24009, W46915, W26713, W4056, W4055, W24011, W24012, W24014, W4048, W3997, W26702, W46969, W4003, W24033, W46974, W3999, W26699, W26705, W24035, W3994, W3992, W26696, W3990, W3989, W4025, W4023, W46948, W4018, W24066, W4016, W46951, W4014, W4008, W24097, W47158, W3811, W3806, W3816, W3800, W3798, W3797, W3796, W3826, W3834, W24087, W3828, W3793, W26648, W3823, W24090, W3821, W26647, W24110, W3768, W24108, W26632, W3776, W3759, W26636, W3792, W24101, W3789, W3788, W24102, W3785, W3783, W47185, W24104, W3778, W3777, W3881, W3889, W3887, W3886, W3885, W24072, W3882, W3890, W26664, W3878, W3877, W3876, W3875, W24075, W3873, W26662, W3907, W24067, W26671, W47066, W47067, W3895, W47074, W3852, W3850, W24083, W3853, W3843, W26655, W47126, W3838, W24086, W3836, W3861, W3870, W24078, W3866, W3864, W3859, W3858, W3856, W24080, W26657, W23936, W23931, W4275, W23932, W26793, W26792, W23937, W4265, W23938, W23940, W23941, W4260, W4259, W4294, W26796, W4292, W4290, W4289, W4288, W4286, W26784, W4284, W4282, W23930, W4278, W4234, W4233, W4232, W4230, W4228, W4227, W4225, W4222, W26770, W4219, W26783, W46733, W4253, W26780, W46739, W23948, W4247, W26779, W26776, W23954, W4236, W23914, W46648, W4349, W4348, W4347, W26808, W4344, W4343, W23910, W4341, W4339, W46661, W26806, W4334, W4361, W4371, W4370, W4369, W4363, W26813, W4333, W23909, W4356, W4353, W4304, W4314, W4309, W23924, W4307, W4305, W4303, W4302, W4301, W4299, W4298, W26797, W4332, W4331, W46664, W4329, W4327, W4217, W26803, W23987, W4124, W4123, W4122, W4121, W26742, W26745, W26740, W4113, W4110, W23992, W26749, W4143, W46833, W4141, W46834, W4137, W23980, W4108, W23982, W26747, W4131, W26746, W4129, W4128, W46895, W4089, W26733, W4085, W23998, W26731, W4081, W46894, W4074, W4073, W4070, W4068, W4107, W4103, W4099, W26751, W46881, W4094, W4093, W4091, W4197, W4196, W4195, W4194, W4193, W4192, W4191, W23965, W4188, W26763, W4183, W23960, W4214, W26768, W23963, W26767, W46786, W4181, W4206, W4203, W4202, W4201, W4200, W4153, W4162, W4159, W4155, W26753, W46817, W4152, W4151, W4149, W4146, W23971, W26761, W4178, W4176, W4175, W4174, W4173, W4168, W46815, W4164, W837, W843, W839, W50148, W25625, W834, W25067, W829, W828, W25051, W869, W866, W865, W864, W862, W825, W25636, W858, W855, W25054, W851, W801, W25080, W799, W798, W796, W25084, W789, W788, W787, W816, W25069, W823, W25619, W25071, W25616, W819, W818, W25613, W808, W915, W923, W921, W919, W917, W25655, W925, W25036, W25648, W943, W941, W25028, W938, W936, W25031, W932, W930, W929, W886, W25047, W880, W50121, W25045, W50123, W876, W873, W896, W25645, W899, W784, W25042, W25642, W686, W25565, W683, W682, W25121, W25122, W676, W673, W696, W25571, W705, W701, W700, W699, W25114, W25126, W695, W690, W25135, W644, W641, W640, W638, W636, W25547, W25140, W658, W666, W25561, W25128, W660, W707, W25558, W25133, W650, W25581, W25582, W754, W50250, W747, W746, W745, W25601, W25600, W778, W25597, W773, W25594, W770, W25591, W766, W724, W722, W719, W715, W714, W713, W712, W25573, W710, W25103, W736, W946, W733, W732, W731, W25578, W729, W24957, W1152, W1150, W1143, W1142, W1177, W1175, W1171, W24949, W25746, W1163, W1161, W1116, W1113, W1112, W1111, W1110, W1109, W1117, W24967, W1105, W1103, W1101, W1138, W1135, W1132, W1178, W1127, W1124, W1123, W49894, W1118, W49774, W1236, W1224, W1223, W1222, W25769, W1219, W25773, W1255, W1253, W25777, W1247, W1244, W49756, W1241, W25771, W24928, W25755, W1194, W1190, W1188, W25764, W25753, W25752, W24944, W1181, W24946, W1206, W1217, W24931, W49796, W1204, W1202, W25765, W1199, W995, W1005, W998, W25690, W1006, W25009, W992, W991, W990, W989, W988, W1023, W24999, W1021, W1020, W25697, W25002, W1016, W25683, W1012, W1011, W1009, W25005, W1007, W955, W25022, W961, W960, W959, W958, W956, W965, W954, W953, W951, W950, W947, W984, W25012, W25675, W25015, W25016, W978, W1024, W25018, W25671, W971, W970, W967, W966, W1079, W1074, W1073, W1070, W24978, W1091, W1099, W1098, W1097, W24969, W24970, W24971, W1061, W1090, W1088, W25724, W1083, W1033, W24987, W1039, W1037, W25706, W1035, W24991, W24993, W25700, W25699, W24997, W24998, W1051, W1060, W24980, W25712, W1054, W1053, W25546, W24983, W49966, W24984, W1045, W24986, W25413, W221, W220, W25419, W217, W215, W222, W210, W208, W207, W206, W203, W200, W231, W240, W234, W233, W25407, W25422, W229, W227, W223, W168, W25280, W25401, W173, W25285, W169, W167, W165, W25289, W25393, W25291, W25392, W25406, W192, W25276, W187, W25278, W182, W291, W25450, W289, W25445, W25444, W283, W281, W25236, W319, W318, W317, W316, W315, W314, W312, W310, W309, W307, W306, W303, W260, W259, W258, W25436, W255, W262, W25254, W247, W246, W25257, W242, W270, W279, W278, W277, W275, W274, W273, W158, W269, W25440, W25248, W265, W263, W60, W25324, W57, W56, W55, W25325, W61, W45, W25370, W25316, W76, W75, W73, W25368, W25321, W10, W21, W25350, W15, W13, W5, W4, W3, W25343, W32, W40, W39, W37, W35, W80, W25330, W28, W25, W24, W25305, W135, W133, W131, W130, W128, W126, W124, W123, W122, W25306, W120, W117, W25298, W141, W89, W25312, W96, W95, W92, W90, W25376, W87, W85, W84, W25372, W81, W25309, W115, W112, W109, W108, W320, W25310, W524, W533, W532, W516, W515, W514, W25167, W552, W25527, W547, W545, W512, W25526, W539, W25169, W536, W484, W25183, W491, W487, W25184, W25506, W478, W25504, W25503, W25180, W510, W507, W505, W553, W500, W499, W25508, W495, W494, W25538, W610, W606, W605, W25540, W25148, W612, W25152, W597, W25153, W25143, W627, W626, W623, W622, W621, W619, W617, W616, W615, W614, W561, W569, W25162, W50445, W25529, W563, W560, W559, W25528, W25165, W555, W580, W25156, W586, W585, W583, W582, W581, W25159, W50437, W575, W574, W572, W368, W25218, W376, W372, W25217, W25222, W365, W364, W363, W362, W361, W396, W395, W393, W392, W25474, W390, W389, W388, W25223, W383, W382, W25216, W25233, W339, W338, W337, W335, W334, W340, W329, W324, W323, W350, W25470, W356, W355, W25469, W353, W347, W25465, W25464, W341, W447, W455, W454, W25194, W25195, W456, W444, W442, W440, W25495, W437, W464, W471, W468, W25499, W462, W461, W458, W457, W408, W25203, W416, W415, W25204, W25488, W412, W409, W25490, W407, W25485, W404, W25479, W435, W431, W430, W429, W428, W1257, W426, W25493, W419, W2093, W26101, W2100, W2098, W2096, W2095, W2102, W2092, W26092, W26091, W2110, W2117, W26103, W2115, W2114, W2113, W2082, W2106, W2105, W2104, W26083, W2056, W24651, W24652, W2051, W2049, W2043, W26080, W2073, W2081, W2079, W2078, W24638, W2076, W24640, W48913, W2067, W2164, W2169, W2168, W26111, W26109, W2161, W2159, W2155, W2191, W26115, W2189, W2185, W2184, W2154, W24615, W2179, W2177, W2174, W24627, W2132, W26106, W2127, W2126, W48877, W2123, W2122, W2121, W2145, W24625, W2151, W2149, W2041, W2144, W2141, W2139, W2138, W1932, W1943, W49055, W26042, W1944, W1930, W24690, W24692, W1924, W1923, W26055, W1961, W1960, W1958, W1957, W1953, W1951, W24681, W26044, W1945, W1889, W1897, W26020, W1895, W24707, W1899, W1888, W24709, W26014, W1880, W26027, W24693, W1919, W1918, W1916, W1914, W1913, W24697, W49029, W24701, W1906, W1903, W26023, W1900, W48969, W2016, W48976, W2011, W2008, W24665, W2006, W24666, W26069, W2003, W2002, W2001, W2031, W2040, W2037, W2036, W2035, W2000, W2026, W2025, W1973, W1982, W1981, W1979, W26063, W1976, W1974, W26064, W1972, W1971, W1967, W26060, W26068, W24669, W24611, W26067, W1988, W1986, W26065, W49007, W2408, W2406, W2404, W48567, W2397, W2395, W2394, W2390, W2417, W2426, W2425, W48553, W2423, W48557, W24538, W24539, W2416, W2415, W48563, W2413, W2410, W26173, W2370, W2359, W24555, W2357, W24557, W2379, W2388, W48602, W26177, W2377, W24551, W48614, W2373, W2372, W2371, W24516, W2489, W2488, W2487, W2486, W26213, W24518, W24519, W2478, W24520, W2475, W2503, W2514, W48469, W2506, W2471, W2497, W2495, W2436, W2445, W2443, W2442, W2439, W2437, W2435, W2434, W26193, W26192, W2459, W2470, W2461, W2352, W2457, W2448, W24599, W2248, W2246, W24597, W2242, W2240, W2249, W2236, W2235, W2234, W2232, W2231, W2269, W24592, W2261, W26135, W2257, W2250, W2204, W48788, W2213, W24610, W2221, W2226, W2225, W2223, W2222, W24603, W48775, W26124, W2215, W2214, W26160, W48670, W2325, W26158, W26152, W2316, W2315, W2312, W24574, W2342, W48645, W2344, W2338, W26167, W24564, W2332, W2278, W2290, W2288, W2287, W2284, W26143, W2280, W2276, W24587, W2273, W24588, W2308, W2307, W2306, W24577, W24578, W1879, W26147, W2295, W2293, W48708, W1465, W24851, W1460, W1457, W1455, W24854, W1453, W1452, W24855, W1449, W25861, W1484, W1483, W1478, W24844, W1446, W1474, W1472, W25853, W1469, W49538, W1418, W1427, W25839, W1425, W24866, W1417, W1416, W1415, W1437, W24858, W1439, W25864, W1435, W1430, W1429, W1535, W1540, W25879, W1537, W1536, W24824, W1529, W1527, W1555, W25890, W24817, W1560, W1559, W25889, W1553, W49448, W1548, W1547, W25881, W1502, W1500, W1499, W1498, W1496, W1492, W24840, W1487, W1523, W25878, W24828, W1409, W24831, W49495, W1311, W1310, W1307, W1306, W1304, W1301, W25790, W1322, W1330, W1329, W1327, W49678, W1325, W24897, W1323, W24898, W1318, W25801, W1316, W25798, W1266, W24913, W24914, W1272, W1271, W1269, W1267, W25787, W1264, W25783, W1260, W1259, W25789, W49715, W24906, W24907, W25802, W1285, W1284, W24908, W1282, W1280, W1278, W24876, W1382, W1381, W1380, W24881, W1389, W1377, W1372, W25815, W1399, W1404, W25830, W1397, W1396, W1395, W1393, W25824, W1340, W25809, W1348, W1347, W1345, W25807, W1342, W24889, W1339, W1338, W1336, W25804, W1333, W25814, W1364, W25813, W1360, W25892, W1357, W1356, W1355, W1353, W1352, W24746, W25971, W1772, W1770, W1769, W1777, W1767, W1765, W24748, W25970, W25969, W49237, W49209, W49199, W1794, W1759, W1787, W1784, W25974, W1779, W1778, W1740, W1738, W1733, W1731, W1741, W1729, W1727, W1724, W25956, W25955, W24753, W1757, W25968, W1753, W1752, W1751, W1745, W1850, W1857, W26005, W1851, W1859, W1849, W1848, W1842, W1878, W1876, W1875, W49116, W1872, W1871, W24713, W1841, W1868, W1864, W26008, W1808, W49174, W49175, W25987, W49178, W24732, W1811, W1810, W1809, W1807, W1806, W25986, W1803, W24734, W1800, W1829, W24721, W26002, W1837, W1833, W1828, W1824, W1823, W1819, W1818, W1621, W1619, W1618, W1617, W25910, W1622, W1612, W1609, W1608, W1602, W1601, W25903, W1639, W1638, W1636, W25915, W25913, W1632, W24795, W1628, W24796, W1624, W1623, W25893, W1580, W1577, W1571, W24813, W1569, W1568, W49426, W1566, W24814, W24808, W1598, W24804, W25901, W25899, W1642, W1589, W1585, W24810, W1701, W1700, W25949, W24766, W24767, W1693, W1703, W1691, W1690, W1688, W25947, W1717, W1716, W1713, W1682, W1711, W1708, W24762, W1706, W1664, W25937, W1662, W24778, W1659, W24779, W1652, W25925, W1645, W25920, W1673, W1681, W1680, W25945, W25942, W1677, W1675, W1674, W4451, W25941, W1671, W25940, W1667, W25938, W27846, W7343, W7342, W7341, W7340, W22893, W27848, W7333, W43568, W7327, W7352, W22886, W7363, W7362, W7361, W7359, W7326, W43547, W7349, W7348, W27850, W7305, W7303, W7302, W43593, W27831, W7306, W43605, W7293, W27827, W7316, W7324, W22898, W7320, W43575, W7318, W43536, W7314, W43580, W7312, W7307, W22869, W27868, W7416, W22867, W7413, W7411, W7420, W7408, W7407, W22870, W22871, W22872, W7402, W27869, W27872, W43462, W7435, W7434, W22859, W7432, W7431, W22861, W7401, W7427, W22863, W7421, W43523, W7382, W22880, W7379, W43513, W43517, W27856, W22885, W7370, W43532, W43535, W7366, W7287, W7385, W22879, W43504, W22878, W27861, W22875, W7392, W7393, W7394, W7397, W7400, W7185, W7192, W7189, W27803, W27800, W27799, W22937, W43679, W7212, W43682, W43683, W22928, W7207, W7205, W22938, W43691, W7201, W43692, W43694, W43695, W7197, W22951, W22947, W7157, W7153, W27792, W7147, W7146, W7141, W7140, W27795, W22939, W7171, W22940, W22941, W43678, W7166, W22945, W7162, W7161, W7160, W22915, W22912, W7266, W7264, W7262, W7261, W7270, W7259, W7257, W7256, W7255, W7254, W7253, W7286, W7285, W22908, W22909, W7277, W7276, W43622, W27826, W27824, W43668, W27812, W22925, W7227, W7226, W27811, W7223, W43669, W43672, W7217, W7215, W43460, W7232, W7234, W7236, W43658, W43657, W7239, W43654, W27815, W7244, W43646, W7250, W7638, W7645, W22784, W7640, W7639, W22785, W7635, W7634, W7633, W27967, W7665, W7663, W7662, W7661, W22777, W43262, W27962, W7652, W43244, W27959, W7648, W43305, W27938, W43301, W7598, W7606, W7595, W7594, W22802, W7591, W7589, W7619, W27956, W27954, W27953, W7621, W7620, W27944, W27942, W7611, W7608, W22757, W27996, W22753, W7720, W27994, W27992, W43173, W27987, W7710, W7708, W27983, W27982, W7731, W7740, W43147, W22748, W43153, W7736, W43155, W27998, W7728, W27997, W7724, W43223, W7686, W7682, W7679, W7678, W7675, W43224, W7671, W7588, W7689, W27977, W22764, W7695, W43203, W7700, W7702, W7482, W7490, W7489, W7486, W27891, W22846, W43411, W7481, W7479, W7478, W7477, W43420, W7508, W7506, W7505, W43395, W7502, W22842, W27893, W7498, W43402, W27892, W7494, W7492, W22857, W43437, W7454, W27880, W43440, W7443, W7442, W7440, W43459, W7458, W22853, W7461, W27885, W7465, W22850, W27889, W43423, W27890, W7559, W22807, W22809, W7563, W7570, W7557, W27927, W22817, W27924, W7550, W7578, W7584, W7583, W7580, W22805, W7576, W7575, W7572, W22806, W7519, W7529, W27911, W22831, W22832, W27908, W27905, W7521, W7515, W7514, W43387, W7531, W27915, W27919, W7535, W22825, W43361, W22820, W7546, W6725, W44187, W6719, W44192, W23100, W6727, W23101, W23102, W6711, W6710, W6709, W27623, W6737, W44158, W44161, W44162, W23092, W27622, W27638, W6732, W6731, W6729, W44181, W44247, W27607, W6679, W6678, W23120, W44255, W6669, W6666, W44263, W6696, W6695, W27615, W6689, W23116, W6687, W27611, W6801, W27655, W6797, W6795, W6794, W6791, W27652, W27650, W23067, W6821, W6817, W23071, W23073, W27648, W27656, W6806, W6805, W6804, W6756, W6765, W6764, W27643, W6760, W23088, W44150, W6753, W6752, W6750, W6749, W6748, W6769, W23084, W6772, W6773, W44131, W6779, W6780, W6782, W6784, W6563, W23153, W44358, W6569, W23154, W27584, W44364, W23152, W6560, W6559, W27579, W6557, W6554, W6589, W23147, W27589, W6582, W27578, W6578, W6577, W44352, W6573, W6534, W6533, W6532, W27574, W6530, W6529, W44388, W23168, W6521, W44393, W27564, W44397, W23171, W6544, W6551, W44375, W6549, W6548, W23161, W23144, W6543, W6542, W6541, W6539, W6538, W6537, W6636, W6644, W44289, W6642, W6638, W6637, W6646, W6635, W6634, W6633, W6632, W6630, W6661, W23125, W23126, W23127, W23128, W6628, W6653, W6652, W23129, W6649, W6647, W6608, W44326, W6604, W6603, W6602, W6601, W27596, W23141, W6594, W6592, W44337, W6614, W6615, W6616, W23133, W6618, W6622, W6623, W44307, W44305, W6626, W43864, W7037, W7033, W7031, W7029, W43848, W7023, W7020, W7018, W7057, W7056, W27754, W7052, W7049, W43843, W7041, W7040, W23008, W6990, W6998, W6987, W6986, W23010, W23011, W7012, W7009, W23003, W43885, W43889, W7002, W27740, W7105, W7113, W7112, W7111, W7109, W7106, W7114, W7103, W7100, W22969, W27765, W7125, W7136, W43756, W7133, W43759, W7129, W7096, W27771, W7120, W7119, W22964, W7067, W22981, W7075, W7074, W27757, W7072, W7069, W22985, W7065, W22986, W7062, W23013, W22978, W7081, W43808, W7083, W7084, W22977, W22975, W7090, W27761, W44029, W6880, W44031, W6877, W6875, W6874, W44035, W23049, W23050, W6867, W44018, W23043, W27695, W6895, W27694, W6892, W23046, W6865, W6888, W6887, W6847, W27683, W6845, W27678, W6842, W6840, W6838, W6848, W6836, W23065, W6899, W23055, W6850, W6851, W6853, W6855, W6857, W27686, W6863, W44041, W27717, W6947, W6946, W43967, W6941, W6939, W27709, W6936, W6965, W6978, W27733, W6974, W6971, W6970, W6969, W43937, W43942, W6959, W27699, W23036, W6910, W6908, W6917, W6904, W6901, W7742, W6918, W6919, W6923, W6924, W43986, W23033, W23032, W27706, W6934, W28255, W22477, W8538, W8536, W8534, W8533, W22481, W8540, W28254, W42364, W8525, W8524, W8523, W8522, W8556, W8554, W8551, W8550, W8549, W8521, W42344, W8546, W8545, W8544, W8493, W8501, W22490, W42385, W8498, W22489, W8491, W8490, W8487, W8486, W8485, W28253, W8519, W8518, W8515, W8514, W8513, W22472, W42372, W8510, W28251, W22456, W8613, W8612, W22453, W8609, W8603, W8602, W8601, W8599, W28270, W8597, W8625, W8631, W22446, W8628, W42267, W8626, W8596, W42274, W22450, W8618, W22451, W8615, W8567, W8576, W8573, W8571, W42324, W8568, W8579, W8566, W42334, W8560, W22471, W8580, W8581, W8582, W8583, W8585, W22464, W22463, W8589, W28268, W42299, W22459, W22458, W42499, W42510, W8386, W8385, W8381, W8379, W22523, W42522, W8403, W8412, W8409, W8407, W8406, W8405, W8375, W8402, W22517, W22518, W8396, W8356, W8355, W8354, W8353, W22530, W8351, W22529, W8347, W8345, W42552, W8343, W8341, W8340, W22524, W8372, W8371, W8368, W22526, W22513, W42534, W8363, W8362, W42536, W22527, W8358, W42423, W8462, W42421, W8459, W8456, W8455, W42430, W42432, W8483, W8480, W8479, W8477, W28239, W8449, W8473, W22495, W8470, W8469, W8468, W8421, W8428, W8427, W8426, W22510, W22511, W8423, W22509, W22508, W8434, W8435, W8439, W22506, W8441, W28231, W22503, W8838, W8845, W8842, W42074, W8839, W8850, W8837, W28373, W8858, W22366, W28387, W8864, W22369, W8859, W8857, W22370, W42056, W42058, W8808, W8803, W42107, W28360, W42109, W8809, W8797, W28359, W8794, W8793, W28358, W42092, W8827, W8826, W8824, W8822, W8821, W28369, W8819, W8817, W28368, W42099, W8811, W28406, W28411, W28408, W8922, W8920, W41988, W8918, W8917, W8915, W8914, W8913, W8911, W22353, W22338, W22354, W28417, W8932, W28412, W8878, W8885, W8884, W22359, W8887, W8877, W22360, W42032, W28392, W8870, W22365, W8888, W42019, W8890, W8892, W8895, W8898, W42003, W28399, W28307, W8689, W8688, W8687, W8686, W42221, W8681, W8691, W8678, W28305, W28302, W8670, W8699, W42200, W22422, W8706, W8705, W28313, W8702, W8701, W8669, W8698, W8693, W8692, W22443, W22440, W42252, W8645, W28281, W28286, W8640, W28279, W8637, W8636, W8652, W8653, W8654, W8655, W22437, W8658, W8662, W8663, W8665, W8766, W8765, W28335, W8763, W8761, W8760, W42144, W8767, W42145, W42146, W8755, W8752, W28331, W22388, W42122, W8787, W22390, W8784, W8783, W28328, W28345, W8776, W8771, W28336, W22402, W22419, W8728, W8726, W22415, W42187, W8721, W22418, W8718, W8717, W8715, W8714, W8713, W8339, W8731, W22411, W22410, W8736, W8737, W8739, W8746, W8747, W28327, W22679, W7941, W22680, W7939, W7938, W42955, W28058, W7943, W42964, W7930, W7929, W7927, W42967, W7925, W7951, W7960, W7958, W28065, W42946, W7950, W7949, W7948, W7947, W28063, W7945, W7897, W22691, W7902, W7901, W28049, W7899, W22694, W42989, W7895, W22696, W7893, W7891, W22687, W42972, W22686, W7921, W7920, W7919, W7918, W7917, W7962, W7914, W28052, W28050, W8018, W8017, W22651, W8013, W8012, W42872, W28082, W22663, W28089, W28090, W22645, W8033, W22647, W42864, W7996, W8026, W8024, W28088, W8021, W8020, W7971, W7977, W28072, W28071, W42926, W42927, W7967, W22673, W7889, W22668, W7982, W22667, W7988, W22666, W28073, W28076, W7993, W7994, W7995, W43093, W7793, W22732, W7790, W28018, W7787, W28016, W43104, W7783, W28012, W22726, W7814, W7813, W43081, W22727, W7802, W7800, W7751, W43135, W7756, W43137, W7753, W28003, W22744, W7749, W22745, W7745, W7743, W7818, W43129, W7767, W7769, W7770, W22738, W7773, W7774, W7775, W28011, W7777, W7779, W7863, W28044, W28041, W7868, W28038, W22704, W7865, W22705, W7861, W7860, W28037, W7857, W43002, W43003, W7886, W7885, W7883, W7855, W7877, W7875, W22700, W7837, W22715, W43055, W22717, W22718, W7823, W7822, W7821, W22721, W7819, W8036, W28033, W22711, W43035, W22708, W7849, W43030, W7852, W28036, W28175, W8245, W42655, W8240, W8238, W22568, W8233, W8232, W8230, W28183, W22557, W8259, W8257, W8228, W8253, W22561, W28180, W8250, W22563, W8199, W28172, W8207, W8206, W8204, W28168, W22574, W8196, W28166, W8191, W8218, W22569, W42670, W8225, W22570, W42673, W8222, W42674, W22571, W8264, W8217, W22573, W8215, W8213, W8212, W8211, W8312, W22540, W42575, W8316, W8315, W8313, W8321, W22541, W8309, W42585, W8329, W8337, W8334, W8333, W28211, W8302, W28209, W8326, W8325, W8324, W8323, W42631, W42616, W8284, W8283, W8280, W42614, W8273, W8270, W8269, W8268, W42633, W8287, W28194, W42609, W8291, W42605, W28199, W28200, W42599, W8297, W22546, W28203, W8093, W8090, W8088, W8087, W42796, W8085, W8094, W8083, W8080, W8077, W8103, W8111, W8110, W42782, W8107, W28125, W28124, W8104, W8102, W8101, W8100, W22617, W8097, W8095, W28096, W28106, W28104, W8051, W8050, W28100, W22631, W8043, W42846, W8040, W28092, W28091, W42824, W28107, W22629, W8062, W42816, W8067, W22627, W22626, W8162, W8167, W22591, W8164, W8172, W8161, W8159, W42733, W28156, W8156, W8155, W28153, W22583, W28164, W22585, W42708, W8182, W22596, W22587, W42723, W8175, W8174, W8173, W42769, W42752, W28145, W28142, W8132, W8129, W8128, W8136, W8121, W42770, W42773, W8117, W8115, W28148, W8138, W22600, W8140, W8144, W8146, W28152, W22597, W8150, W42738, W8152, W6129, W6125, W45569, W6127, W5733, W5484, W6128, W27227, W6130, W5732, W23425, W5226, W44794, W5422, W45443, W5365, W45445, W6117, W5891, W6119, W27438, W23427, W23291, W23511, W5231, W5734, W27129, W23431, W45566, W27230, W44789, W5370, W6140, W23603, W5217, W27232, W6143, W23288, W6145, W6135, W27312, W23289, W5724, W44790, W27179, W6115, W23373, W23599, W5722, W27125, W27310, W45720, W6138, W6139, W6090, W44844, W5469, W44842, W6089, W23515, W5805, W6091, W5741, W6094, W5247, W6073, W44852, W5900, W5744, W6077, W6080, W5249, W27222, W45033, W6082, W27431, W44820, W45699, W5893, W23296, W45570, W5473, W27372, W23295, W6105, W6112, W23595, W45449, W45704, W5737, W5246, W27433, W6097, W23300, W5739, W5489, W27435, W27178, W6102, W23297, W5240, W27305, W45121, W23274, W5182, W27457, W27458, W5184, W27303, W5876, W6196, W27452, W44753, W6183, W27115, W44751, W6185, W6186, W5705, W5875, W5187, W5703, W6190, W6211, W5873, W6207, W5692, W23621, W44714, W45412, W27107, W23441, W6212, W5690, W5168, W27469, W6214, W23624, W27466, W5698, W23270, W23400, W5696, W44718, W5381, W45119, W5501, W27122, W5811, W23606, W23433, W6150, W6155, W23286, W5200, W6157, W6158, W5882, W5371, W5213, W5212, W6146, W6147, W45124, W27368, W5715, W6148, W23604, W23280, W5377, W5495, W23282, W23281, W44765, W27119, W45761, W5193, W5707, W5706, W27446, W6178, W27447, W23610, W27367, W6161, W5881, W6162, W6163, W6165, W6166, W44775, W23435, W5197, W5376, W5710, W23607, W5442, W5970, W23344, W27395, W27396, W27397, W27382, W5975, W5976, W27399, W5351, W27394, W23339, W5979, W27211, W5785, W27340, W23338, W5319, W5324, W5802, W5323, W5321, W5320, W5782, W23363, W5317, W5919, W5966, W45008, W5777, W5993, W27332, W23555, W5353, W5992, W5303, W6000, W5301, W5428, W5449, W5308, W5981, W5915, W5982, W5984, W5985, W23336, W23570, W27393, W5988, W5989, W5990, W5445, W5991, W5307, W5446, W45594, W23354, W23559, W5343, W23353, W5342, W5943, W5341, W44998, W23405, W5339, W5947, W5434, W5435, W5796, W27346, W5927, W5801, W5929, W44996, W5349, W23358, W5933, W44993, W23357, W5346, W5432, W23356, W5798, W27389, W5939, W5441, W5958, W5923, W5330, W5791, W5328, W27383, W5789, W5788, W5325, W23348, W5949, W44976, W27391, W5952, W5334, W23407, W6001, W27206, W23351, W27208, W23361, W23350, W5905, W5360, W6052, W6054, W5275, W5274, W6055, W45161, W23551, W27219, W5462, W5904, W6047, W23519, W27417, W23418, W6046, W23552, W5280, W23317, W45467, W44882, W6050, W5278, W27139, W23587, W45674, W5750, W5749, W5258, W27138, W5254, W5253, W23309, W5748, W5747, W5746, W5901, W45025, W5269, W5267, W6059, W6061, W6062, W27422, W5264, W27140, W23371, W27221, W5295, W5770, W5452, W45641, W5768, W5358, W23328, W23575, W23326, W23324, W5292, W5767, W6018, W6005, W5356, W23332, W23553, W23415, W5771, W23524, W6008, W27153, W23574, W27415, W44902, W6034, W45470, W27326, W45500, W5760, W23369, W23320, W44895, W27218, W44907, W5766, W23323, W23368, W23322, W5289, W44908, W5288, W6025, W23623, W6027, W5765, W6030, W44904, W44903, W6402, W5603, W5052, W6400, W27253, W5844, W5051, W44516, W27279, W6403, W5843, W5050, W23660, W23485, W27528, W5845, W5540, W5541, W5825, W6391, W6392, W5047, W5413, W6394, W6395, W6396, W23205, W5542, W5547, W6423, W5546, W5043, W5041, W6425, W27062, W45314, W5841, W5038, W6428, W5840, W27274, W5400, W5037, W6408, W6410, W45532, W23202, W23201, W27067, W27534, W6418, W45299, W6366, W5620, W23213, W5072, W5071, W44548, W6370, W44542, W27283, W5617, W5068, W44540, W27524, W23492, W23491, W5074, W23217, W45890, W6357, W5823, W45086, W5530, W6375, W5393, W6360, W6361, W27285, W6362, W6363, W5824, W23215, W6387, W5063, W5062, W5847, W5061, W5060, W6385, W27281, W6386, W27185, W23463, W23490, W5609, W27252, W27525, W27527, W23210, W5534, W6378, W5615, W6380, W23544, W5414, W5613, W27359, W6383, W44529, W6487, W5831, W6483, W27049, W27258, W27551, W6492, W27266, W23174, W6470, W6471, W5584, W45328, W6473, W5582, W5016, W6475, W6477, W27189, W5580, W45948, W44406, W5571, W5827, W5007, W5006, W5569, W44403, W6513, W27354, W5566, W6502, W6495, W45336, W44415, W44414, W6469, W5409, W5574, W6503, W6504, W5010, W6505, W6506, W27558, W5553, W44478, W23193, W45322, W5839, W5590, W44473, W5550, W27538, W6447, W27539, W6450, W5031, W27256, W23189, W6434, W23196, W5596, W5401, W45919, W44487, W6432, W23541, W44467, W6435, W6436, W45367, W6438, W5549, W5593, W5592, W23183, W6464, W5558, W23479, W5586, W44456, W27051, W5834, W5585, W23181, W5833, W5836, W5030, W45929, W27541, W5403, W6455, W6456, W27542, W23399, W27056, W6463, W5405, W27297, W44656, W5386, W23637, W5664, W6262, W6263, W44660, W23247, W27496, W45232, W6267, W27296, W44667, W6218, W45249, W27096, W5868, W5666, W5816, W5134, W23380, W5665, W23241, W6280, W5867, W6282, W23240, W5866, W45837, W5660, W5131, W27242, W23639, W45832, W6219, W5872, W5657, W5127, W23242, W5126, W23627, W6230, W6231, W5680, W27476, W45813, W5150, W5149, W45234, W23261, W6224, W5161, W5382, W27302, W5159, W44702, W45236, W5156, W27474, W45411, W27475, W5155, W27101, W5676, W5144, W27299, W45245, W23258, W27481, W5142, W6245, W5509, W27471, W5140, W5385, W23256, W5672, W23633, W27483, W23634, W23628, W23629, W6235, W5146, W27478, W23381, W5145, W44687, W44686, W5384, W27480, W6241, W5392, W6329, W27084, W5091, W5090, W5522, W23225, W23226, W23650, W45083, W6337, W5689, W27516, W5096, W5639, W5095, W44588, W45544, W6324, W27353, W5854, W5637, W6325, W5636, W27288, W44587, W27085, W6327, W27364, W5081, W6350, W45879, W23219, W5626, W5077, W45288, W44560, W27521, W6354, W6355, W44570, W5087, W6342, W5097, W5085, W6345, W5525, W45286, W5628, W5113, W23237, W5112, W6299, W23499, W5651, W6303, W5111, W5108, W6286, W5864, W45265, W5116, W5115, W6292, W6293, W6297, W27184, W27088, W5642, W5102, W5641, W6315, W45858, W5643, W27087, W5099, W6319, W5688, W23383, W23497, W45855, W6309, W6310, W27290, W5859, W5646, W5105, W27510, W5519, W6314, W31492, W28693, W29708, W28193, W27200, W31490, W26840, W25635, W31499, W25633, W26841, W28696, W28698, W25637, W28751, W25713, W31417, W28136, W31414, W26810, W31408, W29675, W27243, W28141, W27244, W25720, W25725, W28755, W30110, W28746, W30089, W30090, W31430, W26816, W25709, W30095, W26815, W26814, W31425, W30099, W31423, W26811, W25711, W28748, W28103, W30118, W27257, W28771, W29659, W25738, W28777, W25741, W28778, W29658, W30115, W25744, W28101, W28779, W29656, W28099, W25750, W31383, W30127, W30129, W28763, W28758, W29666, W30112, W28760, W28761, W27251, W28762, W25705, W25728, W25731, W25732, W25733, W28115, W25736, W26801, W26827, W28177, W31466, W25657, W31465, W29697, W26829, W28176, W30054, W25661, W27216, W27217, W31462, W25663, W28719, W25667, W26823, W26822, W28174, W26832, W27202, W30047, W26836, W28705, W31474, W27203, W28706, W28707, W28708, W26834, W28726, W28713, W31473, W28715, W25650, W26831, W31471, W31470, W25656, W29700, W25693, W28162, W30069, W30071, W27233, W30078, W31441, W29684, W27234, W25696, W30082, W28159, W29680, W26817, W28158, W27239, W31434, W30061, W25669, W26821, W27223, W31454, W28702, W31451, W26820, W25681, W27226, W25684, W27228, W25687, W31448, W27092, W26990, W28322, W26991, W28329, W28505, W27090, W25432, W28498, W31739, W28496, W25427, W27094, W28513, W29808, W28318, W31730, W26983, W25447, W28510, W28509, W29921, W28508, W29809, W28507, W26987, W25410, W25414, W27086, W28487, W29912, W25411, W28491, W28485, W28484, W31761, W29823, W31763, W27089, W29915, W31751, W25423, W25421, W28348, W31754, W28351, W25416, W27108, W31703, W31704, W25472, W25471, W28293, W26959, W31708, W28294, W31711, W25487, W28545, W29943, W25484, W25478, W26960, W31700, W28540, W26954, W28536, W25460, W26973, W28314, W28518, W28315, W26975, W29922, W27102, W26978, W25457, W27098, W26962, W29804, W29934, W28306, W27103, W28308, W31764, W25467, W28522, W26967, W29932, W31719, W25463, W31721, W25367, W28397, W25369, W27033, W31811, W29855, W27054, W28405, W27035, W27052, W29875, W28440, W27026, W31803, W29845, W29883, W31805, W28453, W27024, W27060, W27059, W28451, W27027, W29846, W25371, W28426, W28428, W25354, W25353, W25351, W31822, W27048, W27041, W25347, W25346, W28423, W31815, W28435, W25362, W27038, W28433, W29873, W31801, W31819, W28431, W25358, W29893, W29899, W28370, W28371, W25390, W27007, W31779, W25387, W31784, W27078, W28472, W27077, W25404, W28366, W25402, W29904, W29902, W28367, W31769, W25400, W25386, W31773, W31775, W28479, W31796, W29836, W27019, W29887, W27021, W27070, W28459, W27068, W28389, W28454, W29832, W31789, W28375, W25379, W29891, W31792, W27075, W27072, W29890, W25568, W26879, W30016, W30012, W28227, W31555, W27167, W28646, W27166, W31562, W31566, W27165, W25562, W25572, W31536, W31537, W25574, W31544, W27171, W25570, W25569, W28225, W30020, W28629, W29756, W25550, W25548, W27157, W26898, W28628, W31592, W25545, W31594, W28626, W28641, W31567, W27161, W28232, W28633, W25553, W30001, W28632, W31578, W25607, W27182, W28212, W25611, W26863, W31509, W25605, W26864, W26866, W28214, W28676, W27180, W27188, W25631, W28205, W25630, W26849, W25628, W29718, W25627, W31504, W25599, W25621, W28684, W29721, W28682, W29722, W28659, W27176, W29733, W28662, W31526, W31528, W31525, W28219, W28656, W28221, W25575, W28674, W26868, W25595, W28675, W25587, W25586, W29730, W31520, W25584, W28673, W28672, W28668, W27177, W31661, W28266, W27127, W25507, W31659, W25505, W31668, W28579, W28267, W26931, W28587, W26921, W28262, W31649, W27132, W31652, W28263, W28588, W29783, W28586, W27130, W25510, W28264, W29958, W26941, W29945, W28275, W29796, W26945, W28547, W27124, W31673, W28576, W31674, W28572, W28571, W27135, W29954, W29953, W28560, W28559, W28271, W25498, W25532, W28605, W29865, W26903, W28242, W29762, W28243, W25530, W29981, W31611, W27141, W28616, W28622, W27152, W28620, W25541, W26901, W28617, W28614, W25537, W25536, W27150, W29984, W29959, W31630, W26916, W25519, W29776, W31632, W31629, W31633, W25516, W25514, W27136, W25513, W31636, W26913, W29765, W28600, W31618, W29769, W26844, W28598, W28258, W26914, W31627, W28260, W25524, W27137, W30861, W27749, W26196, W30864, W29428, W27750, W26194, W30445, W26197, W29432, W26562, W27753, W30443, W30870, W27745, W27467, W27744, W29426, W26209, W30859, W29145, W30872, W26205, W26203, W26202, W27746, W29141, W27747, W26201, W27766, W30435, W27764, W29125, W29441, W30433, W29442, W29440, W29123, W29122, W26174, W29445, W26570, W26571, W27769, W26565, W30878, W29132, W30439, W27756, W29424, W27758, W27445, W27759, W27444, W26567, W26185, W26248, W27722, W27725, W27726, W29164, W27728, W27730, W26235, W27702, W27493, W26529, W26532, W30479, W26257, W30819, W27482, W26535, W30475, W29404, W26549, W29419, W26225, W26224, W27470, W30845, W26222, W30847, W26550, W29155, W26217, W30455, W30453, W29417, W30830, W27734, W30464, W29163, W27735, W26230, W29161, W30432, W26229, W27736, W27473, W30835, W29473, W27814, W27429, W29474, W27428, W27817, W27427, W27820, W29084, W30397, W26595, W26132, W29101, W30947, W27434, W29099, W27810, W30396, W29464, W29095, W30955, W30376, W26600, W30974, W30975, W26602, W26604, W29483, W30980, W27421, W26605, W26606, W29066, W27418, W30370, W30993, W27426, W27821, W26114, W29077, W30943, W30970, W29074, W29482, W26108, W27823, W30917, W26577, W29117, W27783, W30427, W29116, W26156, W26155, W27784, W27786, W30918, W30425, W27787, W30919, W29447, W27770, W26572, W30431, W27775, W26170, W27788, W26168, W26165, W29118, W26136, W26141, W26138, W26590, W27437, W26137, W30939, W27801, W30941, W26134, W30423, W26582, W30924, W30420, W26146, W27798, W30412, W30569, W29258, W26371, W30670, W30673, W26367, W26366, W27605, W29246, W30683, W30669, W29267, W30580, W26385, W29265, W27537, W30665, W26380, W27529, W29261, W26377, W30578, W26376, W29259, W26375, W27631, W30707, W27621, W30709, W29358, W27625, W29239, W30710, W27627, W27619, W30560, W30559, W29237, W26347, W29236, W30719, W26346, W29356, W26363, W29245, W30690, W30692, W29244, W27608, W30564, W26469, W29240, W27617, W27582, W29303, W30626, W26414, W26410, W27554, W29321, W27553, W27581, W26415, W29326, W29296, W29294, W30594, W29328, W27586, W27549, W26428, W29311, W30612, W27565, W26406, W29314, W27569, W30616, W26430, W27575, W26420, W26416, W27544, W27592, W30590, W29274, W30649, W30652, W26449, W26453, W27598, W30659, W26396, W27540, W29337, W27601, W27548, W30593, W29287, W30636, W29286, W30592, W26403, W29280, W26446, W30639, W29276, W26447, W26402, W26401, W29335, W29275, W27681, W27508, W30516, W26509, W27685, W26510, W30509, W30506, W30781, W30505, W26511, W26503, W27668, W27670, W29203, W30769, W27674, W29389, W29378, W30526, W30522, W27676, W26294, W29201, W30773, W26522, W26273, W26524, W30808, W30810, W26526, W30803, W30487, W29393, W29172, W26264, W27701, W26263, W26520, W30785, W26514, W30498, W30787, W30495, W30789, W30791, W29181, W30492, W30801, W29179, W27641, W29363, W30733, W27642, W26485, W30736, W26324, W30737, W30739, W30549, W30740, W26495, W27637, W27635, W27636, W26473, W29230, W29372, W29359, W26483, W27640, W27523, W26328, W30534, W26498, W29208, W29207, W30533, W29375, W26501, W26302, W30761, W27661, W26301, W27664, W30765, W30544, W26317, W30743, W27647, W26497, W29216, W26309, W26305, W30540, W26303, W27519, W29210, W31254, W26729, W25874, W27316, W31252, W30216, W25871, W28878, W31250, W28015, W31258, W31259, W26732, W30214, W25880, W30229, W27325, W29595, W31242, W26725, W27322, W30225, W28006, W29603, W28007, W30222, W28010, W27320, W27318, W25876, W30207, W28860, W28859, W25845, W28858, W27308, W26739, W31274, W28028, W30202, W25840, W28855, W28865, W31263, W27314, W25862, W28023, W25852, W31269, W28024, W25848, W30244, W31204, W29572, W31207, W31208, W25909, W27972, W26707, W26708, W25904, W27338, W30253, W25926, W25917, W27968, W28910, W28907, W26701, W31235, W31225, W28887, W26719, W28886, W28885, W26721, W27999, W28883, W31237, W25882, W28000, W26722, W28002, W27329, W29578, W29579, W28892, W31210, W29582, W26715, W27989, W31212, W28890, W31216, W29590, W26777, W31343, W26775, W31345, W25778, W30147, W31348, W25775, W30146, W30145, W31351, W31353, W30140, W31356, W31331, W30166, W25788, W29644, W25786, W28810, W30149, W31369, W25767, W30135, W31371, W28794, W25763, W29654, W27264, W25751, W30131, W31379, W30137, W26781, W31362, W30138, W28077, W29642, W28081, W28084, W25768, W27271, W25823, W26752, W25821, W25819, W28839, W30188, W30187, W29617, W26754, W28836, W28835, W25811, W26757, W28833, W25810, W30201, W25836, W28853, W28851, W25833, W30197, W30195, W28842, W25827, W30174, W29633, W29637, W30176, W27287, W31324, W29639, W28061, W25797, W30172, W28817, W31328, W31330, W26769, W29628, W31308, W31310, W31311, W27293, W31312, W30180, W31316, W25803, W31317, W28824, W27292, W28051, W29016, W31061, W27867, W30331, W30330, W30327, W29511, W29010, W30325, W30322, W26054, W26634, W26072, W31051, W26071, W26633, W31056, W31068, W30341, W29507, W30338, W30336, W31084, W26644, W26645, W26032, W30316, W28998, W28996, W26031, W26030, W27883, W26028, W30308, W26025, W28993, W31088, W28991, W27387, W31073, W27400, W26642, W26043, W29003, W29002, W26035, W27840, W26614, W29057, W26616, W31007, W29054, W26100, W30361, W31009, W27414, W27829, W30365, W26607, W29064, W27828, W30996, W29061, W26088, W26612, W31004, W29059, W27404, W31031, W27406, W29037, W29036, W31042, W26079, W30348, W29498, W29032, W27857, W26077, W27859, W26087, W31014, W26621, W31016, W31021, W31022, W26082, W26626, W27854, W28931, W25957, W28929, W31163, W27357, W27356, W28928, W26679, W27943, W31167, W25953, W27947, W27949, W31170, W31154, W28952, W28950, W26674, W29546, W28947, W25967, W28946, W27355, W28942, W27361, W27360, W25962, W31157, W28941, W25958, W29552, W31184, W31182, W28923, W26690, W30260, W27960, W28919, W26694, W27350, W25935, W26695, W25933, W25931, W30258, W30255, W28915, W29559, W31172, W31173, W25950, W30268, W30267, W25948, W27955, W31177, W31179, W29560, W27352, W31180, W28925, W28980, W27894, W31110, W27895, W27897, W31111, W26659, W28975, W26001, W25999, W26665, W30294, W27906, W30303, W26016, W31096, W26015, W31098, W26011, W31103, W31104, W27379, W30298, W26010, W27374, W25972, W25982, W25979, W28958, W27929, W25977, W29544, W26669, W28957, W31140, W31141, W27934, W31142, W28954, W31118, W25994, W29655, W27920, W30277, W27921, W26666, W27923, W44619, W44594, W44567, W44703, W44699, W44697, W44689, W44666, W44665, W44662, W44469, W44457, W44501, W44497, W44926, W44942, W44940, W44922, W44911, W44988, W44995, W44990, W44989, W44884, W44949, W44947, W44774, W44766, W44814, W44760, W44755, W44748, W44742, W44863, W44821, W43981, W44007, W43999, W43982, W44015, W43957, W44088, W44086, W44083, W44071, W44053, W44034, W43818, W43845, W43838, W43832, W43825, W43819, W43815, W43813, W43798, W43932, W43930, W43928, W43926, W44091, W43884, W43862, W44336, W44312, W44231, W44391, W44386, W44383, W44166, W44163, W44143, W44141, W44135, W44096, W44092, W44225, W44214, W44185, W44182, W45822, W45821, W45792, W45788, W45779, W45907, W45902, W45861, W45853, W45836, W45656, W45639, W45625, W45718, W45715, W46135, W46124, W46110, W46079, W46078, W46218, W46213, W46164, W45988, W45984, W45977, W45951, W45920, W46053, W45206, W45171, W45302, W45296, W45281, W45278, W45262, W45254, W45089, W45078, W45102, W45049, W45149, W45141, W45135, W45125, W45114, W45108, W45504, W45490, W45488, W45469, W45468, W45456, W45590, W45587, W45585, W45580, W45571, W45543, W45529, W45371, W45365, W45364, W45437, W45409, W45387, W45383, W42259, W42254, W42242, W42239, W42236, W42233, W42228, W42307, W42345, W42317, W42306, W42302, W42300, W42296, W42288, W42139, W42108, W42104, W42220, W42218, W42203, W42175, W42172, W42171, W42164, W42578, W42573, W42541, W42660, W42653, W42640, W42630, W42380, W42414, W42382, W42361, W42360, W42358, W42352, W42351, W42520, W42515, W42490, W42477, W42450, W42439, W41720, W41718, W41712, W41704, W41699, W41690, W41680, W41678, W41675, W41671, W41670, W41666, W41664, W41778, W41775, W41774, W41763, W41762, W41757, W41754, W41661, W41744, W41734, W41732, W41589, W41587, W41582, W41577, W41576, W41543, W41656, W41650, W41648, W41609, W41607, W41973, W41994, W41992, W41981, W41978, W41974, W41997, W41955, W42064, W42049, W42033, W42030, W42029, W41877, W41842, W41880, W41829, W41825, W41819, W41805, W41945, W41939, W41930, W41905, W41900, W41889, W43377, W43414, W43404, W43398, W43380, W43373, W43465, W43453, W43439, W43276, W43288, W43236, W43232, W43353, W43319, W43732, W43710, W43684, W43681, W43786, W43766, W43765, W43652, W43757, W43755, W43750, W43557, W43556, W43555, W43542, W43538, W43511, W43492, W43618, W43645, W43643, W43637, W43635, W43631, W43630, W42838, W42857, W42823, W42822, W42893, W42928, W42922, W42908, W42901, W42900, W42891, W42890, W42881, W42739, W42731, W42717, W42707, W42699, W42805, W42797, W42791, W42790, W42786, W42778, W42754, W43142, W43122, W43119, W43103, W43100, W43186, W43216, W43208, W43205, W43075, W43176, W42979, W42983, W42981, W42976, W42958, W43054, W43051, W43025, W43022, W43017, W49437, W49433, W49527, W49276, W49379, W49368, W49341, W49687, W49816, W49570, W49668, W49660, W49634, W48848, W48836, W48803, W48790, W48777, W48936, W48915, W48908, W48899, W48669, W48664, W48739, W48717, W48706, W48695, W49087, W49086, W49234, W49190, W48963, W48958, W49068, W49839, W50563, W50539, W50072, W50059, W49893, W50116, W50242, W50225, W50198, W46966, W47004, W46987, W46985, W46826, W46812, W46811, W46793, W46888, W46886, W46848, W47274, W47260, W47226, W47369, W47041, W47180, W47162, W46425, W46517, W46475, W46299, W46241, W46239, W46378, W46372, W46369, W46335, W46325, W46714, W46707, W46764, W46753, W46748, W46734, W46732, W46729, W46561, W46555, W46544, W46531, W46621, W46641, W46638, W46635, W46624, W46589, W48183, W48234, W48226, W48022, W47993, W48114, W48106, W48073, W48577, W48540, W48537, W48322, W48396, W48395, W47584, W47565, W47539, W47531, W47665, W47649, W47626, W47611, W47414, W47404, W47375, W47514, W47510, W47458, W47919, W47897, W47860, W47854, W47933, W47689, W47824, W47768, W34941, W34963, W34957, W34956, W34952, W34948, W34947, W34939, W34937, W34932, W34921, W35042, W35041, W35035, W35033, W35019, W35016, W34999, W34968, W34810, W34807, W34801, W34794, W34789, W34784, W34768, W34767, W34752, W34743, W34892, W34890, W34885, W34883, W34878, W34865, W34850, W34848, W34844, W34841, W34834, W34828, W34822, W35204, W35247, W35243, W35234, W35228, W35225, W35224, W35215, W35199, W35198, W35194, W35185, W35177, W35312, W35282, W35281, W35174, W35276, W35265, W35260, W35255, W35077, W35105, W35101, W35100, W35088, W35087, W35084, W35114, W35074, W35063, W35059, W35054, W35144, W35172, W35166, W35160, W35158, W35155, W35146, W35139, W35138, W35134, W35133, W35130, W35129, W34366, W34392, W34387, W34384, W34379, W34376, W34372, W34362, W34356, W34355, W34343, W34339, W34450, W34447, W34417, W34330, W34412, W34410, W34408, W34404, W34400, W34395, W34261, W34260, W34257, W34255, W34254, W34248, W34238, W34264, W34230, W34219, W34211, W34207, W34205, W34302, W34326, W34322, W34320, W34317, W34309, W34303, W34288, W34273, W34622, W34646, W34642, W34640, W34632, W34626, W34625, W34647, W34612, W34596, W34594, W34593, W34674, W34702, W34696, W34694, W34692, W34688, W34672, W34667, W34657, W34653, W34650, W34649, W34501, W34493, W34484, W34482, W34481, W34479, W34471, W34466, W34457, W34553, W34583, W34578, W34569, W34567, W34564, W34562, W34560, W34557, W35330, W34549, W34543, W34540, W34534, W34526, W34524, W36079, W36073, W36070, W36067, W36065, W36092, W36061, W36047, W36164, W36161, W36157, W36149, W36143, W36139, W36133, W36042, W36121, W36106, W36104, W35929, W35958, W35956, W35950, W35946, W35963, W35925, W35923, W35921, W35912, W35903, W36004, W36040, W36037, W36031, W36023, W36017, W36016, W36002, W35993, W35976, W35972, W35968, W36403, W36399, W36396, W36405, W36342, W36329, W36480, W36474, W36470, W36463, W36460, W36456, W36453, W36327, W36433, W36418, W36413, W36411, W36252, W36248, W36247, W36240, W36235, W36226, W36211, W36210, W36201, W36255, W36196, W36194, W36187, W36186, W36180, W36294, W36309, W36302, W36299, W36267, W36264, W35534, W35565, W35564, W35563, W35539, W35566, W35529, W35509, W35508, W35596, W35638, W35631, W35629, W35627, W35624, W35601, W35597, W35585, W35580, W35359, W35391, W35388, W35386, W35373, W35362, W35354, W35348, W35335, W35453, W35469, W35468, W35466, W35465, W35449, W35443, W35432, W35803, W35824, W35823, W35822, W35815, W35814, W35809, W35826, W35802, W35797, W35781, W35771, W35893, W35875, W35869, W35867, W35769, W35862, W35853, W35848, W35844, W35840, W35839, W35827, W35703, W35701, W35694, W35692, W35690, W35686, W35683, W35706, W35672, W35670, W35664, W35655, W35646, W35645, W35763, W35761, W35759, W35755, W35754, W35751, W35747, W35745, W35733, W35729, W35719, W35710, W32637, W32667, W32665, W32660, W32656, W32653, W32648, W32641, W32640, W32669, W32635, W32633, W32621, W32618, W32617, W32616, W32719, W32769, W32768, W32753, W32731, W32725, W32722, W32720, W32708, W32695, W32694, W32689, W32688, W32530, W32512, W32495, W32532, W32480, W32479, W32473, W32463, W32461, W32458, W32455, W32604, W32599, W32595, W32585, W32575, W32570, W32568, W32566, W32565, W32772, W32533, W32976, W32972, W32970, W32961, W32949, W32947, W32943, W32942, W32933, W32923, W32909, W32907, W32904, W32903, W32902, W32899, W33038, W33036, W33030, W33018, W33016, W33005, W32997, W32992, W32837, W32824, W32819, W32815, W32810, W32808, W32806, W32842, W32794, W32789, W32784, W32783, W32781, W32780, W32779, W32774, W32897, W32889, W32888, W32885, W32883, W32878, W32875, W32453, W32864, W32863, W32862, W32861, W32859, W32854, W32097, W32087, W32077, W32075, W32071, W32069, W32101, W32066, W32053, W32052, W32040, W32036, W32028, W32177, W32164, W32131, W32114, W32109, W32106, W32104, W31927, W31925, W31917, W31914, W31912, W31910, W31901, W31899, W31934, W31881, W31872, W31855, W31842, W31834, W31984, W32015, W31995, W31987, W32188, W31982, W31981, W31978, W31976, W31963, W31959, W31938, W32390, W32386, W32383, W32379, W32374, W32367, W32364, W32363, W32397, W32351, W32347, W32344, W32343, W32334, W32330, W32423, W32448, W32443, W32440, W32436, W32434, W32426, W32425, W32424, W32324, W32422, W32416, W32402, W32400, W32399, W32254, W32250, W32248, W32242, W32236, W32235, W32232, W32258, W32230, W32216, W32213, W32211, W32205, W32291, W32320, W32318, W32306, W32305, W32299, W32293, W32292, W33049, W32290, W32289, W32285, W32270, W32269, W32265, W32263, W33819, W33864, W33855, W33853, W33843, W33839, W33837, W33834, W33826, W33821, W33811, W33925, W33921, W33916, W33903, W33887, W33714, W33704, W33702, W33701, W33699, W33695, W33685, W33671, W33669, W33781, W33774, W33764, W33761, W33755, W33754, W33934, W33742, W33741, W33728, W33726, W33722, W34120, W34106, W34100, W34099, W34094, W34092, W34128, W34088, W34083, W34075, W34066, W34167, W34195, W34194, W34186, W34183, W34179, W34170, W34168, W34165, W34144, W34136, W34129, W33967, W34000, W33994, W33992, W33983, W34004, W33966, W33961, W33958, W33944, W33942, W33938, W33936, W34035, W34053, W34048, W34047, W34040, W34037, W34032, W34030, W34024, W34014, W33262, W33281, W33280, W33276, W33274, W33273, W33272, W33271, W33268, W33264, W33256, W33254, W33242, W33238, W33311, W33348, W33338, W33323, W33314, W33312, W33308, W33301, W33300, W33299, W33291, W33288, W33086, W33122, W33117, W33105, W33101, W33093, W33128, W33085, W33078, W33077, W33070, W33064, W33060, W33055, W33161, W33211, W33205, W33200, W33186, W33174, W33172, W33159, W33154, W33147, W33137, W33133, W33575, W33574, W33558, W33557, W33551, W33547, W33577, W33535, W33527, W33525, W33518, W33613, W33645, W33644, W33635, W33624, W33623, W33619, W33612, W33609, W33584, W33399, W33425, W33424, W33422, W33411, W33409, W33407, W33401, W33394, W33389, W33379, W33375, W33373, W33369, W33365, W33364, W33499, W33498, W33497, W33488, W33486, W33485, W33466, W33463, W33461, W33457, W33448, W33447, W39790, W39785, W39778, W39764, W39762, W39736, W39728, W39725, W39714, W39871, W39840, W39807, W39611, W39605, W39618, W39587, W39574, W39572, W39566, W39693, W39691, W39686, W39680, W39880, W39661, W39660, W39636, W39625, W40080, W40079, W40078, W40048, W40047, W40045, W40039, W40032, W40160, W40194, W40190, W40180, W40179, W40174, W40167, W40158, W40156, W40148, W39958, W39944, W39936, W39971, W39921, W39895, W39893, W40026, W40009, W40008, W40000, W39988, W39978, W39974, W39973, W39138, W39137, W39129, W39154, W39114, W39101, W39099, W39098, W39193, W39216, W39208, W39202, W39196, W39089, W39181, W39176, W39171, W38979, W39025, W39024, W39021, W39015, W39013, W39009, W38995, W38992, W38982, W38962, W38952, W38951, W39065, W39088, W39086, W39059, W39055, W39050, W39042, W39034, W39465, W39459, W39432, W39479, W39415, W39406, W39403, W39379, W39555, W39550, W39547, W39528, W39514, W39505, W39491, W39484, W39257, W39289, W39288, W39267, W39264, W39260, W39256, W39242, W39241, W39235, W39233, W39354, W39352, W39344, W39341, W39328, W39304, W41128, W41071, W41035, W41031, W41198, W41176, W41173, W41165, W41142, W40927, W40911, W40905, W40904, W40889, W40885, W40866, W40860, W40848, W40992, W41018, W41009, W41002, W40986, W40970, W40952, W40951, W40945, W41410, W41403, W41400, W41397, W41393, W41523, W41512, W41497, W41387, W41475, W41473, W41469, W41463, W41454, W41453, W41265, W41298, W41282, W41276, W41270, W41252, W41245, W41236, W41234, W41233, W41229, W41342, W41382, W41380, W41374, W41363, W40412, W40386, W40377, W40371, W40484, W40519, W40516, W40514, W40513, W40479, W40478, W40470, W40461, W40266, W40257, W40256, W40249, W40225, W40216, W40196, W40336, W40326, W40324, W40322, W40319, W40315, W40308, W40303, W40292, W40291, W40285, W40764, W40758, W40776, W40737, W40839, W40830, W40800, W40797, W40787, W40783, W40608, W40604, W40577, W40565, W40616, W40532, W40526, W40687, W40686, W40680, W40675, W40673, W38939, W40646, W40639, W40630, W37321, W37364, W37362, W37341, W37324, W37323, W37313, W37280, W37266, W37455, W37453, W37448, W37440, W37425, W37405, W37404, W37392, W37388, W37373, W37151, W37174, W37165, W37164, W37162, W37158, W37140, W37112, W37220, W37263, W37257, W37256, W37253, W37200, W37197, W37190, W37183, W37628, W37680, W37679, W37657, W37651, W37621, W37611, W37610, W37713, W37744, W37738, W37737, W37726, W37723, W37715, W37588, W37712, W37706, W37703, W37702, W37698, W37694, W37518, W37515, W37514, W37506, W37499, W37524, W37483, W37469, W37466, W37465, W37464, W37586, W37585, W37567, W37553, W37106, W37551, W37543, W37542, W37541, W37540, W37527, W36664, W36666, W36665, W36710, W36659, W36654, W36652, W36650, W36648, W36640, W36764, W36749, W36746, W36745, W36733, W36726, W36723, W36717, W36556, W36539, W36572, W36524, W36502, W36501, W36499, W36598, W36634, W36630, W36617, W36770, W36596, W36593, W36587, W36586, W36580, W36579, W36577, W37008, W37037, W37025, W37023, W37022, W37019, W37017, W37016, W37003, W37000, W36995, W36989, W36988, W37071, W37099, W37094, W37073, W37056, W36824, W36819, W36806, W36804, W36797, W36832, W36790, W36788, W36780, W36779, W36773, W36772, W36959, W36931, W37745, W36886, W36884, W36872, W36858, W36846, W38593, W38590, W38566, W38563, W38560, W38598, W38556, W38631, W38681, W38680, W38675, W38670, W38640, W38622, W38613, W38608, W38601, W38424, W38418, W38416, W38412, W38389, W38384, W38381, W38377, W38356, W38519, W38506, W38491, W38479, W38464, W38455, W38454, W38449, W38446, W38435, W38842, W38867, W38855, W38851, W38845, W38844, W38869, W38824, W38821, W38816, W38809, W38923, W38921, W38915, W38912, W38908, W38907, W38807, W38893, W38887, W38879, W38878, W38872, W38708, W38735, W38724, W38717, W38744, W38707, W38703, W38702, W38698, W38695, W38770, W38805, W38785, W38782, W38776, W38772, W38353, W38761, W38754, W38752, W38751, W38748, W37973, W37969, W37968, W37967, W37966, W37964, W37961, W37958, W37952, W37939, W37938, W37937, W37917, W38037, W38034, W38033, W38022, W38015, W38006, W38004, W38002, W37977, W37822, W37821, W37810, W37803, W37798, W37779, W37773, W37770, W37762, W37866, W37904, W37896, W37889, W37878, W37869, W38043, W37856, W37844, W37840, W37836, W38239, W38282, W38276, W38271, W38264, W38253, W38288, W38230, W38226, W38223, W38220, W38219, W38213, W38352, W38351, W38349, W38346, W38341, W38340, W38333, W38209, W38320, W38298, W38297, W38102, W38091, W38089, W38088, W38087, W38084, W38082, W38078, W38075, W38067, W38061, W38050, W38046, W38172, W38187, W38186, W38185, W38184, W38181, W38171, W38168, W38161, W1, W38141, W4512, W4500, W4501, W4504, W8145, W8143, W4511, W18875, W13185, W13180, W18872, W4516, W18865, W8139, W8137, W8153, W4487, W4489, W13171, W18896, W4491, W18893, W4493, W4525, W13173, W4496, W13176, W8149, W8148, W13178, W8133, W18837, W13203, W13205, W13208, W13209, W13210, W4543, W18840, W4545, W18829, W18827, W4548, W13217, W18824, W18822, W13219, W4532, W18856, W13192, W18852, W4529, W13194, W18850, W13195, W18847, W13168, W13196, W4535, W18844, W18842, W4537, W13198, W4538, W4539, W18954, W13148, W18963, W18962, W18959, W18957, W8180, W4435, W18956, W4436, W13146, W4437, W8179, W18952, W13154, W4444, W13156, W4449, W4421, W8187, W13137, W13138, W18980, W18979, W8185, W4420, W4450, W4422, W4424, W8184, W8183, W13143, W18910, W4465, W18923, W18920, W4467, W18916, W4468, W8168, W4478, W4462, W18909, W8160, W18907, W8158, W13166, W4483, W4485, W13167, W18932, W18944, W8176, W18942, W18941, W8171, W18937, W4456, W13161, W13220, W18931, W18930, W8170, W4459, W18928, W18927, W4460, W13281, W4633, W18696, W8105, W8099, W4634, W13278, W13273, W13282, W18686, W18680, W18678, W18676, W18675, W18709, W18721, W18716, W8109, W18713, W13260, W13261, W4620, W13266, W4627, W8106, W4630, W18703, W13272, W18702, W18700, W18640, W8079, W13303, W13308, W4663, W18638, W8078, W8076, W4668, W18633, W13310, W8074, W8089, W18673, W4646, W13289, W13290, W13292, W4649, W18669, W18667, W13259, W18662, W18661, W8082, W4656, W18652, W18650, W13235, W13228, W8124, W4574, W4576, W18780, W18778, W18793, W18777, W8120, W4582, W13240, W4584, W13242, W13245, W4556, W4558, W18816, W13222, W13225, W8127, W18809, W18804, W18768, W4562, W18801, W13227, W4567, W18795, W18794, W8126, W18736, W18745, W18744, W4598, W8113, W4601, W4606, W8112, W8116, W18734, W4612, W18729, W13256, W18725, W13257, W18767, W8119, W18763, W4592, W18760, W13248, W18759, W13132, W4593, W13249, W8118, W18752, W18748, W13251, W4248, W4244, W13050, W4245, W8252, W13052, W19213, W13053, W19208, W4246, W19217, W13054, W19203, W19202, W19201, W19200, W13055, W19198, W19235, W8260, W8258, W19230, W19227, W19226, W13040, W13044, W19220, W4242, W13048, W13071, W8244, W13067, W19180, W19177, W19175, W19173, W13070, W4270, W19170, W4276, W4277, W8243, W13074, W4261, W19196, W4251, W4252, W13058, W8247, W4256, W4257, W4258, W13033, W13059, W19190, W4264, W19187, W19186, W13064, W4268, W4269, W12990, W4167, W19286, W19285, W19281, W12987, W8288, W19280, W19279, W19288, W4177, W12996, W4179, W12997, W12998, W4182, W8285, W19301, W8292, W12982, W4156, W4157, W4160, W4161, W8290, W19303, W13000, W19300, W19294, W19293, W4163, W19291, W4165, W19290, W8289, W19245, W4212, W19248, W19247, W8267, W4218, W4220, W8263, W4223, W13021, W8261, W19243, W13025, W13026, W19240, W13028, W13032, W13011, W19269, W13001, W19265, W4189, W8281, W19263, W8279, W4205, W4207, W4208, W19257, W8277, W4209, W13019, W8274, W8200, W8203, W19049, W19048, W4366, W4367, W4372, W19043, W4374, W19041, W4364, W4376, W4380, W4385, W4387, W19031, W19029, W19063, W19069, W13107, W4354, W8210, W19067, W8208, W8205, W19064, W19027, W13112, W19057, W4359, W19055, W19053, W4408, W13124, W4400, W8192, W4402, W4404, W19003, W13125, W18996, W8193, W13128, W18993, W18989, W18988, W13129, W8189, W18986, W19017, W4393, W19026, W19024, W19022, W19021, W19019, W19070, W8197, W4395, W19013, W8195, W19012, W8194, W4397, W19119, W19131, W19129, W4308, W19124, W13081, W8231, W13085, W4313, W4316, W8229, W19117, W8227, W19113, W4319, W8226, W19152, W4280, W4281, W4283, W4285, W4287, W19157, W19156, W4293, W19109, W19150, W19146, W19144, W8237, W13076, W13077, W8236, W19134, W4342, W13100, W4337, W4338, W19080, W13102, W8216, W19089, W19076, W4345, W4346, W13104, W19072, W8214, W4350, W4326, W19108, W4321, W4323, W4324, W19098, W13092, W8223, W4670, W8221, W4328, W19096, W8219, W4335, W19094, W13095, W19090, W13545, W13540, W13541, W4954, W4956, W13543, W13544, W18147, W4957, W18162, W18145, W4958, W18138, W4959, W4960, W18137, W4961, W13549, W4939, W4925, W4927, W13529, W18182, W4931, W13531, W13532, W7935, W4965, W18177, W4943, W4945, W4947, W18164, W7932, W13575, W4976, W4978, W4979, W18112, W4981, W18110, W4983, W7911, W7910, W4985, W7909, W18105, W13579, W4993, W4994, W13561, W13555, W13557, W18124, W4966, W4968, W4969, W18185, W18116, W13563, W4970, W4972, W7915, W13571, W7913, W4975, W7964, W13494, W18257, W4891, W18254, W18249, W13499, W18248, W18260, W7963, W4900, W18241, W18235, W18234, W18233, W7969, W7970, W18275, W18274, W13487, W18270, W13488, W18268, W4884, W4901, W4885, W4886, W13489, W4888, W7968, W7966, W18199, W4918, W18205, W7946, W13517, W4920, W18203, W13520, W7952, W18197, W18196, W13524, W13525, W7937, W18187, W13527, W4908, W4902, W4903, W18226, W7957, W7956, W13504, W13505, W7955, W18101, W4909, W18216, W4912, W4915, W7953, W4916, W13516, W5059, W17997, W5048, W17995, W13629, W5054, W17988, W17987, W7870, W13632, W18000, W17982, W7864, W17976, W13634, W5066, W5067, W5069, W17969, W18020, W13621, W18018, W5039, W5040, W18015, W18014, W18013, W17967, W18010, W5042, W13628, W18007, W18005, W18004, W7873, W13656, W5086, W17937, W5089, W17933, W7846, W13655, W13647, W7845, W5092, W5100, W17922, W17921, W17950, W13635, W5073, W17960, W17959, W7858, W17953, W7876, W5076, W13638, W7851, W13643, W7850, W13644, W5084, W13598, W18074, W5009, W5011, W18070, W18069, W13597, W7898, W13600, W18062, W5015, W13601, W5018, W18057, W18099, W13583, W13584, W13585, W13586, W5002, W18091, W18090, W13602, W18087, W13588, W18085, W18084, W7904, W18079, W13595, W13614, W18042, W18039, W5028, W7884, W13612, W18031, W13613, W18043, W7881, W13615, W7880, W7879, W5034, W7878, W5022, W18055, W5019, W7896, W7894, W18051, W7892, W18049, W5021, W7972, W5024, W18048, W7888, W5026, W18047, W18046, W5027, W18494, W18504, W13359, W13361, W4740, W18502, W4741, W18499, W18498, W13365, W13368, W18489, W13369, W8037, W18486, W13374, W8046, W4725, W18530, W18527, W8053, W8052, W8049, W18484, W18515, W4731, W18512, W18511, W18510, W18509, W13357, W18508, W13394, W8028, W13391, W8027, W18463, W13393, W18461, W4777, W4768, W18457, W4778, W4779, W4781, W13398, W18453, W8031, W18483, W4750, W18482, W13377, W13381, W4754, W4756, W4757, W18535, W18475, W18474, W13386, W4763, W18469, W13388, W4766, W4767, W18596, W13323, W18605, W18604, W8069, W4691, W18602, W18601, W8066, W18597, W4687, W13327, W18594, W4695, W4696, W13329, W18590, W18589, W18620, W4673, W13311, W18629, W8073, W4678, W13312, W4682, W8071, W4683, W13320, W8070, W13321, W4686, W18548, W13344, W18556, W18555, W18554, W4717, W13348, W18550, W4718, W18557, W18546, W4719, W4722, W4723, W18541, W18539, W18536, W4724, W8059, W4705, W8064, W4706, W13332, W8063, W13336, W18572, W18450, W4712, W8057, W18565, W8056, W13341, W8055, W4840, W4842, W4843, W7987, W18337, W7984, W4845, W18343, W13465, W7983, W18327, W7981, W18323, W13467, W4851, W18352, W13452, W13453, W18361, W4833, W7991, W18355, W13457, W18354, W7980, W7990, W4837, W7989, W18344, W18286, W4866, W18297, W18294, W18293, W4869, W18288, W4875, W18301, W18282, W18280, W18279, W7973, W18277, W13484, W13474, W18318, W18317, W13470, W4855, W13473, W18310, W18365, W18308, W18307, W13475, W7978, W13478, W4864, W4865, W13418, W4798, W18425, W4799, W13412, W13413, W4802, W13417, W18428, W4804, W8010, W13424, W13425, W18414, W4811, W13427, W18438, W18447, W13408, W4791, W4793, W4795, W18442, W18440, W4797, W18410, W13409, W18437, W18436, W18435, W18433, W13410, W7998, W18384, W4824, W18381, W13436, W18380, W7999, W4827, W13435, W13442, W13443, W13444, W4828, W13445, W13446, W7997, W13451, W4818, W4814, W8006, W8005, W13430, W4816, W8004, W18398, W18395, W4820, W18394, W8003, W13433, W18388, W18387, W18385, W3469, W3461, W3462, W20275, W12503, W12504, W3467, W12505, W12506, W3460, W3470, W8598, W8595, W3471, W3473, W8594, W3474, W3475, W3451, W20294, W20293, W20292, W3447, W12497, W20291, W3449, W20289, W20263, W12498, W3453, W3454, W20281, W3457, W12502, W20279, W8586, W20240, W8588, W20238, W20237, W12522, W20233, W20232, W12526, W12520, W3499, W8584, W8578, W12528, W3503, W12532, W12533, W20222, W3482, W20261, W20260, W12508, W3479, W12509, W12510, W12511, W12512, W12519, W8591, W3484, W3487, W20247, W3404, W12467, W3399, W20358, W20357, W8621, W3401, W12470, W20364, W20341, W8619, W8617, W12475, W3411, W3412, W8616, W8632, W12456, W12457, W3377, W3378, W12459, W20383, W3382, W3384, W12476, W3386, W8629, W8627, W20376, W8622, W3394, W3395, W20365, W20305, W20313, W8608, W3436, W3437, W12489, W20307, W8605, W3440, W3433, W20303, W20301, W3444, W20300, W20298, W12493, W3445, W12496, W20322, W12477, W20330, W3417, W20328, W12478, W8614, W20326, W20324, W8575, W12480, W3420, W20321, W3424, W12482, W8610, W3428, W20099, W12582, W20105, W3594, W8541, W20104, W3595, W12586, W12588, W12590, W20111, W3602, W3604, W20095, W3607, W20091, W12595, W20126, W20125, W3577, W20118, W12574, W3583, W12596, W8548, W12577, W8543, W3587, W3591, W12580, W20058, W12611, W12612, W8528, W3629, W12616, W3636, W20062, W20059, W12609, W8526, W20054, W8520, W3642, W20050, W3645, W12603, W12599, W12601, W3613, W20086, W8532, W3614, W20084, W20129, W12605, W3619, W3622, W20078, W20076, W20074, W8530, W8570, W3520, W3524, W3527, W20194, W3528, W20190, W8572, W3531, W12543, W3535, W3537, W20182, W3538, W3539, W8569, W3512, W20217, W3507, W20214, W20213, W12535, W20210, W3509, W3510, W20177, W20206, W20204, W8574, W12538, W20200, W3517, W3518, W12560, W20152, W12561, W20151, W3566, W3567, W12564, W12556, W20146, W3571, W20142, W8561, W8559, W20137, W12569, W8557, W3555, W8564, W20176, W12549, W12550, W3553, W20167, W12454, W12552, W20163, W3559, W3560, W12553, W12554, W20156, W20625, W20636, W20634, W20631, W20630, W8729, W8727, W3205, W3206, W12360, W8732, W3207, W3208, W20623, W3211, W20619, W20618, W3212, W3214, W3193, W20661, W3187, W20655, W20653, W3191, W20652, W3192, W20614, W12355, W20648, W20646, W3195, W20643, W3196, W8738, W8735, W8704, W20595, W20592, W20590, W20589, W3233, W20581, W12370, W20574, W8703, W3241, W20570, W20569, W12382, W8700, W3221, W12367, W3215, W20609, W8720, W3216, W20607, W3220, W20606, W12352, W3222, W3224, W20601, W20600, W8712, W20598, W20597, W3230, W8774, W20728, W20725, W12311, W3142, W3146, W12312, W3148, W20719, W20730, W8772, W8768, W20713, W3155, W20710, W8764, W20709, W12298, W3129, W20749, W8781, W20747, W12300, W3160, W8780, W20739, W20736, W20735, W20734, W3140, W20733, W20732, W12346, W12333, W12337, W8749, W20681, W8748, W20680, W20679, W3177, W20683, W20674, W8743, W12349, W3179, W20666, W20665, W3181, W3182, W20695, W3161, W12317, W8757, W20697, W3162, W3245, W20694, W3165, W12328, W20691, W20687, W3172, W3326, W20459, W3330, W3331, W8659, W12434, W20451, W20462, W3337, W8657, W3341, W20442, W3343, W8656, W20433, W20432, W3320, W20482, W20481, W20480, W12427, W20474, W20472, W20471, W20470, W20431, W20468, W20467, W3321, W3322, W20465, W3324, W20464, W3325, W3370, W3361, W3362, W20403, W3363, W12451, W3369, W8639, W20398, W20395, W3371, W8635, W20389, W8633, W8647, W20429, W20428, W3345, W8650, W12437, W8649, W8648, W12441, W20483, W20416, W3355, W20415, W8646, W12447, W8643, W20409, W8641, W8684, W8694, W20541, W20540, W3269, W3272, W3273, W3275, W12396, W3264, W20532, W20529, W20528, W3280, W20525, W12399, W20518, W12401, W3258, W3253, W20564, W20561, W20560, W3254, W12387, W3255, W3281, W20553, W20551, W12388, W12389, W3260, W20545, W3262, W8695, W20490, W20498, W20497, W3298, W8673, W20493, W3305, W20499, W8671, W3309, W20486, W12424, W3312, W3313, W8667, W8666, W12404, W20514, W20513, W20512, W8680, W12405, W3286, W12406, W8517, W8679, W20507, W8677, W20506, W12412, W3294, W20503, W19572, W3974, W3975, W3976, W8374, W19580, W8373, W3978, W3979, W12860, W8376, W12862, W19567, W12863, W8370, W3984, W19562, W12867, W12845, W8382, W3962, W12851, W3964, W19595, W19593, W19555, W8380, W19591, W8377, W19590, W19588, W12854, W3972, W4007, W19530, W8360, W19527, W8359, W19525, W12891, W19523, W12892, W12884, W19520, W12894, W12896, W8352, W4012, W4013, W8349, W12873, W12876, W12877, W3995, W19547, W12878, W8389, W8366, W8365, W19539, W12879, W8364, W12882, W3906, W19678, W3902, W3903, W3904, W19671, W19667, W8400, W19666, W19664, W3909, W8395, W3911, W12818, W12819, W12821, W19700, W19698, W12797, W8410, W12799, W8408, W3894, W19649, W3897, W8404, W19683, W19682, W8401, W19681, W19680, W12810, W12836, W3941, W19623, W3942, W3943, W8391, W3947, W19613, W19628, W3950, W19612, W3952, W3953, W3956, W19609, W19608, W3923, W19648, W19646, W3915, W3916, W12823, W3921, W19511, W19631, W3929, W12826, W12829, W12831, W3938, W19629, W19397, W8314, W4098, W4100, W4101, W19391, W12936, W4104, W4105, W4095, W8310, W8308, W8307, W19377, W4111, W19374, W8305, W12929, W4078, W12922, W12925, W19415, W19414, W8322, W8320, W19413, W12930, W4084, W19407, W8318, W4090, W19403, W19399, W8295, W4130, W4133, W19331, W4134, W19330, W4135, W4138, W4127, W8294, W4140, W19323, W8293, W4145, W19356, W19367, W19364, W8304, W19358, W8301, W8327, W12952, W12962, W19351, W4119, W19343, W8300, W4120, W12968, W19476, W19485, W4029, W12903, W4032, W4033, W4036, W12904, W4037, W19477, W4028, W19474, W4038, W19473, W8332, W4046, W19467, W19496, W19508, W12899, W8348, W4021, W8346, W19502, W19501, W4047, W19494, W4026, W12902, W8344, W4027, W19488, W19487, W12916, W19437, W4062, W19433, W4066, W4067, W4069, W19428, W4072, W19421, W19420, W19419, W4076, W8328, W4077, W19456, W8331, W4050, W19460, W19459, W12909, W19457, W12910, W4054, W12795, W4058, W19452, W19451, W12912, W19447, W19446, W4059, W19441, W8466, W3718, W19940, W3722, W3723, W19934, W19930, W8467, W19942, W19923, W12682, W19922, W3728, W12684, W19916, W19915, W19954, W19966, W19964, W19962, W8484, W3703, W8482, W19956, W12676, W19949, W3711, W19948, W19946, W3714, W19944, W19889, W19897, W8457, W19895, W12689, W3753, W19890, W3747, W12691, W12693, W3755, W19880, W19876, W19908, W3734, W12685, W3735, W3737, W19909, W3738, W19967, W3739, W12686, W8460, W3746, W8458, W19903, W19902, W12639, W20023, W20022, W20020, W20019, W3658, W3662, W20017, W20016, W3664, W20025, W3666, W3667, W8504, W20013, W8503, W8502, W20046, W20044, W20041, W20039, W12644, W20035, W8508, W12635, W20029, W8507, W3655, W8506, W3693, W12657, W19985, W25342, W12661, W12667, W12668, W12656, W3694, W19974, W3695, W3697, W3699, W3701, W19997, W20009, W20008, W3673, W20006, W3674, W20004, W12645, W12646, W12696, W12650, W3677, W8497, W12652, W19989, W8495, W3841, W19765, W12761, W19764, W8420, W19761, W12762, W19759, W8422, W3842, W19757, W19753, W19751, W8417, W19745, W19787, W8430, W3824, W19792, W3825, W12745, W12746, W12747, W12748, W19744, W12749, W12751, W8425, W19780, W19773, W12756, W3869, W12787, W19714, W19713, W12789, W3867, W19712, W3868, W12790, W19708, W12791, W3879, W3880, W3888, W8415, W19742, W19741, W12765, W12771, W12772, W3844, W19735, W12777, W3819, W12779, W3848, W12782, W19725, W12785, W3857, W3860, W19844, W8450, W19853, W19850, W19848, W12707, W3772, W12708, W8447, W3770, W12715, W3779, W3780, W12716, W19842, W19840, W3784, W12721, W19865, W3758, W19873, W8453, W8452, W19869, W3762, W19867, W3763, W8451, W3765, W3766, W3767, W3769, W3813, W8433, W19807, W19806, W19805, W12734, W3809, W3812, W12731, W19802, W3815, W19800, W3817, W12738, W12741, W3818, W3799, W12724, W19834, W19832, W3794, W19828, W8440, W5101, W19821, W19814, W12728, W8438, W8437, W19808, W6376, W6377, W14518, W7252, W6379, W15918, W15917, W7248, W15928, W6382, W6384, W14522, W15907, W7246, W14525, W6393, W14499, W15952, W15951, W6349, W7272, W14493, W15946, W6353, W6359, W15902, W14501, W6368, W14510, W14514, W7260, W15930, W15929, W15871, W15870, W15869, W15864, W15863, W15862, W14536, W6411, W15856, W15854, W15853, W6412, W6413, W14539, W6415, W6398, W14528, W15898, W7243, W15894, W7242, W6404, W15891, W7273, W15888, W14533, W7241, W15882, W6406, W15879, W15876, W14474, W7290, W7288, W14472, W6307, W14473, W6308, W7291, W15995, W7283, W15994, W6316, W15989, W6317, W6318, W16023, W14455, W14456, W14458, W6283, W6284, W14460, W6320, W6288, W16018, W6289, W6290, W6291, W6295, W14461, W7292, W7278, W6335, W7280, W14485, W15963, W15962, W6338, W6340, W14484, W15958, W14488, W7275, W6346, W15956, W6347, W6348, W6328, W14476, W6321, W14477, W6322, W15982, W6323, W14478, W15845, W14479, W6331, W15976, W6332, W14482, W15972, W15971, W15969, W15726, W15744, W7214, W6489, W15739, W15737, W15734, W7211, W6493, W15728, W15746, W7210, W6494, W6496, W15721, W7208, W6482, W15765, W15762, W15756, W15755, W14572, W15717, W15751, W14573, W15750, W15749, W6485, W6486, W14578, W15674, W14597, W15685, W15684, W6512, W15681, W6514, W7198, W15689, W15673, W14603, W6516, W15669, W6518, W6522, W6523, W14594, W6498, W15714, W15710, W15708, W6500, W15706, W14590, W15701, W6479, W14596, W6507, W7200, W6508, W15693, W15692, W6511, W7228, W6437, W15820, W14545, W6439, W14546, W6440, W7229, W6441, W14543, W6443, W6444, W15810, W15809, W14549, W15807, W15806, W15805, W7231, W6416, W6417, W6419, W15843, W15840, W15839, W6420, W15804, W6424, W6426, W6429, W15830, W14541, W15829, W6431, W15828, W14568, W6461, W6462, W6465, W15782, W6466, W7222, W15778, W6460, W15775, W15774, W14569, W15772, W6468, W6474, W7219, W6478, W14554, W14550, W15801, W15800, W14551, W15799, W15797, W6277, W14555, W6453, W14556, W15793, W6457, W7224, W15786, W6459, W7364, W6124, W14367, W16311, W6132, W14374, W16298, W7365, W16296, W7368, W6136, W14375, W16292, W14377, W16291, W6141, W14378, W6144, W14360, W16339, W16338, W16336, W14356, W14358, W16331, W6114, W6118, W6149, W14361, W16324, W16323, W16321, W6122, W16317, W6123, W6176, W16260, W16259, W6173, W6174, W16255, W6175, W16247, W14384, W16246, W7347, W6179, W7346, W6181, W16232, W16285, W6152, W6153, W14379, W16278, W16277, W14382, W6108, W16273, W7356, W16268, W6168, W6169, W6171, W16262, W6067, W7390, W14316, W14318, W14322, W16419, W6064, W16416, W16428, W14334, W14335, W16401, W7381, W7380, W16396, W16395, W6078, W16436, W16452, W16449, W16448, W16442, W14306, W16440, W16439, W16389, W6053, W16433, W16432, W6056, W6057, W7391, W6060, W16429, W6098, W16362, W6099, W14345, W14347, W6104, W14351, W7374, W16345, W14354, W16343, W6107, W6086, W6079, W7376, W16387, W6084, W16381, W16379, W6085, W14389, W6087, W7375, W16374, W6092, W16372, W6095, W14341, W14342, W16090, W16095, W7311, W6246, W6247, W16094, W6249, W14431, W14434, W16097, W14435, W16085, W16084, W7309, W6253, W6254, W6255, W14438, W6229, W14418, W6232, W14419, W6234, W6236, W16109, W6237, W16108, W6239, W14423, W14424, W6243, W14425, W16100, W14428, W14453, W16049, W16048, W14452, W16046, W16053, W6274, W6275, W16039, W16037, W16036, W16035, W16033, W6264, W14439, W16073, W6256, W6257, W7308, W14444, W16069, W6261, W14417, W6265, W16061, W7298, W14447, W6269, W7297, W6197, W16205, W6193, W6194, W16201, W14393, W16198, W7336, W16196, W14395, W6192, W6198, W6199, W16183, W16180, W16179, W6200, W7329, W16175, W16221, W6184, W16231, W6188, W7339, W16227, W16226, W16223, W16172, W16218, W16216, W16215, W6189, W16212, W14392, W14411, W16138, W14409, W6215, W6217, W16131, W16139, W6221, W7317, W6222, W6223, W6225, W6226, W7315, W14416, W6205, W16171, W7325, W16160, W16156, W14407, W16151, W16150, W6204, W14610, W6206, W6208, W16147, W16144, W6209, W16142, W16141, W14819, W15167, W6830, W15166, W15164, W15163, W6831, W15157, W7034, W6829, W15154, W15153, W15152, W6834, W14821, W7028, W14822, W15184, W6814, W6816, W6818, W14810, W7043, W7042, W6824, W6841, W6825, W15179, W15176, W15171, W15170, W14839, W15120, W6856, W14837, W15118, W15117, W6859, W7024, W7022, W6861, W6862, W15104, W6864, W6866, W14840, W6868, W6844, W15144, W6843, W15139, W7027, W14828, W15134, W6813, W14830, W14832, W7026, W6852, W15129, W15127, W15124, W14787, W14782, W6763, W6766, W6767, W15252, W6768, W14784, W14786, W7068, W6775, W15243, W15242, W14790, W6781, W15266, W15273, W14768, W15272, W7071, W15271, W15270, W15269, W14770, W6785, W14774, W14776, W15264, W15263, W6757, W15261, W7070, W15259, W14805, W7051, W15210, W15209, W15206, W15203, W6802, W6803, W15215, W14806, W7047, W15200, W6809, W15196, W15195, W15194, W15193, W15226, W14793, W7060, W6789, W15233, W14796, W15228, W6792, W15227, W6869, W15224, W15220, W6796, W7054, W15218, W6798, W7053, W14950, W6953, W14960, W14959, W6954, W14954, W14953, W14887, W6991, W14962, W6957, W14889, W14949, W14947, W6989, W14891, W6938, W14984, W6940, W14876, W14982, W6948, W6949, W14940, W14973, W14972, W14969, W6995, W14968, W14966, W14883, W6952, W6985, W14921, W14920, W6975, W14899, W6979, W6980, W14916, W6981, W6973, W14902, W14906, W6982, W6983, W6984, W14903, W14904, W14894, W14939, W6958, W14937, W14892, W14936, W14893, W6961, W6962, W14989, W14895, W6964, W14896, W14933, W14926, W6988, W14898, W14923, W6894, W15071, W14843, W14848, W6889, W14850, W6890, W7014, W6891, W6893, W6886, W14855, W6897, W15049, W15046, W15045, W6903, W6905, W15083, W6870, W15094, W15092, W15090, W15089, W7019, W6873, W15040, W14841, W6878, W15080, W6879, W6881, W6882, W7017, W14868, W15016, W15014, W7003, W6927, W15004, W6930, W14998, W15019, W14996, W14995, W14994, W14871, W14874, W14991, W14990, W6935, W15027, W14856, W15039, W14857, W7008, W6907, W14858, W6911, W7073, W6912, W7007, W6915, W14860, W6920, W7005, W15538, W15551, W15549, W6606, W15545, W15544, W14652, W15542, W14654, W15536, W15533, W7169, W15528, W15527, W15526, W7168, W14639, W6590, W7175, W15567, W15566, W15565, W15564, W6595, W15563, W14662, W14640, W15561, W15560, W6597, W15559, W14642, W6600, W15554, W14677, W6625, W6627, W14670, W14672, W7163, W15488, W15487, W15495, W15485, W14678, W6640, W7158, W14679, W7156, W6641, W15479, W15516, W15524, W14663, W7167, W14667, W6617, W6619, W15517, W15569, W15513, W15508, W15507, W15504, W6621, W15501, W6624, W15497, W15633, W14620, W15641, W6553, W15639, W15638, W6556, W6558, W6561, W15634, W15644, W15632, W15630, W15628, W15626, W6562, W15623, W14616, W15660, W6525, W7193, W7191, W6528, W15652, W6565, W6531, W15650, W14618, W6545, W6546, W15646, W6547, W6550, W15580, W15593, W6574, W6575, W14631, W6576, W15591, W7179, W15585, W14632, W14636, W6586, W15575, W7176, W14638, W15605, W15621, W15619, W7183, W15615, W6568, W15478, W14628, W7182, W15603, W6571, W15602, W15597, W6572, W14733, W14734, W6708, W15339, W15338, W14736, W15337, W6705, W7091, W15325, W6718, W7087, W15317, W7097, W15367, W15366, W15365, W15361, W7099, W6693, W6697, W6699, W14741, W15351, W6701, W15350, W6703, W7093, W15346, W15345, W6704, W14752, W14756, W15290, W14757, W15286, W6742, W14762, W6745, W15293, W14765, W15279, W6746, W15278, W14766, W6747, W14767, W6734, W6722, W6723, W15315, W15309, W6728, W6730, W6733, W15368, W14745, W6735, W15303, W15299, W6736, W7078, W15428, W7139, W6659, W7137, W7135, W7134, W15434, W15430, W15440, W14695, W7131, W15419, W15416, W15415, W6668, W14699, W15461, W7155, W6643, W7152, W15465, W15464, W7149, W6654, W15452, W6657, W7143, W15441, W7142, W15384, W15393, W6677, W7116, W7115, W15391, W15389, W15385, W15394, W6683, W6685, W14722, W14723, W15373, W7104, W15369, W15409, W7124, W15413, W7122, W14709, W6672, W14711, W15410, W16453, W15408, W7118, W15406, W15405, W14713, W15401, W6676, W15398, W13885, W17473, W7696, W5402, W7694, W5406, W7693, W7691, W13880, W17464, W17461, W13886, W5415, W17458, W7688, W7685, W7684, W17451, W17494, W13875, W5394, W7699, W17491, W5395, W17487, W17484, W17450, W17483, W17482, W17481, W5397, W5399, W7697, W5436, W17414, W5427, W17413, W7674, W17411, W7673, W5430, W17405, W17416, W7669, W17402, W13904, W5437, W5438, W17391, W17390, W17434, W17449, W17447, W17445, W17444, W17441, W7680, W5421, W5390, W17431, W17430, W5423, W17425, W5424, W17418, W17535, W5345, W5347, W17543, W7713, W17539, W5352, W17536, W13847, W13853, W17534, W5357, W17531, W13855, W7709, W13857, W7715, W7721, W17566, W17563, W13835, W7718, W7716, W13838, W17561, W5362, W17557, W13840, W5338, W17555, W17554, W17553, W13843, W7714, W13872, W13870, W17504, W5374, W7704, W5375, W7703, W5380, W7701, W17501, W17500, W17499, W5388, W17498, W13873, W17496, W5389, W17513, W17525, W5364, W5366, W13862, W17516, W5367, W7666, W5369, W5372, W13866, W17508, W17507, W5373, W5512, W5504, W5505, W17284, W13951, W17277, W5507, W17273, W5511, W17271, W5503, W17268, W5513, W5514, W7624, W13956, W5516, W5499, W13947, W17307, W17305, W17304, W7629, W17298, W17266, W17296, W17293, W17291, W17290, W17289, W7628, W13950, W17286, W17234, W13973, W5535, W17242, W5536, W17241, W13977, W5538, W17233, W7616, W7615, W5544, W17231, W7614, W17229, W17228, W5521, W17265, W13958, W5520, W17261, W17260, W17259, W13960, W5496, W13961, W17253, W5526, W7618, W5529, W17249, W5532, W5464, W13915, W13920, W13921, W17359, W5463, W17354, W17353, W17351, W17363, W17350, W13922, W17348, W7647, W13923, W5467, W7646, W5454, W17389, W5443, W13910, W7659, W7656, W7654, W17382, W7653, W5470, W5455, W17379, W17377, W5456, W17375, W17374, W17371, W17370, W17319, W5483, W17329, W5487, W17327, W13935, W5490, W17320, W13933, W17318, W5491, W17316, W7632, W13942, W13943, W5493, W13946, W17335, W5471, W17343, W5474, W5475, W17340, W13928, W5476, W7644, W5329, W13929, W17334, W5478, W17332, W7643, W5480, W13932, W7810, W13713, W13715, W7817, W17814, W7816, W5180, W5181, W7811, W5183, W5177, W17806, W13722, W7809, W17801, W13727, W17798, W17794, W5188, W17831, W17837, W5164, W17835, W5166, W13706, W17832, W5167, W7825, W5170, W17829, W5171, W7824, W5173, W7820, W13712, W5176, W17756, W17766, W5203, W17763, W7797, W5205, W17759, W17758, W17754, W13739, W5208, W13741, W13743, W5209, W5214, W17777, W5190, W7805, W17784, W17782, W5192, W7804, W17780, W17840, W5196, W17775, W17774, W13730, W5199, W5201, W17770, W7799, W17886, W5123, W5124, W5125, W7835, W5128, W17890, W13676, W17889, W5122, W17884, W7834, W5130, W17881, W17879, W5132, W5133, W13667, W13661, W5106, W17916, W13662, W17915, W13663, W5114, W17913, W13670, W17909, W7840, W17904, W13674, W17903, W5121, W7836, W17847, W13690, W13694, W13695, W5157, W17850, W17849, W17848, W5153, W17846, W17845, W5160, W13705, W17841, W17866, W17873, W5136, W5137, W7831, W17870, W17867, W13684, W17738, W17865, W17863, W17857, W7829, W5148, W13689, W17855, W5296, W7738, W5287, W17641, W5290, W17640, W5291, W5293, W17636, W5294, W5285, W17631, W7737, W17628, W17626, W7733, W5302, W13813, W5273, W7755, W5265, W17653, W5268, W17651, W5271, W7752, W17621, W7748, W5279, W7747, W5283, W7746, W5284, W17580, W17589, W13832, W5316, W17587, W17584, W17583, W7722, W7723, W17579, W17578, W5326, W17575, W5327, W17572, W17571, W17568, W17601, W13814, W17615, W17614, W17613, W17607, W17606, W5306, W5262, W13818, W13820, W7726, W17595, W5313, W5314, W13827, W7776, W17716, W13758, W17712, W13759, W17709, W7778, W17708, W5228, W5229, W7780, W5232, W17701, W5234, W5236, W17697, W17694, W17693, W7788, W7791, W17736, W7789, W17732, W17730, W17728, W17727, W13750, W5216, W7786, W7785, W7784, W7782, W5220, W7781, W5221, W17668, W17674, W7761, W7759, W5255, W13784, W17672, W17671, W5256, W5257, W17665, W13791, W17663, W17661, W5260, W5261, W17681, W17691, W17690, W13770, W17688, W13771, W17685, W13774, W7764, W13983, W7763, W17680, W5242, W17679, W13777, W13778, W5245, W17677, W16705, W5890, W5894, W16716, W5895, W16715, W16713, W16710, W7462, W14207, W14210, W7459, W16704, W16703, W14216, W16699, W16698, W7455, W14206, W14200, W7468, W5879, W14202, W16735, W5880, W14219, W16733, W5883, W5884, W5885, W5886, W7466, W16724, W5922, W7450, W5917, W5921, W14232, W5914, W5924, W16659, W14234, W5926, W5930, W5931, W7448, W16689, W16696, W5902, W14220, W5906, W7453, W7452, W16690, W7469, W5908, W5910, W14225, W14227, W5913, W16680, W16679, W16807, W5826, W7499, W5828, W5829, W16814, W16813, W14165, W16810, W14167, W14161, W16806, W14168, W5837, W16800, W5846, W14170, W5815, W14154, W16841, W16840, W16839, W16838, W5812, W14155, W16836, W16833, W5818, W16827, W16826, W5819, W16821, W5821, W5870, W5861, W5862, W5863, W16759, W16755, W5869, W16764, W16746, W14184, W14186, W14187, W14196, W7485, W5851, W16792, W5852, W16791, W16783, W7488, W5856, W7487, W5935, W5858, W16776, W16775, W16770, W16766, W6022, W16526, W14288, W6019, W16520, W7414, W16516, W6021, W16528, W6023, W16512, W14291, W14294, W6026, W6028, W16555, W6006, W16549, W6010, W6011, W16545, W6029, W6012, W6013, W16532, W6015, W16469, W14299, W16479, W14300, W7403, W16473, W6045, W16470, W7404, W16468, W16463, W16461, W14302, W16458, W16454, W6048, W6049, W6036, W7410, W16503, W16502, W7409, W16500, W14297, W6035, W16497, W7406, W16496, W6039, W16489, W16488, W6040, W6041, W16484, W16609, W5954, W16619, W5955, W16617, W16616, W5956, W16611, W16610, W7438, W5957, W7436, W14256, W7433, W14258, W14259, W14261, W5937, W14239, W16642, W7445, W16640, W14244, W5944, W16638, W16604, W14246, W5946, W5948, W14247, W16631, W16628, W16627, W14249, W16570, W14269, W14270, W5983, W16573, W5986, W16571, W5987, W16579, W16568, W5994, W14273, W7424, W5996, W16565, W5997, W14276, W16594, W16603, W14263, W5963, W14264, W16597, W14265, W7509, W16592, W7428, W16587, W16586, W16584, W5973, W14048, W17106, W14044, W14045, W5630, W17101, W17100, W14046, W17097, W5632, W14040, W7568, W17092, W5635, W5638, W14056, W17089, W17088, W14034, W17122, W17121, W5618, W14035, W17117, W5647, W5619, W5621, W7577, W17112, W5623, W7573, W5674, W5668, W17059, W5670, W17056, W17055, W17054, W5671, W5673, W5663, W5675, W5677, W5678, W17047, W17046, W14074, W5681, W17044, W17079, W7566, W14060, W5652, W14061, W5653, W17081, W17080, W5612, W5655, W17077, W5656, W14067, W5661, W14068, W14069, W17065, W17193, W17191, W17188, W7601, W14002, W7599, W17179, W5568, W7602, W5570, W7597, W5575, W17165, W17163, W7592, W17161, W5578, W7610, W17222, W17220, W7607, W5559, W5561, W14008, W5562, W13996, W17203, W17202, W7603, W17194, W5608, W5602, W14023, W7582, W17140, W17139, W17138, W5607, W5601, W17136, W17135, W14025, W17130, W17129, W14033, W17151, W14010, W17158, W5587, W7590, W17152, W14017, W5682, W5589, W5591, W14018, W5595, W7585, W5598, W5599, W14022, W16901, W5758, W16911, W5761, W5762, W16906, W7518, W14137, W5769, W16902, W5757, W5773, W16894, W16893, W16889, W16887, W7513, W14125, W5743, W5745, W14123, W16932, W16930, W16929, W5752, W16928, W5778, W16926, W16925, W7523, W16914, W14127, W14128, W7522, W5806, W16867, W7511, W16865, W5800, W16861, W5797, W16858, W5807, W16856, W16855, W5808, W16851, W16850, W16849, W16876, W16883, W7512, W5781, W14146, W5784, W14147, W16880, W16875, W14148, W16874, W14149, W5792, W5793, W5794, W14150, W5702, W17015, W5697, W14089, W14090, W17012, W14091, W17009, W17008, W5701, W5704, W5708, W5709, W7541, W5711, W17000, W7540, W17031, W14075, W7551, W5684, W17037, W7549, W14081, W17034, W16995, W17030, W5691, W5693, W17026, W17022, W17020, W7545, W16949, W14108, W14110, W14114, W16956, W5730, W16953, W5731, W16951, W14117, W16945, W16940, W5735, W16936, W5740, W5742, W16981, W16994, W16993, W16991, W16988, W7538, W5716, W5717, W20185, W14102, W16979, W16971, W7534, W16967, W5720, W16966, W14105, W22911, W22902, W9466, W1669, W1668, W1666, W22904, W1665, W10552, W24576, W1663, W9963, W11306, W544, W1658, W24572, W22918, W10553, W10554, W9471, W9473, W22921, W22922, W551, W1651, W1650, W22890, W9451, W9454, W24590, W9455, W11322, W537, W24585, W1692, W10547, W9460, W22884, W1685, W22888, W1684, W1679, W1678, W11317, W10549, W22897, W9463, W11313, W543, W10551, W22900, W9465, W1634, W1633, W566, W9480, W567, W1630, W24554, W10561, W11281, W24552, W11280, W9481, W1615, W565, W22972, W1614, W11275, W11274, W1610, W1607, W9482, W22983, W9484, W1603, W24550, W11266, W22943, W556, W1649, W11299, W1648, W22931, W22932, W11297, W24566, W557, W22936, W558, W9478, W22865, W22944, W9479, W22946, W1643, W1641, W11293, W22950, W564, W22954, W1635, W22956, W11292, W24620, W22792, W1749, W22793, W10533, W22794, W10535, W1748, W11363, W520, W22796, W22797, W24622, W24621, W11362, W9419, W9426, W22801, W22803, W22808, W1746, W22811, W1744, W1743, W1742, W11360, W9429, W22814, W22815, W1763, W509, W11377, W11375, W1774, W9410, W9412, W22769, W9414, W1768, W9973, W513, W521, W1762, W1761, W22776, W1760, W1758, W22778, W9417, W11367, W22781, W22783, W22786, W1754, W9418, W24633, W9447, W529, W22840, W22841, W11340, W1718, W10545, W9441, W9445, W1714, W1712, W11337, W9446, W11334, W24596, W22838, W534, W24593, W11329, W11328, W1702, W9449, W11327, W1699, W22856, W22858, W11326, W11324, W9435, W24616, W1735, W22822, W9430, W22826, W1734, W22827, W10536, W22828, W11351, W10537, W522, W1599, W10538, W11346, W523, W22833, W24606, W11345, W22834, W525, W526, W1725, W22837, W527, W11341, W9970, W9553, W9550, W23130, W23132, W23134, W608, W10580, W23136, W11202, W9552, W11200, W609, W24494, W23149, W11196, W23151, W23155, W1508, W23156, W1507, W9557, W11189, W1504, W9558, W23164, W604, W23098, W1531, W9532, W1525, W9534, W9537, W9539, W1520, W1519, W23110, W23111, W1518, W1503, W24502, W23114, W23117, W607, W9548, W1515, W24500, W23119, W23121, W23122, W23123, W10588, W11154, W630, W23191, W1477, W23194, W24483, W10590, W631, W1476, W23199, W24479, W11155, W9567, W11148, W23208, W1470, W1468, W23211, W1466, W23218, W9569, W1463, W23224, W9570, W11171, W11186, W23165, W10583, W1497, W1495, W9937, W10585, W1493, W9559, W23169, W625, W11183, W9561, W11172, W1532, W1488, W1486, W1485, W23176, W9562, W23177, W629, W1480, W9564, W23184, W10586, W23185, W9936, W578, W24537, W24536, W9498, W9500, W23026, W1582, W1581, W23027, W9501, W1578, W23029, W23030, W1586, W579, W11246, W23031, W24535, W11245, W11244, W24533, W23034, W587, W588, W589, W573, W9960, W11265, W1596, W22996, W9488, W11263, W9489, W23002, W9490, W23006, W23007, W570, W571, W11258, W1593, W9504, W23014, W576, W11255, W9494, W10564, W23017, W11253, W1591, W11251, W24544, W9956, W9495, W23021, W24542, W596, W23068, W9516, W11226, W9517, W1549, W594, W9518, W1543, W9520, W23078, W23079, W24514, W1541, W23081, W1539, W593, W23083, W9524, W9525, W598, W23087, W23089, W10574, W599, W23091, W23094, W1534, W600, W24511, W23056, W23042, W23045, W590, W9508, W23048, W23051, W1565, W11237, W23053, W9509, W1564, W24527, W1775, W9512, W1562, W23058, W10571, W9514, W1557, W1556, W11232, W24522, W1554, W1552, W9515, W9318, W10481, W410, W10483, W1983, W10007, W413, W414, W1978, W11505, W9325, W1977, W406, W22448, W1975, W11503, W9327, W9328, W1969, W10004, W22462, W22465, W11502, W22469, W22430, W9303, W9304, W9306, W10476, W11515, W9308, W10477, W22425, W22427, W22428, W22470, W22431, W11514, W10478, W1992, W1991, W9313, W1990, W22434, W22435, W10479, W1987, W405, W11511, W1935, W10488, W9337, W9338, W22512, W1941, W10489, W11475, W24729, W9341, W22522, W1936, W22531, W11470, W11469, W11466, W22535, W22536, W22537, W11465, W1929, W22542, W22543, W1928, W11464, W1954, W1966, W1964, W10002, W421, W11497, W11495, W10485, W11492, W11490, W1956, W24738, W1996, W22486, W11487, W11486, W22491, W10486, W1949, W22494, W424, W24733, W24731, W10487, W1948, W11484, W22500, W11560, W11569, W379, W9270, W22345, W10018, W22349, W22351, W11564, W2061, W2060, W10456, W24780, W11558, W22357, W11557, W22358, W2055, W22362, W24776, W385, W2053, W11551, W386, W22328, W2077, W22316, W22318, W2075, W2074, W11580, W24788, W11578, W22320, W11577, W22324, W22326, W24787, W22327, W24772, W9264, W22330, W11572, W22333, W22335, W22336, W377, W10449, W22337, W10450, W22339, W9267, W22340, W24763, W22393, W2020, W11527, W2018, W22395, W2017, W2015, W9294, W398, W22398, W2013, W2012, W22391, W2010, W399, W22404, W2007, W22405, W2005, W11522, W11519, W1999, W10475, W22412, W1997, W22368, W11546, W22371, W2047, W10016, W11542, W22373, W11541, W10465, W9286, W10013, W2034, W9343, W2032, W22382, W11538, W9287, W11536, W2029, W9288, W11531, W2027, W10012, W2022, W9291, W11528, W11409, W11418, W483, W22675, W486, W11417, W22676, W1822, W1821, W11416, W11415, W1817, W9385, W1816, W1815, W10520, W482, W22685, W22688, W22689, W488, W24663, W490, W9388, W11406, W9389, W493, W1836, W22637, W1845, W10513, W1844, W1843, W22641, W24679, W1840, W22644, W1838, W24677, W11427, W24657, W481, W10516, W24676, W22659, W1834, W11425, W1831, W9982, W11424, W1830, W9383, W11395, W9405, W11392, W11391, W9976, W22743, W11388, W502, W22747, W22749, W11387, W22752, W1785, W11384, W9975, W1782, W9409, W10529, W24635, W506, W11381, W22759, W1776, W11379, W22724, W22702, W24656, W22703, W22706, W1804, W11401, W22710, W22714, W1802, W22720, W9395, W22723, W496, W497, W22729, W24653, W9399, W9400, W22730, W9401, W24649, W10525, W11396, W1795, W501, W22589, W24715, W1901, W438, W439, W1896, W22580, W22581, W22582, W10497, W1894, W443, W24708, W1892, W22590, W446, W11451, W10499, W24705, W1887, W22595, W1886, W11449, W10500, W22599, W450, W1884, W24722, W22545, W1926, W1925, W1922, W1921, W1920, W1917, W24725, W11462, W22555, W24723, W11448, W1911, W1910, W22558, W1909, W436, W1908, W9345, W24719, W22562, W11456, W1904, W24716, W9365, W24687, W22615, W1863, W11438, W466, W9989, W1861, W22619, W469, W22620, W24685, W470, W22614, W472, W1858, W9366, W11436, W1855, W473, W1854, W9367, W1852, W22633, W476, W11429, W1846, W10512, W11446, W451, W22602, W452, W453, W1882, W1881, W9992, W1877, W24699, W9356, W459, W460, W23228, W1873, W463, W10504, W24691, W22608, W9358, W22609, W1869, W10506, W1866, W9360, W22613, W9872, W9756, W10873, W1066, W1065, W9758, W10694, W24240, W23790, W1063, W10695, W10870, W23793, W1068, W23796, W23798, W1059, W9760, W776, W10864, W23805, W9871, W10863, W1056, W767, W1085, W9748, W10889, W9875, W765, W23768, W10886, W10692, W9750, W10884, W23775, W24251, W1075, W23778, W24248, W24243, W10880, W10878, W772, W23785, W9859, W23841, W1038, W23847, W10851, W23850, W23852, W9857, W10850, W1034, W23856, W23857, W1041, W792, W1031, W24218, W9768, W10704, W24215, W1029, W794, W9771, W10847, W1027, W795, W781, W23813, W23816, W23819, W10862, W1052, W1050, W24228, W10699, W1049, W23823, W780, W23824, W1048, W23827, W1047, W10859, W23829, W782, W24225, W10857, W23831, W1044, W785, W24223, W1156, W748, W23680, W24286, W10683, W1154, W750, W1153, W751, W1149, W23688, W1148, W744, W23692, W1146, W1145, W23694, W10920, W23695, W23698, W10684, W23702, W1140, W752, W23704, W10919, W1139, W23668, W9727, W10934, W1168, W23662, W23663, W10933, W24298, W10931, W1165, W9884, W9728, W753, W1162, W24296, W1160, W23670, W23671, W1159, W9883, W23674, W10679, W741, W1158, W23678, W10681, W9876, W10908, W9877, W1104, W23741, W24260, W10907, W1102, W761, W10905, W24259, W10902, W10901, W10900, W23739, W1093, W23750, W10898, W23752, W10689, W10691, W764, W23755, W10895, W23758, W1089, W10894, W9747, W23760, W1129, W10917, W10685, W23709, W23710, W10686, W24270, W1133, W1130, W756, W9737, W9738, W10687, W24267, W1125, W23722, W24265, W9882, W1121, W1120, W1119, W1114, W9743, W759, W1108, W10910, W1107, W907, W10778, W10777, W912, W24031, W24032, W847, W909, W24139, W10773, W24039, W24041, W24028, W848, W906, W905, W24047, W904, W903, W24137, W24136, W24135, W24134, W901, W900, W10767, W10787, W10794, W937, W840, W24159, W23999, W24000, W24001, W24157, W10792, W24006, W9807, W931, W10788, W9827, W24017, W842, W24019, W920, W918, W844, W10783, W24151, W24146, W24144, W9829, W10779, W10752, W879, W9824, W857, W24088, W877, W859, W24089, W24091, W875, W9820, W24093, W24094, W10744, W874, W881, W10745, W9821, W24099, W871, W10749, W863, W24109, W10748, W868, W10747, W24113, W897, W24059, W24060, W24131, W850, W10765, W24068, W10764, W10763, W10759, W24071, W891, W23996, W9826, W10757, W889, W888, W887, W853, W24127, W884, W854, W10753, W10742, W10743, W24121, W10721, W9848, W23906, W23907, W1000, W9786, W10718, W804, W805, W10720, W23918, W996, W23921, W23903, W24202, W993, W24201, W809, W23927, W810, W23928, W10722, W10723, W9847, W814, W23933, W10725, W987, W24209, W24212, W9851, W10842, W9775, W23870, W10838, W1015, W23875, W23878, W1014, W23881, W1013, W10707, W9844, W23883, W23884, W10710, W23887, W9850, W10831, W23890, W1003, W23893, W23894, W24207, W23898, W1002, W23902, W10804, W974, W831, W972, W969, W968, W24169, W24168, W10806, W832, W24167, W833, W23975, W963, W835, W24164, W24174, W962, W957, W10803, W23985, W10801, W944, W24161, W838, W940, W23993, W10736, W10795, W10818, W9839, W23939, W982, W23943, W23944, W824, W826, W23949, W23950, W10935, W981, W23953, W23955, W23956, W10729, W979, W24178, W23961, W977, W976, W9836, W9924, W23364, W11087, W677, W9617, W9618, W678, W9619, W9620, W23367, W11079, W23372, W1370, W23374, W1375, W9623, W1368, W23382, W11073, W1367, W1366, W24408, W23389, W10625, W680, W11096, W23330, W11109, W669, W670, W23331, W9612, W23334, W11102, W671, W23337, W23340, W1387, W1359, W9613, W9614, W9616, W23352, W11091, W1378, W23359, W24413, W11089, W672, W9925, W23434, W1320, W23421, W1319, W23422, W1317, W23423, W9639, W11043, W9917, W10633, W23432, W1321, W23436, W23438, W23439, W23443, W24389, W9911, W1308, W1305, W11039, W1341, W23395, W1354, W24406, W9630, W24405, W1350, W1349, W23404, W24404, W11063, W1344, W10626, W23411, W24420, W1337, W23412, W1335, W11058, W1332, W11055, W10632, W687, W9637, W688, W11052, W23420, W10598, W11134, W11133, W24464, W1442, W23253, W11131, W1441, W1440, W646, W1438, W10601, W9582, W9931, W1436, W23264, W1434, W11130, W1433, W10602, W24456, W10603, W649, W651, W11144, W24477, W9572, W24474, W23231, W632, W633, W10592, W1461, W635, W10593, W24471, W1458, W23238, W24470, W9933, W24467, W1456, W9576, W23245, W11138, W1450, W643, W9579, W24465, W1400, W23294, W661, W23298, W1406, W23301, W10609, W24430, W24429, W9606, W662, W23306, W1402, W10611, W11114, W23293, W23312, W23313, W24425, W664, W11111, W23316, W665, W1394, W24422, W10619, W10620, W668, W24438, W652, W1426, W653, W9591, W9929, W24450, W10605, W10606, W23273, W9596, W24446, W1421, W23276, W11036, W24434, W1413, W1412, W9928, W23279, W9600, W9601, W10608, W1410, W9603, W1407, W23292, W1209, W9699, W10663, W10973, W23577, W1211, W9702, W720, W10665, W10666, W23580, W24324, W24323, W9697, W10962, W23585, W9707, W9709, W10960, W10956, W723, W9711, W23594, W10952, W23596, W1201, W10951, W709, W23548, W23550, W1229, W10997, W10995, W24343, W9690, W24341, W1227, W1226, W711, W1221, W23567, W24335, W10658, W24329, W10988, W717, W718, W10987, W24328, W10982, W23569, W24327, W9694, W1182, W24309, W9721, W10670, W730, W23640, W735, W23644, W1174, W23646, W23648, W23649, W737, W10940, W10672, W24299, W10938, W23651, W23652, W23654, W23655, W738, W23656, W1170, W1189, W9713, W23600, W9890, W1198, W24319, W1195, W10667, W24318, W10947, W1192, W24317, W1191, W23612, W1230, W23616, W10946, W10944, W23619, W23620, W726, W1186, W727, W728, W23630, W23631, W1184, W1183, W10644, W23471, W11015, W23474, W1288, W1287, W1283, W1281, W1279, W23483, W9664, W9665, W24367, W10643, W11019, W703, W23488, W1274, W9668, W1273, W23493, W704, W1268, W9669, W23502, W23450, W11033, W11032, W24387, W9648, W24384, W692, W23455, W24380, W11028, W1297, W9908, W694, W1295, W23465, W1294, W11026, W697, W23467, W9659, W11021, W23470, W1248, W1246, W23527, W23528, W10651, W23529, W1242, W9681, W11004, W10653, W1237, W23534, W9897, W23536, W1235, W24347, W9683, W23539, W9684, W23542, W10998, W23543, W9686, W1231, W23546, W23512, W1265, W1263, W23504, W1262, W1261, W24358, W11009, W23507, W23508, W1256, W24357, W23509, W23510, W8782, W1254, W24356, W1252, W24355, W24354, W23517, W24353, W23518, W23520, W10648, W10650, W21340, W8965, W2737, W8967, W2736, W142, W2734, W12032, W10298, W21351, W21352, W25105, W2731, W21356, W21339, W8971, W21364, W8973, W12030, W12029, W12028, W144, W145, W2727, W25099, W12024, W12037, W12042, W10295, W25118, W2756, W21313, W21315, W2753, W138, W2747, W2746, W25115, W12038, W21321, W21372, W2743, W8960, W25113, W2742, W25112, W2740, W2739, W10124, W21332, W21333, W2738, W21336, W2689, W21404, W150, W151, W152, W8987, W10114, W8989, W12001, W154, W2695, W8992, W2692, W149, W156, W11997, W11995, W25082, W11994, W8993, W157, W2684, W159, W2683, W21429, W10116, W12023, W21376, W25096, W21378, W21380, W8981, W2719, W12015, W8983, W2709, W10292, W12012, W2707, W12011, W25094, W148, W8985, W12006, W21400, W25093, W2704, W21402, W21403, W21221, W2809, W2808, W21225, W8924, W12072, W21231, W2805, W2802, W12071, W2799, W8925, W21235, W8926, W2796, W21239, W2795, W2793, W110, W25149, W111, W113, W2790, W2789, W2788, W2787, W2819, W8908, W21193, W2827, W2826, W103, W21198, W2824, W104, W21200, W25164, W21201, W25163, W10132, W12082, W21208, W12077, W106, W107, W2814, W2812, W8916, W8919, W8921, W2811, W25157, W21292, W21275, W127, W129, W2770, W21281, W8943, W8944, W21287, W21289, W12048, W10128, W8946, W10284, W21293, W21294, W134, W8947, W12045, W21296, W12044, W2766, W21300, W21301, W25124, W12043, W2779, W12066, W114, W8930, W116, W21254, W8931, W10281, W25145, W21255, W2782, W12062, W25144, W2780, W21257, W11991, W118, W119, W21259, W8934, W12059, W21268, W21270, W25138, W2776, W8937, W10282, W121, W21589, W2562, W21575, W195, W2561, W21579, W21580, W10340, W25025, W10086, W11933, W25024, W9046, W196, W11932, W21587, W21590, W2554, W2552, W2549, W9054, W10347, W21600, W9055, W21601, W2547, W21605, W10082, W2574, W21544, W21545, W10090, W10332, W10087, W11942, W11941, W25034, W25033, W2576, W2575, W21551, W11923, W2573, W2572, W2571, W193, W9040, W2569, W194, W9042, W11936, W25029, W9044, W25027, W21654, W11915, W2532, W2531, W216, W25007, W218, W11914, W2526, W10359, W25006, W9067, W2524, W21651, W2523, W11911, W21644, W9068, W219, W10361, W11909, W11907, W21660, W25003, W21662, W2516, W2515, W21667, W211, W2542, W21610, W11922, W21612, W2541, W10348, W11920, W21615, W21617, W202, W21624, W204, W10349, W2538, W10091, W10352, W11918, W21632, W25010, W2536, W2535, W214, W21637, W21638, W9064, W11916, W10357, W2533, W25063, W175, W11977, W25064, W2658, W2656, W21466, W21467, W21468, W21469, W9007, W11974, W2650, W176, W2649, W2660, W2643, W177, W2640, W10098, W2639, W9011, W178, W2637, W25056, W10097, W180, W25053, W2668, W161, W2676, W8996, W21436, W25076, W164, W11988, W11986, W10105, W2670, W11985, W10101, W8999, W11964, W9002, W2666, W174, W2663, W10318, W21454, W21455, W2662, W25065, W9004, W10099, W21459, W9005, W21524, W9025, W9026, W11953, W185, W2602, W21519, W11952, W2599, W2598, W25038, W2597, W21521, W11951, W2613, W11950, W2591, W9027, W9028, W21534, W9029, W11945, W2586, W11944, W21541, W21542, W21543, W2584, W11957, W21487, W2631, W2630, W2629, W2628, W2625, W2623, W2622, W21494, W11958, W2619, W12088, W2618, W25044, W21504, W2616, W11956, W21509, W25041, W9024, W21511, W2614, W25040, W20885, W25272, W20874, W20876, W3034, W20878, W8823, W20881, W25270, W10170, W12239, W10169, W20883, W20884, W25266, W8818, W3032, W20887, W20888, W20889, W20892, W8825, W42, W3024, W20895, W20896, W8828, W3023, W3055, W8812, W25290, W3062, W20854, W10209, W27, W30, W10177, W25283, W3058, W20859, W12248, W12247, W12235, W12246, W12244, W3050, W3049, W3048, W10175, W10173, W12242, W20869, W3044, W10212, W20870, W3042, W51, W20928, W2994, W2993, W2992, W20931, W25255, W12222, W10230, W20936, W20938, W20939, W2988, W8836, W8844, W2987, W2982, W20940, W12221, W2978, W12219, W12216, W2973, W20951, W12212, W47, W20900, W10221, W8831, W12230, W3018, W3017, W20905, W3016, W10226, W20910, W20911, W3015, W3012, W3010, W8810, W3008, W3006, W10167, W20916, W12226, W20923, W12225, W25256, W8834, W10166, W3103, W20777, W3113, W8, W12282, W3111, W20779, W12281, W9, W11, W12280, W8795, W3105, W8796, W8790, W12278, W10183, W3100, W3099, W12275, W25328, W14, W10197, W25327, W3095, W10182, W25337, W20755, W12293, W20757, W3128, W20758, W12291, W20760, W2, W6, W3127, W8788, W3093, W20764, W20767, W12286, W12285, W20771, W10191, W3117, W12284, W20772, W20775, W10184, W20843, W3078, W3077, W10204, W3074, W12259, W20832, W20833, W22, W3073, W8805, W3071, W20838, W20827, W25297, W20845, W12255, W12254, W3068, W10207, W12252, W25293, W3065, W20847, W20850, W10203, W25323, W12273, W10199, W3090, W20800, W8801, W25314, W8802, W8804, W12211, W25311, W12267, W25308, W20815, W12265, W3083, W12264, W19, W20819, W20824, W2882, W21102, W2881, W82, W21115, W10141, W21120, W8891, W21121, W21122, W21123, W12127, W25201, W12122, W25198, W25197, W2872, W25193, W25192, W12118, W21131, W21132, W21134, W2867, W25189, W10250, W2900, W21073, W12154, W21077, W12153, W21078, W10252, W8874, W10260, W21087, W25211, W21136, W12139, W72, W2889, W25210, W10146, W2886, W25207, W25206, W78, W10266, W21179, W21168, W21169, W21170, W2838, W25178, W21171, W25177, W21173, W21176, W2837, W8904, W8905, W10276, W25175, W12093, W2840, W21180, W10277, W25172, W12091, W21183, W8906, W97, W98, W2830, W2828, W101, W25187, W8896, W12110, W12107, W2862, W21143, W21144, W2861, W2860, W12104, W21152, W12103, W12158, W25186, W25185, W12100, W10272, W8901, W2856, W21157, W21161, W2852, W8902, W12097, W2846, W21006, W2956, W20993, W8854, W25243, W2952, W20995, W2951, W25242, W10235, W12198, W8856, W25241, W10157, W2945, W21007, W2944, W12193, W25240, W10154, W2933, W25239, W21013, W10153, W12188, W20974, W20957, W2971, W2970, W10164, W8846, W20961, W2969, W20962, W20966, W25251, W20970, W8849, W8851, W12185, W2968, W20979, W20980, W2967, W54, W2963, W20985, W25247, W2958, W58, W12204, W10158, W21055, W10247, W25231, W25230, W10249, W12169, W21046, W12167, W2915, W21048, W2914, W2911, W12166, W21042, W12164, W21056, W21057, W67, W68, W21063, W21064, W2907, W12161, W21067, W12160, W8871, W2930, W12183, W21018, W21020, W21021, W21023, W2926, W12179, W21026, W21027, W2923, W21029, W22314, W21031, W12177, W12176, W2922, W10242, W21035, W25235, W10245, W21039, W21041, W10246, W2175, W11775, W2268, W11629, W22136, W11704, W11773, W11630, W10054, W11772, W11626, W2362, W22062, W24923, W2176, W11768, W2360, W11705, W2358, W11767, W22059, W21897, W11621, W11777, W21894, W2368, W352, W9227, W282, W21895, W21896, W11766, W2367, W21898, W24925, W11623, W2216, W11624, W2366, W22200, W24826, W293, W290, W11761, W21920, W2182, W9219, W21923, W24911, W2186, W24910, W21925, W9220, W24837, W21926, W346, W9216, W2274, W2348, W311, W2347, W10396, W287, W11631, W11632, W11764, W21913, W2180, W21914, W24920, W24919, W348, W24868, W21916, W11633, W22055, W2354, W9130, W2272, W22191, W10390, W24940, W9119, W22076, W21859, W11794, W10026, W22219, W21860, W2263, W24818, W2264, W2162, W2386, W359, W266, W2385, W10027, W10435, W267, W9116, W2258, W2156, W10388, W22223, W11696, W360, W10434, W2259, W9117, W9185, W11670, W2262, W10060, W11798, W2218, W11796, W2265, W2166, W22211, W22073, W11618, W22071, W22070, W2266, W21883, W10057, W21881, W22066, W10056, W22065, W11619, W2375, W24927, W2374, W22215, W11788, W21870, W2383, W21872, W268, W271, W11639, W10058, W357, W2163, W21877, W2381, W24933, W11781, W11780, W2378, W22009, W22048, W2199, W11734, W11733, W22004, W10034, W2283, W24880, W2201, W2310, W11664, W11729, W9201, W11728, W22147, W22150, W22151, W21998, W21990, W298, W24885, W2282, W9145, W21995, W2321, W21996, W10412, W10409, W2320, W21999, W300, W2319, W2318, W24882, W9203, W2317, W301, W302, W22026, W22027, W22028, W2298, W11724, W22032, W9163, W22023, W2297, W2208, W2209, W304, W22153, W11719, W2292, W2210, W2294, W2305, W11667, W9149, W2303, W2302, W22045, W9166, W2212, W2203, W24847, W21989, W22159, W2300, W11716, W2289, W9199, W10413, W2299, W2211, W21953, W11753, W21947, W2340, W10404, W2339, W21951, W11752, W22144, W11714, W2343, W9209, W11749, W21957, W21960, W22179, W10033, W11747, W22177, W21937, W21931, W345, W11711, W2346, W22184, W11759, W22183, W21935, W2345, W11743, W11713, W22143, W21938, W10048, W9213, W11757, W332, W10399, W9136, W9212, W10416, W24893, W2196, W297, W21980, W22165, W9206, W9142, W2279, W24892, W22050, W21977, W342, W24891, W21985, W11738, W2323, W24890, W22162, W21673, W24888, W9168, W21965, W22052, W11650, W24839, W11742, W11741, W11654, W9141, W2158, W21971, W11655, W24894, W22171, W21972, W2328, W343, W24869, W2327, W2112, W21730, W10077, W9194, W22102, W24800, W21731, W24982, W22101, W24981, W21734, W373, W2108, W2116, W21735, W2480, W22099, W22098, W11597, W24979, W24859, W11892, W2119, W2245, W9256, W21719, W22291, W228, W22122, W2483, W21723, W2244, W11896, W10373, W24794, W2107, W21725, W21726, W21727, W2481, W24797, W22288, W21729, W2247, W2228, W10378, W11885, W2125, W2463, W11883, W2460, W21762, W21763, W10379, W2466, W2458, W9189, W9081, W24974, W22273, W22271, W21767, W21768, W2472, W2477, W22124, W2476, W10377, W9249, W235, W22277, W21748, W2484, W10074, W11889, W21752, W2469, W2468, W2467, W22275, W9190, W11586, W2238, W22308, W11686, W2508, W2239, W2507, W24790, W2087, W2505, W24996, W2241, W11901, W9073, W24791, W21696, W2088, W21697, W2084, W327, W2511, W9193, W10446, W21675, W21676, W21677, W11581, W2504, W21681, W25000, W9262, W11902, W21684, W2085, W2086, W2509, W21689, W21693, W2494, W2099, W21705, W21708, W22296, W21709, W22295, W2499, W2498, W21714, W9077, W21704, W11684, W11899, W10368, W2492, W2491, W2490, W22104, W10078, W2103, W2090, W2502, W21699, W22301, W2089, W2501, W225, W22300, W2500, W9084, W22106, W11688, W10079, W2094, W11685, W9075, W9259, W328, W21703, W10429, W9107, W22244, W2414, W9109, W10386, W251, W2254, W9195, W9239, W24951, W22242, W11836, W21832, W22239, W2227, W9238, W22238, W24809, W252, W2409, W10067, W21834, W11842, W11608, W22248, W249, W11844, W250, W22129, W22247, W2422, W24811, W2421, W9105, W21817, W2142, W11838, W21822, W21824, W21826, W2400, W21844, W254, W2256, W22232, W22133, W2401, W22083, W2152, W11672, W2399, W24815, W21850, W10423, W11611, W22227, W21851, W2398, W11674, W11691, W22131, W11823, W367, W24812, W24862, W2147, W9235, W22127, W22085, W2148, W253, W11610, W11820, W11816, W2402, W11815, W11814, W24805, W22264, W2449, W10382, W9089, W2447, W11859, W24965, W22263, W239, W11861, W2131, W21785, W10071, W370, W22089, W10383, W9093, W11854, W11599, W2453, W10441, W24803, W238, W10380, W21769, W22092, W11868, W21772, W241, W371, W22091, W11600, W21774, W11865, W10381, W11602, W2130, W321, W21797, W11604, W2433, W21793, W2441, W9094, W2136, W11605, W24959, W21796, W2135, W22252, W11851, W22251, W21799, W24958, W9188, W11850, W11848, W11847, W245, W10385, W244, W2438, W2440, W21789, W22259, W24807, W24961, W2133, W43882, W10159, W40902, W10155, W40712, W7396, W7389, W7006, W41036, W9869, W7174, W7395, W9874, W9870, W41069, W7423, W10180, W9832, W10023, W9831, W10179, W10014, W7425, W10181, W40881, W7199, W10178, W9835, W7418, W7203, W7419, W6993, W9834, W10011, W43477, W9833, W7422, W6992, W40704, W7430, W43914, W7429, W10022, W7187, W7188, W10020, W7190, W10185, W10187, W40875, W7196, W43910, W40696, W40871, W10017, W7195, W7194, W10031, W7001, W7213, W9853, W7000, W7405, W43488, W6999, W40720, W43896, W10001, W10035, W7216, W7177, W43886, W7004, W9867, W9849, W7178, W9864, W7399, W9858, W9845, W10133, W41058, W40709, W7184, W40864, W43482, W10176, W43709, W43903, W7417, W6994, W10009, W6997, W7180, W7209, W40718, W10030, W10029, W43685, W7412, W7206, W10028, W7204, W43898, W6996, W10171, W10172, W7323, W7127, W40991, W10100, W10104, W7066, W10108, W7128, W7126, W7064, W10109, W10111, W7063, W7130, W10113, W7271, W7268, W7117, W43579, W40789, W40788, W10095, W40785, W7279, W7328, W7121, W40988, W7319, W7274, W7321, W9926, W7322, W40936, W7335, W10062, W40995, W10117, W7337, W7058, W7258, W40938, W43831, W40768, W9922, W7251, W7138, W7249, W43644, W43835, W9918, W7263, W7061, W10065, W7330, W43633, W7265, W7132, W9965, W43566, W9966, W7331, W43638, W9968, W7092, W40805, W43611, W9952, W40956, W7295, W10080, W7101, W7089, W43801, W7284, W7088, W9939, W43604, W9949, W9943, W7095, W7094, W43793, W9950, W7294, W40799, W40806, W9951, W7098, W9942, W7289, W9940, W7282, W7079, W9935, W9961, W10092, W10093, W7077, W7080, W7310, W7110, W7281, W7076, W9932, W7299, W10084, W7086, W7085, W43807, W7102, W40976, W43592, W7300, W7301, W7304, W43587, W7107, W7108, W7082, W7373, W41024, W7230, W7170, W9985, W9986, W10140, W10042, W40844, W7021, W9991, W40845, W7369, W10134, W7233, W9981, W10043, W10136, W41021, W9889, W10137, W10148, W10138, W9983, W7371, W43526, W7372, W7384, W7378, W10039, W10151, W7013, W7220, W7383, W7377, W9996, W7011, W7387, W10152, W7388, W10037, W7010, W7015, W43726, W7172, W43518, W40740, W10041, W7225, W43516, W10150, W7173, W41030, W9994, W43722, W9995, W9879, W7044, W7350, W10055, W7151, W40934, W40826, W9903, W40932, W7045, W7154, W10127, W43742, W10053, W9900, W7351, W40759, W9898, W7353, W7144, W9915, W7145, W40822, W9914, W7338, W7247, W10118, W7050, W7048, W7148, W7344, W10126, W7245, W43746, W7345, W9909, W7046, W9907, W43842, W9892, W10047, W10046, W10045, W7360, W9894, W7238, W7358, W7164, W7030, W7237, W7367, W7165, W9978, W7235, W9980, W10050, W7354, W7036, W7240, W7355, W43541, W7159, W10049, W41015, W7357, W7035, W10131, W41792, W9120, W9122, W42570, W41788, W8319, W8330, W8317, W8311, W41784, W42580, W8306, W9111, W9100, W9101, W9102, W9104, W41808, W8338, W9123, W9113, W9139, W8286, W9140, W8278, W9143, W9144, W8276, W42629, W8275, W8271, W8266, W9129, W8303, W41780, W42594, W9125, W42595, W9127, W8299, W8298, W8296, W9131, W9132, W42602, W9133, W9135, W42606, W9069, W42478, W41855, W8411, W9063, W9066, W41851, W41856, W9070, W9071, W8399, W8398, W8397, W8394, W8416, W9045, W8424, W9047, W41866, W9048, W9049, W8419, W8418, W41861, W8393, W9056, W42470, W9058, W8414, W9060, W8413, W8361, W42527, W9085, W8367, W42529, W41828, W41827, W9086, W8369, W9090, W42540, W9092, W8357, W42542, W8350, W9097, W8384, W9076, W9078, W42508, W8390, W8388, W8387, W8265, W8383, W41839, W42518, W42521, W9079, W41833, W9274, W8135, W8134, W9265, W9266, W8131, W9269, W9273, W9263, W8130, W9275, W9276, W8125, W8123, W8122, W9253, W8169, W9243, W8166, W8165, W8163, W9245, W9246, W8157, W9251, W9252, W8154, W8151, W9258, W8147, W42745, W9260, W8142, W9321, W8098, W8096, W9309, W9311, W9317, W8091, W41620, W8084, W42788, W41616, W8081, W9323, W8075, W9329, W8072, W9295, W9280, W9281, W42771, W41647, W9283, W9285, W42772, W41643, W9290, W8114, W9242, W9297, W9300, W8108, W9301, W42783, W9302, W8224, W8241, W8239, W9187, W42658, W8235, W8234, W9184, W9192, W8220, W9197, W9165, W8256, W8255, W9152, W9153, W8254, W9157, W9159, W42681, W8248, W42648, W9171, W8246, W9176, W9179, W9182, W9183, W9225, W8186, W9229, W9231, W8181, W9233, W9222, W9234, W8178, W42719, W8177, W9241, W9207, W9200, W9202, W8202, W9204, W8201, W42693, W8198, W9211, W9217, W9218, W41698, W8190, W8660, W8853, W42245, W8855, W8651, W42251, W8860, W8661, W8644, W8642, W8862, W8863, W8638, W8634, W8865, W8866, W8867, W8668, W8682, W8835, W8840, W8843, W8676, W8675, W8674, W8672, W42044, W8847, W8848, W42237, W42065, W8852, W42063, W8664, W8889, W8604, W8600, W8882, W8883, W8886, W8893, W8894, W8897, W8868, W42042, W8624, W8623, W42273, W8620, W8869, W42276, W8872, W8873, W8875, W8876, W8879, W8881, W8607, W8744, W8753, W8751, W8750, W8799, W42156, W42111, W8800, W8745, W42106, W8742, W8741, W8740, W8806, W8807, W8734, W8733, W8770, W8785, W8786, W8779, W8777, W8775, W8773, W8789, W8769, W8791, W8792, W8762, W8759, W8756, W42147, W42150, W8697, W42089, W42198, W42199, W8708, W8707, W42206, W8710, W8696, W8830, W8832, W42080, W8685, W8723, W8730, W42177, W42180, W8725, W8813, W8724, W8593, W8814, W8722, W8815, W42094, W8719, W8816, W8716, W8820, W8481, W8994, W8478, W42404, W8476, W8995, W8997, W8998, W8475, W8474, W8472, W8471, W9003, W8979, W8500, W8980, W8982, W8499, W8496, W8984, W8494, W42419, W8492, W8489, W8986, W8988, W8991, W8443, W8436, W9030, W9031, W9033, W9035, W8445, W8431, W42452, W9036, W9041, W42453, W42454, W9043, W8429, W41870, W9006, W8461, W9008, W9009, W9010, W8454, W8976, W9016, W41894, W9017, W9018, W42431, W8448, W8446, W8927, W8910, W8912, W42322, W45809, W41990, W42327, W41986, W42320, W8928, W8563, W8929, W8562, W41976, W8558, W8555, W8553, W8900, W8592, W42006, W8590, W42305, W8587, W8903, W42311, W8552, W8577, W41998, W8907, W8909, W8516, W8958, W42359, W8959, W8529, W8963, W42362, W42363, W8964, W42366, W42367, W42369, W8531, W8512, W8511, W8509, W8968, W8969, W8970, W8972, W8974, W8975, W8505, W8539, W8935, W8547, W8939, W42346, W8542, W8940, W8941, W8942, W8945, W8535, W42354, W8948, W8951, W8954, W9692, W9693, W7630, W7631, W9700, W41221, W7627, W9704, W7626, W7625, W7623, W9673, W7658, W7657, W7655, W41248, W7651, W7650, W7649, W41210, W9674, W9676, W41242, W41241, W9677, W9682, W43251, W7641, W7637, W7636, W41194, W9726, W7596, W7593, W43311, W41196, W7587, W9730, W41193, W7586, W9731, W9733, W41190, W41189, W7581, W9734, W41187, W7579, W7622, W9715, W7617, W9716, W9717, W7613, W7612, W7660, W7609, W9722, W43291, W7605, W7604, W41201, W7719, W7717, W9622, W43178, W41300, W9625, W7712, W9627, W7711, W41284, W9629, W7706, W41281, W41316, W9605, W41314, W7735, W7732, W9631, W7729, W7727, W9607, W9610, W41305, W7725, W41302, W43221, W9651, W9652, W7687, W7681, W9657, W41256, W7677, W9663, W9666, W7672, W41251, W7670, W7668, W7667, W41279, W7705, W41278, W9632, W9636, W41273, W9641, W9644, W41186, W9646, W43200, W7692, W9649, W7690, W9799, W41110, W7495, W7493, W7491, W41106, W7496, W7483, W41104, W7480, W43417, W9800, W7476, W7475, W9784, W9785, W9787, W7510, W7507, W9792, W43394, W7474, W7504, W7503, W7501, W7500, W9793, W9795, W7497, W7451, W9815, W7449, W43448, W7447, W7446, W9816, W7444, W9819, W7441, W7439, W41076, W43432, W9805, W9806, W7473, W7472, W7471, W7470, W7467, W41095, W43431, W9783, W9811, W7464, W7463, W41091, W9812, W7456, W41171, W41170, W7556, W7555, W7554, W7553, W7552, W9749, W41164, W43344, W7558, W9751, W7548, W41160, W7547, W43352, W7544, W7569, W41185, W9736, W41182, W7574, W7571, W9739, W9740, W9741, W9759, W9742, W7567, W9744, W7565, W7564, W7562, W7561, W9764, W9765, W9766, W7524, W7520, W7525, W9772, W7516, W9773, W9774, W43386, W9780, W43389, W9782, W41127, W7543, W7542, W41152, W7539, W7537, W9761, W7536, W9602, W43365, W7533, W7532, W43369, W7530, W7528, W9763, W7526, W41517, W7976, W42918, W7974, W42921, W9411, W9408, W9421, W7965, W9422, W9394, W8000, W9386, W42895, W9387, W9391, W42898, W9393, W7992, W7961, W9398, W7986, W9403, W9404, W41526, W7979, W7924, W7936, W9440, W7934, W7933, W41485, W7931, W7928, W7926, W7923, W9456, W41478, W9457, W9459, W42950, W9424, W7959, W7954, W42945, W41499, W7944, W9434, W8001, W7942, W7940, W9436, W9438, W41492, W9439, W8041, W42833, W9344, W8048, W8047, W42841, W8045, W8044, W9346, W8042, W9347, W9349, W42847, W8039, W9350, W9351, W8038, W9353, W9354, W9330, W9331, W9333, W8068, W41601, W9335, W8035, W8065, W9336, W9339, W8061, W8060, W8054, W9342, W42831, W8009, W8016, W41565, W8015, W9368, W9369, W8011, W9370, W9371, W9372, W8008, W8007, W9375, W9377, W9382, W8002, W42889, W8029, W8034, W42854, W8032, W9355, W42860, W41575, W9357, W42862, W7922, W41573, W8025, W9359, W9362, W9364, W42869, W8023, W8022, W8019, W41370, W7806, W7803, W41365, W7801, W7798, W7807, W41359, W7796, W43094, W43095, W7795, W7794, W9566, W41356, W9540, W9541, W7828, W9546, W7827, W43062, W7826, W9547, W9549, W9555, W7815, W9556, W7808, W41329, W9588, W7760, W7758, W7757, W43136, W9589, W9590, W9593, W9587, W7754, W9595, W9597, W7750, W9598, W7744, W7741, W43120, W43110, W41350, W41349, W43113, W9574, W7772, W43117, W7771, W7768, W9533, W7766, W9577, W9578, W41343, W9580, W9583, W7762, W43128, W9475, W41452, W42999, W41450, W7890, W7887, W43004, W41446, W41456, W9487, W7874, W9491, W43012, W7872, W9492, W9493, W7871, W7869, W7867, W9461, W7916, W9462, W7912, W7908, W7907, W9470, W41465, W7906, W9472, W7905, W7903, W42993, W7900, W9474, W9519, W9513, W7843, W7842, W7841, W7839, W7838, W7844, W41401, W9522, W7833, W7832, W9526, W9527, W7830, W41392, W9503, W7866, W7862, W7859, W9496, W7854, W7853, W9823, W41422, W9505, W43033, W7847, W9510, W2349, W2350, W2351, W2353, W2355, W2356, W2361, W2363, W2364, W2365, W2369, W2329, W2330, W48663, W2331, W2333, W2334, W2335, W2376, W2336, W2337, W2341, W2391, W2392, W2393, W2396, W2403, W2405, W48569, W2407, W2411, W2412, W48600, W2380, W2382, W2384, W2387, W2389, W2253, W2229, W2230, W2233, W2237, W2243, W2252, W2255, W2260, W2267, W2219, W2200, W2202, W2205, W2206, W2207, W2217, W2220, W2224, W2314, W2301, W2304, W2309, W2311, W2313, W2322, W2324, W2326, W2281, W48727, W2270, W2271, W2275, W2277, W2285, W2286, W2291, W2296, W48705, W2559, W2560, W2564, W2565, W2566, W2567, W2577, W2578, W2579, W48389, W2580, W2582, W48437, W2539, W2540, W2583, W2544, W2545, W2548, W2558, W2635, W2633, W2634, W2620, W2638, W2641, W2648, W2653, W2596, W2585, W2587, W2589, W2593, W2595, W2601, W2606, W2611, W2612, W2615, W2617, W48541, W2444, W48535, W2446, W2450, W2432, W2451, W48523, W2452, W2454, W2418, W2419, W2420, W48558, W48556, W48554, W2424, W2427, W2455, W2428, W2429, W48545, W2430, W2431, W2519, W2512, W2513, W2518, W48478, W2520, W2525, W2528, W2534, W2456, W2462, W2465, W2473, W2479, W2482, W2485, W2493, W2496, W49078, W1902, W1905, W1907, W1912, W1898, W1915, W1927, W1931, W1933, W1934, W1865, W1867, W1870, W1874, W1937, W1883, W1885, W1890, W1891, W1893, W1959, W1962, W1963, W1965, W1968, W1970, W49018, W1980, W1947, W1938, W1939, W1940, W1942, W1946, W1862, W1950, W1952, W1955, W49037, W1799, W1792, W1793, W1796, W1797, W1798, W1791, W1801, W1783, W1773, W49220, W1780, W1781, W1786, W1788, W1789, W1790, W1835, W1839, W1847, W1853, W49133, W1856, W1860, W1820, W1805, W1812, W1813, W1814, W1825, W1826, W1827, W1832, W2153, W2134, W2137, W2140, W2143, W2146, W2150, W2157, W2160, W2118, W2091, W2097, W2101, W2109, W2165, W2120, W2124, W2128, W2129, W48872, W2190, W2183, W2187, W2188, W2192, W2193, W2194, W2195, W2197, W2198, W48828, W2167, W2170, W2171, W2172, W2173, W2178, W48818, W2181, W2023, W2009, W2014, W2019, W2021, W2024, W2028, W2030, W2033, W2038, W1984, W1985, W1989, W1993, W2039, W1995, W1998, W2004, W2062, W2063, W2064, W2065, W2066, W2068, W2069, W2070, W2071, W2072, W2080, W2083, W2052, W2042, W2044, W2045, W2046, W2048, W2050, W2659, W2054, W2057, W2058, W2059, W3202, W47758, W3203, W3209, W47787, W3178, W3186, W3189, W3194, W3198, W3199, W3200, W3201, W3265, W3250, W3252, W3257, W3259, W3244, W3274, W3276, W3277, W3279, W3238, W3229, W3232, W3234, W3235, W3176, W3239, W3240, W3242, W3243, W3115, W3116, W3120, W3121, W3126, W47853, W3112, W3130, W3132, W3089, W3091, W47886, W47884, W3092, W3096, W3098, W3136, W3101, W3109, W3110, W3171, W3163, W3164, W3166, W3168, W3173, W3174, W3137, W3141, W3149, W3151, W3153, W3154, W3156, W3157, W47518, W3439, W3442, W3443, W3446, W3452, W3455, W3458, W3464, W3468, W47504, W47501, W3406, W3408, W3410, W3413, W3415, W3419, W3477, W47547, W3426, W3438, W3506, W3500, W3501, W3502, W3504, W3498, W3508, W3511, W3514, W3516, W3519, W3478, W3480, W3405, W3495, W3497, W3334, W3314, W3316, W3327, W47632, W3311, W3336, W3339, W3340, W47624, W3344, W3350, W47675, W3282, W3283, W3284, W3288, W3291, W3292, W3293, W3352, W3295, W3297, W3299, W3303, W3306, W3307, W3388, W3380, W3381, W3385, W3376, W3390, W3392, W3396, W3398, W3400, W3403, W3354, W3356, W3357, W3358, W3359, W3364, W3365, W3375, W2791, W2778, W2781, W2783, W2784, W2785, W48181, W2792, W2797, W2801, W2806, W2807, W2768, W2763, W2764, W2767, W48207, W2769, W2772, W2773, W2774, W2775, W2835, W2836, W2849, W2850, W2854, W2858, W2834, W2859, W2863, W2823, W2815, W2817, W2818, W2822, W2831, W2833, W48136, W2686, W2687, W2696, W2697, W2698, W2699, W2700, W2703, W2706, W2672, W2664, W2667, W2669, W2708, W2673, W2675, W2680, W2685, W48231, W2733, W48235, W2744, W2748, W2755, W2759, W2760, W2725, W2711, W2713, W2716, W2722, W2723, W2865, W2726, W2728, W2729, W2730, W3005, W2990, W2991, W2995, W2996, W2998, W47968, W3001, W3002, W2989, W3019, W3021, W2957, W2959, W2962, W2965, W47994, W2972, W2975, W2977, W2979, W3061, W3063, W3064, W3067, W3070, W3082, W3084, W3085, W3087, W3088, W3045, W3030, W3033, W3037, W3038, W3046, W3051, W2897, W2887, W2890, W2891, W2892, W2893, W2895, W2896, W2899, W2902, W2904, W2906, W2877, W2869, W2871, W2875, W2879, W2883, W2885, W2946, W2929, W2931, W2932, W2936, W2937, W2940, W2942, W2947, W2948, W2953, W2954, W2918, W2909, W2916, W2917, W1771, W2919, W2921, W2924, W618, W601, W602, W603, W611, W613, W50410, W620, W624, W628, W591, W577, W584, W592, W595, W679, W663, W667, W674, W675, W657, W681, W684, W685, W634, W637, W639, W642, W645, W568, W647, W648, W654, W655, W656, W485, W477, W479, W480, W489, W492, W498, W503, W449, W434, W441, W445, W448, W504, W465, W467, W474, W475, W548, W535, W538, W540, W541, W542, W546, W531, W549, W550, W554, W562, W519, W508, W511, W517, W518, W689, W528, W530, W817, W820, W821, W822, W827, W830, W815, W836, W841, W845, W846, W800, W791, W793, W797, W849, W802, W803, W806, W807, W811, W812, W813, W895, W883, W885, W890, W892, W893, W50105, W894, W882, W898, W902, W908, W910, W852, W856, W860, W861, W867, W790, W870, W872, W878, W716, W708, W721, W725, W691, W693, W734, W698, W702, W706, W771, W760, W762, W763, W768, W769, W774, W775, W777, W779, W783, W743, W739, W740, W742, W749, W755, W757, W758, W139, W125, W132, W136, W137, W140, W143, W91, W79, W83, W86, W88, W147, W93, W94, W99, W100, W102, W105, W184, W186, W188, W189, W190, W191, W197, W198, W199, W201, W153, W155, W160, W162, W163, W166, W50909, W170, W171, W172, W179, W181, W34, W26, W29, W31, W33, W36, W38, W41, W43, W0, W7, W12, W44, W16, W17, W18, W20, W23, W62, W63, W64, W65, W66, W69, W70, W71, W74, W77, W53, W46, W48, W49, W50, W52, W205, W59, W374, W366, W369, W358, W50627, W375, W378, W380, W325, W326, W331, W333, W381, W344, W349, W351, W354, W402, W403, W411, W417, W418, W420, W422, W423, W425, W427, W432, W433, W397, W384, W387, W391, W394, W322, W400, W401, W248, W236, W243, W232, W256, W257, W261, W224, W209, W212, W213, W264, W226, W230, W305, W50698, W299, W308, W313, W272, W276, W280, W284, W285, W286, W911, W288, W292, W294, W295, W296, W1490, W1491, W1494, W1489, W1505, W1506, W1509, W1510, W1464, W1467, W1471, W1473, W1475, W1511, W49528, W1479, W1481, W1482, W1533, W1538, W1542, W1544, W1530, W1545, W1546, W1550, W1551, W1512, W1513, W1514, W1516, W1517, W1521, W1522, W1524, W1526, W1528, W1401, W1388, W1390, W1391, W1392, W1398, W49615, W1403, W1405, W1411, W1384, W1373, W1374, W1376, W1379, W1383, W1385, W1386, W49624, W1451, W1443, W1444, W1445, W1448, W1454, W1459, W49549, W1462, W1423, W1414, W1419, W1420, W1422, W1424, W1428, W1431, W1432, W1696, W1697, W1698, W1704, W1695, W49293, W1705, W1707, W1709, W1710, W1715, W1676, W1660, W1661, W1670, W1672, W1683, W1686, W1687, W1689, W1694, W1737, W1739, W1747, W1736, W1750, W1755, W1756, W1764, W1766, W1726, W1719, W1720, W1721, W1722, W1723, W1728, W1730, W49262, W1583, W1584, W1587, W1588, W1590, W1592, W1579, W1594, W1595, W1558, W1561, W1563, W1567, W1597, W1570, W1572, W1573, W1574, W1575, W1576, W49362, W1637, W1640, W1644, W1646, W49353, W1647, W1653, W1654, W1655, W1656, W1657, W1600, W1604, W1605, W1606, W1611, W1613, W1371, W1616, W1620, W1625, W1626, W1627, W1629, W1631, W1064, W49942, W1067, W1069, W1071, W1072, W1076, W1077, W1078, W1040, W1042, W1043, W1046, W1055, W1080, W1057, W1058, W1062, W1115, W1122, W1126, W1128, W1106, W1134, W1136, W1137, W1141, W1144, W1092, W1081, W1082, W1084, W1086, W1087, W1094, W1095, W1096, W1100, W945, W948, W949, W952, W964, W942, W973, W975, W980, W927, W913, W914, W916, W922, W924, W983, W928, W933, W934, W935, W939, W1017, W1018, W1019, W1022, W1025, W1026, W1010, W1028, W49987, W1030, W1032, W1036, W997, W985, W986, W994, W1147, W999, W1001, W1004, W1008, W1292, W1277, W1286, W1289, W1290, W1291, W1276, W1293, W1296, W1298, W1299, W1300, W1251, W1238, W1239, W1240, W1243, W1245, W1249, W1250, W1258, W1270, W1275, W1358, W1331, W1334, W1343, W1346, W1351, W1328, W1361, W1362, W1363, W1365, W1369, W1309, W1302, W1303, W1312, W1313, W1314, W1315, W1324, W1326, W1187, W1176, W1179, W1180, W1185, W1193, W1196, W1197, W1200, W1151, W1155, W1157, W1203, W1164, W1167, W1169, W1172, W1228, W1216, W1218, W1220, W1225, W1215, W1233, W1234, W1205, W1207, W1208, W3523, W1210, W1212, W1213, W1214, W5787, W5772, W5774, W5775, W5776, W5779, W5780, W5783, W5764, W5790, W5795, W5799, W5809, W45179, W5736, W5738, W5751, W5810, W5753, W5754, W45165, W5755, W5756, W5759, W5860, W5848, W5849, W5850, W5853, W5855, W5857, W5842, W45075, W5865, W45068, W5822, W5814, W5817, W45111, W5830, W5832, W5838, W5650, W45269, W45267, W45264, W5654, W5658, W5659, W5649, W45255, W5667, W45251, W5669, W45237, W5622, W5624, W5625, W5627, W5629, W5683, W5631, W5633, W5634, W5640, W5644, W5645, W5648, W5719, W5712, W45205, W5713, W5718, W45209, W5721, W5723, W5725, W5726, W5727, W5728, W5729, W5685, W5686, W5687, W45225, W5694, W5695, W5699, W5700, W45211, W6031, W6014, W6016, W6017, W6020, W6024, W6032, W6033, W44901, W6037, W6038, W6042, W6043, W5978, W5968, W44950, W5971, W5972, W5974, W5977, W6044, W5999, W6002, W6003, W6004, W6007, W6065, W44862, W44861, W6066, W6069, W6070, W6071, W6072, W6074, W44864, W6075, W6076, W6081, W6088, W6093, W44836, W6051, W5965, W6058, W44868, W6063, W5903, W5896, W5898, W5899, W5892, W5907, W5909, W45018, W5911, W5912, W5877, W5871, W5874, W5878, W5887, W5888, W5889, W5959, W5950, W44974, W5953, W5945, W5960, W5962, W5932, W5916, W5918, W5920, W5925, W44999, W5934, W5936, W5938, W5940, W5941, W5942, W5348, W5336, W5337, W45595, W5340, W5344, W5350, W5354, W5355, W5361, W5322, W5309, W5310, W5311, W5312, W5315, W5331, W45606, W5333, W5335, W5396, W5398, W45533, W5404, W5407, W45525, W5408, W5410, W5411, W45559, W45574, W5363, W5368, W45564, W45558, W5378, W5379, W5383, W5387, W5238, W5230, W5233, W5237, W45710, W5239, W45693, W45692, W5241, W5243, W5219, W45732, W5215, W45728, W45726, W5218, W5222, W5223, W5224, W5225, W45714, W5227, W5299, W5286, W5297, W5298, W5300, W5304, W5305, W5259, W5244, W5248, W5250, W5251, W5252, W45679, W45678, W5412, W5263, W5266, W5270, W5272, W5276, W5277, W5554, W45373, W5539, W5545, W5551, W5552, W5555, W5556, W5557, W5506, W5508, W5510, W5517, W5560, W5523, W5524, W5528, W5531, W5533, W5600, W5581, W5583, W5588, W5594, W5597, W5579, W5604, W5605, W5610, W5611, W5614, W5616, W5567, W5563, W45349, W5565, W5502, W5572, W5573, W45337, W5576, W5577, W5439, W5440, W5444, W5447, W5448, W5433, W5450, W5451, W5453, W5457, W5458, W5419, W45517, W5416, W5417, W5418, W5460, W5420, W5425, W5426, W5429, W5431, W5494, W5488, W5492, W45429, W45426, W5486, W5497, W5498, W5500, W45413, W5468, W45463, W5461, W5465, W5466, W6096, W5477, W5479, W5481, W5482, W6692, W6682, W6684, W44226, W6686, W6688, W6690, W6691, W6681, W6698, W6700, W44209, W6702, W6675, W44249, W6671, W44246, W6673, W6674, W44241, W44239, W6680, W6743, W6740, W44167, W6741, W6744, W44159, W6751, W44154, W44153, W6754, W6720, W6706, W6712, W6715, W6716, W44190, W6721, W44183, W6726, W6607, W6609, W6610, W6611, W6612, W6613, W6620, W6587, W6579, W44348, W6581, W6583, W6584, W6585, W6588, W6591, W6593, W6596, W6598, W6599, W6663, W6658, W6662, W6656, W6664, W6665, W44261, W6667, W6670, W6631, W6639, W44296, W44293, W44292, W6755, W6645, W6648, W6650, W6655, W6922, W6909, W6913, W6916, W43992, W6921, W6925, W6926, W6928, W6929, W6931, W6932, W6872, W6876, W6885, W44024, W44023, W43976, W6896, W6898, W6900, W6902, W6906, W44004, W6967, W43947, W6960, W6966, W6968, W6972, W6976, W6977, W6933, W6937, W6942, W6943, W6944, W6950, W6871, W6951, W43958, W6955, W6956, W43950, W44120, W6790, W6793, W6787, W6799, W6807, W6808, W6810, W6811, W6770, W6758, W6759, W6761, W6762, W44139, W6812, W6771, W6774, W44132, W6776, W6777, W6778, W6786, W6846, W6835, W6837, W44064, W6839, W6833, W6849, W6858, W6860, W6828, W6815, W6819, W6820, W6822, W6823, W6826, W6827, W44077, W44075, W6832, W6251, W44682, W6244, W44680, W6248, W6250, W6242, W6252, W44668, W6258, W6227, W6203, W6210, W6216, W6220, W6259, W44698, W6228, W44694, W6233, W6238, W6240, W6279, W6285, W6287, W6294, W6296, W6298, W6278, W6301, W6302, W6304, W6305, W44603, W6311, W6312, W6268, W44655, W6260, W6266, W44647, W44646, W44645, W6270, W6272, W6273, W6133, W6120, W6126, W6131, W6116, W6134, W6137, W6142, W6151, W6154, W6156, W6109, W6100, W6101, W6103, W44824, W6106, W6159, W6110, W44816, W6111, W6113, W44812, W6195, W44735, W6201, W6202, W44763, W6164, W6167, W6170, W6172, W6313, W44762, W6177, W6182, W6187, W6481, W44441, W6484, W6488, W6490, W6480, W6491, W6497, W6499, W6458, W6442, W44474, W6445, W6446, W6448, W6451, W6452, W6454, W6467, W6476, W6526, W6527, W44384, W6536, W6540, W6552, W6555, W6524, W6566, W6567, W44359, W6570, W6501, W6509, W6515, W6517, W6519, W6520, W6365, W6351, W44561, W6352, W6356, W6358, W6364, W6367, W6369, W44545, W6371, W6334, W44590, W6326, W6330, W44581, W6333, W6372, W6336, W6339, W6341, W6343, W6344, W6414, W6405, W6407, W6409, W44504, W6401, W6422, W6430, W44486, W6433, W6388, W6373, W6374, W6381, W44531, W5211, W6389, W6397, W6399, W4083, W4086, W4087, W4088, W4092, W4096, W4097, W4102, W4106, W4109, W46867, W4112, W4114, W4115, W4053, W46914, W4060, W4061, W4064, W4071, W4116, W4075, W4079, W4080, W4082, W4144, W4147, W4148, W4150, W4154, W4158, W4142, W4166, W46814, W4169, W4170, W4171, W4172, W4125, W46860, W46858, W4117, W4118, W46852, W4052, W4126, W4132, W46841, W4136, W46836, W4139, W3987, W3980, W3982, W3983, W3985, W3986, W3988, W3991, W3993, W3996, W3998, W4000, W47010, W3958, W3959, W4001, W47008, W3963, W3966, W3967, W3970, W3971, W3973, W4030, W4017, W4019, W4020, W4022, W4024, W4015, W4039, W4040, W4041, W4043, W4045, W4049, W4051, W4002, W4004, W46968, W4005, W4006, W4009, W4010, W4011, W4340, W4330, W4336, W46660, W4325, W4351, W4352, W4355, W4297, W4300, W4306, W4310, W46686, W4357, W4311, W4312, W46681, W4317, W4320, W4322, W4405, W4406, W4407, W4411, W4401, W4416, W4417, W4418, W4419, W4425, W4426, W4378, W4358, W4360, W4362, W4365, W4368, W4373, W4375, W4296, W4389, W46617, W4396, W4398, W4399, W4210, W4211, W46776, W4213, W4215, W4216, W46769, W4221, W4224, W4229, W4231, W4235, W4237, W4238, W4239, W4204, W4184, W4185, W4186, W4187, W4190, W4198, W4199, W4274, W4262, W4263, W4266, W4267, W4271, W4272, W4273, W46709, W46708, W4279, W4291, W4295, W46754, W4240, W4241, W4243, W4249, W4250, W4254, W4255, W3675, W3665, W3668, W3669, W47309, W47308, W3670, W3672, W3657, W3676, W47296, W3678, W3637, W3641, W3648, W3679, W3649, W3650, W3656, W3719, W3705, W3706, W3713, W3720, W3726, W3729, W3680, W3681, W3682, W3683, W3685, W47287, W3687, W3689, W3631, W3690, W3691, W3692, W3698, W3702, W3573, W3563, W3564, W3570, W3572, W3562, W3579, W3580, W3586, W3545, W3526, W3533, W3534, W3540, W3542, W3543, W3548, W3551, W3554, W3557, W3561, W3620, W3609, W3611, W3612, W3618, W3624, W3626, W3627, W3628, W47381, W47388, W47385, W47384, W3593, W3597, W3598, W3599, W3601, W3603, W3606, W3863, W3851, W47105, W3854, W3855, W3862, W3865, W3871, W47090, W3872, W3874, W3883, W3884, W3835, W3837, W3839, W3840, W47122, W47120, W3891, W47117, W3845, W3846, W3847, W3925, W3913, W3918, W3919, W3922, W3931, W3932, W3933, W3935, W3940, W3944, W47027, W3898, W3892, W3893, W3896, W3833, W3899, W3900, W3905, W3908, W47057, W3910, W3773, W3761, W3764, W3771, W47195, W3760, W3774, W3775, W3781, W3782, W3750, W3730, W3732, W3733, W3736, W3740, W3745, W47227, W3786, W3751, W3754, W47216, W3757, W3820, W3822, W47145, W3827, W3829, W3831, W3832, W3804, W3787, W3790, W3801, W3802, W3803, W46582, W3805, W3807, W3808, W3810, W3814, W4950, W4951, W46030, W46029, W4952, W46025, W4948, W4963, W4964, W4921, W4922, W4923, W4924, W4932, W4935, W4936, W4938, W4941, W4944, W46036, W5003, W4996, W4997, W4999, W5000, W45964, W5004, W5008, W45953, W5013, W4974, W46005, W4967, W45999, W4971, W4973, W4984, W4986, W4991, W4992, W4860, W4861, W46137, W4862, W4867, W4868, W4857, W46122, W46121, W46119, W4878, W4844, W4836, W4839, W4879, W4847, W4848, W4849, W4850, W4853, W4854, W4856, W4914, W4905, W4906, W4907, W4913, W4917, W4893, W4881, W4882, W4887, W4890, W4894, W4896, W4898, W4899, W46091, W5162, W5147, W45811, W5154, W12659, W5158, W5143, W5163, W5169, W5174, W5129, W45845, W5120, W45841, W5175, W5135, W5138, W5139, W5141, W5195, W45758, W5198, W5202, W45751, W5194, W5204, W5206, W5207, W5210, W5178, W5179, W45776, W5185, W45771, W5186, W5189, W45766, W5191, W5049, W5035, W45918, W5036, W5044, W5045, W5046, W45922, W5053, W5055, W5056, W5058, W5064, W5065, W5017, W5020, W5023, W5025, W5029, W5032, W5033, W45925, W45924, W45923, W5103, W45867, W5093, W5094, W5098, W5104, W5107, W5109, W5110, W5117, W5118, W5119, W45895, W5070, W5075, W45884, W45883, W5078, W5079, W5080, W5082, W5083, W5088, W4597, W4586, W4587, W4589, W4591, W4594, W4595, W4600, W4611, W4613, W4614, W4615, W4570, W4559, W4560, W4561, W4566, W46459, W4568, W4617, W4571, W4572, W4573, W4578, W4581, W46443, W4655, W4647, W4648, W4650, W4651, W4653, W4654, W4643, W4657, W46377, W4658, W4660, W4662, W4664, W4619, W4623, W46411, W4625, W4629, W4631, W4557, W46402, W4636, W4638, W4639, W4641, W4486, W4457, W4463, W4474, W46546, W4476, W4477, W4480, W4488, W4490, W4445, W4427, W4429, W4430, W4431, W4434, W4438, W4440, W4446, W4447, W46560, W4455, W4531, W4534, W4536, W46489, W4540, W46480, W4546, W4549, W4550, W4553, W46509, W4498, W4499, W46518, W4507, W4508, W46512, W4510, W4518, W4519, W4521, W4523, W4524, W4526, W4528, W4790, W4782, W4783, W4785, W46233, W4787, W4789, W4780, W4796, W4800, W4801, W46215, W4755, W4758, W4760, W4761, W4764, W4769, W4772, W4774, W4775, W4776, W46176, W4822, W4823, W4826, W4829, W4830, W4831, W46168, W4803, W4805, W4808, W4812, W46203, W4753, W4815, W46197, W4817, W46193, W4821, W4694, W4701, W4702, W4704, W4708, W4709, W4710, W4711, W4714, W4715, W46355, W4666, W4677, W4679, W4681, W46357, W46353, W4684, W4689, W4690, W4692, W4693, W4745, W4734, W4735, W4737, W4739, W46282, W4743, W4733, W4748, W46277, W4749, W4751, W46317, W46313, W4726, W43917, W4727, W4729, W4730, W20337, W20338, W20339, W20345, W20334, W30428, W20362, W30424, W20366, W20367, W20370, W20318, W20310, W30472, W20312, W30468, W20315, W30465, W30461, W20323, W20327, W30454, W20402, W20405, W20406, W30381, W30380, W20413, W30391, W30375, W30374, W30372, W20419, W20420, W20385, W30414, W30413, W20378, W20380, W20384, W20309, W30405, W30403, W30402, W20387, W20391, W20393, W20399, W20252, W20235, W30561, W20236, W30557, W30554, W20244, W20248, W20251, W30548, W30547, W20254, W30543, W20256, W30538, W20259, W20224, W30588, W30587, W20211, W20215, W20219, W20221, W20223, W20264, W30574, W20225, W30572, W30570, W20228, W20230, W30567, W30566, W20296, W20282, W30503, W20288, W30501, W30499, W30497, W30496, W30508, W20297, W20302, W30476, W20272, W20265, W30530, W30529, W20267, W20270, W30524, W20273, W20274, W20276, W30514, W20280, W20603, W20588, W20596, W30196, W30193, W20599, W20602, W30183, W20608, W20611, W20616, W30232, W30227, W20566, W20617, W20572, W20576, W20580, W20582, W20584, W30132, W30144, W30142, W20637, W20638, W30139, W20642, W20650, W20635, W20651, W30128, W20659, W30121, W30120, W30119, W30170, W20620, W30167, W30165, W30164, W20624, W30161, W20554, W20627, W30151, W20632, W30312, W20466, W30328, W20469, W30320, W20484, W20485, W20463, W30310, W30309, W20488, W30304, W20492, W20494, W20445, W20425, W20426, W20427, W30357, W20438, W20439, W20443, W30351, W20495, W30346, W30345, W20453, W30343, W20455, W20456, W20460, W30261, W20533, W20534, W20537, W20538, W30252, W20527, W30248, W20542, W20543, W30243, W20546, W20547, W20550, W30291, W30289, W20505, W20508, W20510, W20209, W20511, W30273, W30272, W20515, W20524, W20526, W30266, W30900, W30913, W30912, W30911, W30910, W30908, W30905, W19921, W19911, W19927, W30893, W19935, W30888, W19937, W30932, W19885, W19888, W19891, W19892, W19894, W30935, W30933, W19899, W19904, W30925, W19905, W19906, W19907, W19910, W19973, W19976, W19977, W30844, W30842, W30850, W19983, W19984, W19986, W30832, W19987, W19988, W19990, W30827, W19957, W19943, W30876, W30874, W30873, W19950, W19951, W19883, W30862, W30857, W30853, W30851, W31023, W31034, W19801, W31027, W19804, W31025, W31036, W31019, W31018, W31015, W19810, W19811, W19812, W19823, W31058, W19782, W31055, W31054, W31052, W19789, W19790, W19827, W19791, W19794, W31041, W31038, W19849, W19851, W19854, W19856, W19860, W19846, W19863, W19864, W19868, W19871, W30952, W19881, W30997, W19835, W19841, W30991, W19992, W30985, W30983, W19845, W20140, W20123, W30672, W20132, W20139, W20141, W20148, W20150, W30654, W30653, W20153, W30691, W30700, W30699, W20107, W20110, W20113, W20114, W30689, W30688, W30687, W30686, W20115, W30684, W20117, W30682, W20183, W30617, W20184, W20187, W20188, W20189, W20191, W30607, W30606, W30619, W20195, W30603, W20198, W20199, W30597, W20168, W20155, W20158, W20159, W30642, W20161, W20165, W30704, W20170, W30631, W20179, W30623, W20180, W20181, W20015, W20018, W30786, W20026, W20027, W20028, W20030, W20033, W30797, W20036, W20040, W30771, W20042, W20052, W20010, W19993, W30822, W20000, W20002, W30818, W20007, W30759, W30806, W20012, W30804, W30802, W20092, W30726, W30724, W30722, W20089, W20090, W20080, W20094, W30715, W30712, W20096, W20098, W30708, W20100, W20101, W20068, W30758, W30756, W30753, W30752, W20063, W20065, W20066, W20663, W30742, W20069, W20071, W20072, W30738, W30735, W30732, W21299, W29481, W21288, W29475, W21279, W21309, W29458, W21314, W21260, W21248, W29512, W21251, W21252, W21256, W29504, W29502, W21316, W21263, W21265, W29494, W29493, W29489, W21277, W29486, W21367, W21363, W21365, W29425, W29409, W29408, W21368, W29406, W21371, W29402, W21375, W21377, W29397, W21328, W21317, W21319, W21320, W21323, W21324, W21325, W21326, W21247, W29439, W21341, W21348, W21349, W21178, W29599, W29588, W29587, W29586, W29584, W29580, W21182, W21184, W29576, W29575, W29573, W21187, W21146, W29630, W21135, W29627, W21140, W29621, W29571, W21148, W21153, W21154, W29608, W21238, W21223, W21230, W29534, W21233, W29530, W21237, W21222, W29526, W21240, W29523, W29521, W21242, W21244, W21246, W21207, W21195, W21199, W29562, W21202, W29558, W29557, W21209, W21210, W29549, W29547, W21215, W21217, W21522, W21512, W21516, W21518, W21520, W29255, W29249, W21526, W29247, W21527, W21535, W29242, W21540, W21493, W21486, W29290, W21489, W21492, W29284, W29283, W21495, W29279, W29278, W21499, W21505, W21507, W21584, W29211, W21567, W21569, W29200, W21582, W21583, W29212, W29195, W29190, W21598, W21599, W21550, W29231, W21549, W29225, W29224, W21553, W21554, W21557, W21560, W29213, W21423, W29366, W21411, W29361, W21412, W21417, W21420, W29368, W21432, W21433, W29346, W21435, W21382, W21383, W21386, W29388, W21392, W21395, W21437, W29381, W29380, W29379, W21401, W21406, W21407, W21475, W29316, W29310, W21471, W21473, W29318, W21476, W21478, W29300, W21479, W21482, W21483, W21484, W21451, W21440, W21442, W21443, W29334, W21450, W21130, W21452, W21453, W21458, W21460, W21461, W20806, W29966, W20795, W20797, W20798, W20799, W20804, W29957, W20793, W20807, W20811, W29947, W20829, W20830, W29978, W29988, W29987, W29986, W20782, W20787, W29940, W20788, W20790, W29971, W20791, W20868, W20861, W20862, W20863, W20865, W29900, W29898, W29895, W20871, W20872, W20873, W20879, W29923, W29939, W20836, W20837, W20839, W20840, W29926, W29925, W29924, W20852, W29916, W20856, W20858, W30076, W20690, W30086, W30085, W30084, W30083, W20692, W30077, W20689, W20696, W20698, W20700, W30070, W20701, W30067, W20708, W30105, W30116, W20668, W30111, W20671, W20672, W30108, W20675, W30060, W20676, W30100, W30098, W30097, W30096, W20685, W30093, W30091, W30009, W20741, W20748, W20751, W20752, W20753, W30017, W30014, W20756, W30011, W30028, W30007, W20763, W30004, W20770, W29997, W29996, W29995, W20724, W30058, W20717, W30055, W20721, W20723, W20882, W30045, W30042, W30040, W30036, W30032, W30029, W29709, W29724, W21036, W21037, W21038, W29717, W29716, W21044, W21047, W21049, W21053, W29704, W29702, W21061, W21065, W29693, W21066, W29757, W21008, W29753, W21009, W29751, W21010, W29748, W21014, W29744, W21016, W29742, W21019, W21025, W29734, W21028, W29727, W21119, W29663, W21096, W21099, W21101, W29657, W21108, W21113, W29665, W21124, W21125, W21126, W21128, W29636, W29635, W29677, W21068, W21070, W21071, W21074, W29679, W21081, W21004, W21082, W21085, W21090, W29669, W21091, W21092, W21093, W20925, W20913, W20914, W20915, W29844, W29841, W20924, W29837, W29849, W29829, W20932, W20935, W29820, W20902, W29882, W29880, W20894, W20897, W20898, W20899, W20901, W29861, W20903, W20904, W29857, W20909, W29852, W20912, W29850, W20991, W29782, W29781, W20986, W20988, W20989, W20990, W29773, W20992, W20997, W20999, W21000, W21003, W20959, W29814, W20946, W29806, W29805, W19781, W20960, W20967, W20969, W20973, W20975, W29785, W18492, W18477, W32353, W18479, W18480, W32349, W18485, W18487, W18488, W18491, W32355, W18495, W18497, W18501, W32328, W18503, W32323, W18471, W18465, W18467, W18468, W32373, W32372, W32371, W32370, W32368, W18473, W32365, W18476, W32359, W18549, W32283, W32281, W32280, W32277, W32275, W18545, W18564, W18567, W32266, W18570, W32262, W18573, W18575, W18507, W32319, W18513, W18517, W18518, W18519, W18522, W18464, W32304, W18533, W32294, W18543, W18544, W18404, W18391, W32462, W18392, W32460, W18393, W32457, W18397, W18399, W32452, W32451, W18390, W18412, W32442, W18413, W32439, W18372, W18366, W32487, W32485, W18367, W18369, W18371, W32437, W18376, W18377, W32477, W32476, W18379, W32472, W18383, W32468, W32392, W32405, W32404, W32403, W18445, W18449, W18452, W32406, W18455, W18456, W32388, W32387, W18460, W18462, W18415, W18416, W18417, W18419, W18420, W18576, W18426, W18429, W18430, W32420, W18439, W32411, W32408, W32407, W18746, W32093, W18754, W32086, W18769, W32099, W18772, W18775, W18776, W32065, W18708, W18710, W18711, W18712, W32119, W32061, W18727, W18731, W18737, W18740, W32103, W32100, W18832, W32027, W32026, W18830, W32022, W18821, W32017, W18834, W18841, W32007, W32006, W18802, W32060, W32057, W32056, W18798, W18800, W32049, W32048, W32046, W32042, W18814, W18815, W18817, W18819, W32035, W18820, W18627, W18616, W32221, W32220, W18621, W32217, W18623, W18624, W32212, W18631, W32209, W32208, W18632, W18634, W32203, W18595, W32256, W18578, W18581, W32249, W32247, W18593, W18635, W18600, W32237, W18607, W18608, W18691, W32166, W18672, W32155, W32153, W18689, W32149, W18695, W18697, W18699, W32138, W32136, W32135, W18704, W18637, W18639, W18644, W32189, W18649, W32185, W32491, W18656, W18657, W18658, W32174, W32171, W32169, W18671, W18061, W18063, W32804, W18064, W18067, W32796, W32795, W32809, W18075, W18076, W18077, W18081, W18083, W18086, W32776, W32823, W18029, W18034, W18035, W18037, W32832, W32826, W18050, W18053, W32811, W32748, W18115, W32743, W32740, W32738, W32749, W32734, W18118, W18121, W18122, W18125, W18127, W32762, W18093, W18094, W32771, W18095, W18096, W18100, W32765, W32764, W18104, W18028, W18106, W32756, W32755, W18108, W32750, W32920, W32928, W17934, W17935, W32925, W17938, W17939, W32921, W17931, W32919, W32914, W32913, W32912, W17946, W32946, W32957, W17914, W32951, W17917, W17919, W17949, W32945, W17920, W17923, W17926, W32936, W32934, W17930, W17996, W32871, W32870, W18002, W18008, W17992, W18021, W32850, W18022, W18025, W32845, W32844, W32843, W17952, W32906, W17954, W32900, W17965, W32895, W17971, W17973, W17974, W17980, W32887, W17984, W17985, W17986, W32882, W32881, W32576, W32589, W32577, W18278, W18289, W18291, W32608, W18230, W18231, W32622, W18240, W18243, W18244, W18300, W32606, W18255, W32600, W18258, W18259, W18261, W32592, W32510, W18329, W18332, W32519, W32514, W18340, W18342, W18326, W18345, W18349, W32503, W32498, W18357, W18360, W32494, W32492, W18305, W32554, W32553, W32552, W18303, W18304, W32545, W18229, W18309, W18311, W18312, W32534, W32531, W32529, W18321, W18169, W18158, W18160, W32692, W32690, W18167, W18156, W18173, W18174, W18178, W18179, W18140, W18130, W18132, W18133, W18134, W18135, W18136, W32716, W32715, W32714, W32707, W18148, W18151, W18153, W18154, W18215, W18208, W18210, W32643, W18212, W18213, W18214, W32649, W18217, W18220, W18221, W32630, W18222, W18223, W18192, W18183, W32672, W32671, W18191, W32003, W18193, W18194, W18198, W18201, W18202, W32654, W32651, W18204, W31382, W19453, W31375, W19458, W31370, W19462, W31368, W31367, W19450, W31363, W19468, W31360, W31357, W19478, W19479, W19417, W31411, W31409, W19423, W31402, W19424, W19480, W31398, W19430, W19436, W19442, W31387, W31384, W19516, W19517, W31315, W19519, W31313, W19522, W31318, W19526, W19529, W19531, W31299, W19535, W31297, W31295, W19536, W19500, W19481, W19484, W31344, W19489, W31338, W19503, W19504, W19507, W19512, W19513, W19333, W31496, W31494, W19329, W31489, W19332, W31486, W19327, W19336, W31482, W31481, W19337, W19338, W19339, W31477, W19341, W19309, W19289, W31524, W19292, W31515, W19306, W31513, W19308, W19350, W31510, W19310, W19313, W19315, W31506, W19321, W19322, W31502, W19325, W19404, W31438, W19395, W31435, W19389, W19406, W19408, W31416, W19371, W19352, W19353, W19362, W19363, W19537, W19375, W31452, W19376, W19379, W19383, W31447, W31445, W19386, W19693, W19696, W31133, W31132, W19704, W31128, W19709, W31123, W31121, W31178, W31176, W19665, W31171, W19670, W31168, W31166, W31120, W19676, W31162, W19677, W31159, W19679, W31155, W31152, W31151, W31076, W19738, W19739, W31091, W19740, W31085, W31078, W19758, W31074, W19762, W19766, W19770, W19771, W19778, W31119, W31117, W31115, W19716, W31113, W19719, W19723, W31108, W31106, W31100, W19732, W19734, W31097, W31247, W19581, W31257, W31256, W19582, W19583, W31253, W19587, W31261, W19597, W19598, W19601, W19602, W19603, W31234, W31291, W19548, W19549, W31281, W31280, W19552, W19604, W31270, W19565, W31267, W19568, W19573, W19576, W19641, W31202, W19633, W19636, W19630, W19643, W19644, W19645, W19656, W19657, W19658, W31230, W19607, W31228, W31226, W19610, W31223, W31221, W19614, W19617, W19625, W19626, W31844, W18984, W31851, W31850, W31846, W18994, W19001, W31841, W19004, W19005, W19007, W19008, W18968, W31890, W31888, W31885, W31880, W18964, W18967, W31871, W18972, W18975, W18976, W19047, W31793, W19051, W19054, W31788, W19056, W19058, W19066, W31774, W19068, W19071, W31768, W31765, W19073, W19033, W19011, W31829, W31827, W31820, W31817, W31816, W19028, W31891, W19036, W19039, W19040, W19042, W19045, W18886, W18877, W31971, W31970, W31968, W31967, W18883, W18888, W18890, W31957, W31955, W31952, W18859, W18846, W18849, W18851, W31994, W31950, W18862, W18863, W18864, W18869, W31980, W18874, W31977, W18876, W31903, W31920, W18929, W18936, W31911, W18939, W31907, W18943, W18924, W18946, W18947, W18949, W31898, W18950, W18951, W31894, W18906, W31949, W18898, W18899, W18900, W31944, W31940, W31937, W18911, W31933, W31930, W18915, W18918, W31924, W31596, W31613, W19223, W31609, W19228, W31604, W19233, W31600, W19238, W19221, W31595, W19242, W31587, W31586, W31585, W31584, W19209, W31644, W19195, W31642, W31637, W19205, W19207, W31583, W19214, W19215, W31621, W31619, W31617, W31616, W31545, W31557, W31556, W19264, W19268, W19271, W19273, W31559, W31542, W31541, W31540, W31535, W31534, W19249, W19251, W19254, W19255, W31576, W31573, W31572, W31570, W31569, W19260, W31564, W31563, W19262, W31560, W31717, W19105, W19106, W19107, W19110, W19111, W31724, W19120, W31733, W19121, W19122, W19123, W19127, W19128, W31707, W19133, W31755, W19085, W31750, W19095, W31742, W31741, W31740, W19102, W19171, W19176, W31663, W19182, W19183, W31672, W19184, W19188, W19191, W19192, W31650, W19193, W31647, W19141, W31699, W19143, W31697, W31696, W19154, W19155, W21603, W19159, W31684, W19160, W19161, W19162, W31678, W19167, W31675, W24128, W26624, W26623, W24117, W24118, W24122, W24125, W26613, W26625, W24133, W26603, W24140, W26599, W26593, W24096, W24081, W24082, W24085, W26649, W26646, W24156, W26640, W24098, W26638, W26635, W26631, W26628, W26627, W26548, W26559, W24192, W24199, W24200, W26553, W26552, W26551, W26560, W26547, W24203, W24204, W24206, W26540, W26539, W26537, W26576, W26587, W26586, W24160, W24162, W24163, W24165, W24166, W26658, W26573, W26569, W24179, W26564, W24183, W23997, W23986, W23990, W23994, W26734, W23983, W24004, W26726, W24007, W24010, W24015, W26720, W24018, W24024, W26759, W23964, W26766, W23967, W23970, W26760, W26714, W23972, W23974, W26756, W26755, W23976, W23978, W26748, W24049, W24050, W26681, W26680, W24055, W24062, W24064, W26685, W24069, W26668, W24073, W26663, W24076, W26661, W24077, W24025, W26712, W26706, W24030, W26704, W26698, W24036, W24040, W24042, W24044, W26370, W26383, W24366, W26374, W24363, W24381, W24388, W26361, W26360, W26357, W26405, W26418, W24326, W26413, W24338, W26356, W26394, W24352, W24418, W24421, W26318, W26315, W24427, W24431, W26308, W26307, W26306, W24433, W24447, W24448, W26344, W24393, W26353, W24399, W24401, W26348, W26345, W26419, W26340, W26339, W26338, W26334, W24411, W24412, W26331, W24238, W26502, W24241, W24246, W26493, W26491, W26490, W24252, W26505, W26486, W26484, W24258, W26482, W26476, W24220, W26523, W24221, W26475, W26518, W26515, W24226, W26513, W26512, W24231, W24232, W26507, W24307, W26448, W26445, W26444, W26442, W26440, W26439, W24295, W26435, W26433, W24311, W24313, W24314, W24320, W24322, W26462, W26474, W24261, W26470, W24268, W24282, W23959, W24285, W26459, W26458, W24293, W27105, W27121, W27118, W23609, W23611, W23614, W27111, W23602, W23625, W27100, W23636, W27095, W23638, W27091, W23589, W23579, W23581, W23583, W23586, W23590, W23591, W27134, W27131, W23597, W27128, W27126, W23684, W23677, W27046, W23679, W27044, W27039, W23682, W23683, W27032, W23691, W27028, W23693, W27025, W27065, W27083, W27081, W27074, W23657, W27071, W23658, W27149, W27064, W27063, W23665, W23667, W27057, W23669, W27055, W23675, W23498, W23503, W27238, W27235, W23506, W27247, W27229, W27224, W23516, W27220, W27213, W23526, W23468, W23469, W27269, W27267, W23472, W23473, W27261, W27210, W23484, W23486, W27248, W23568, W27173, W23563, W27168, W23565, W27164, W27162, W23558, W27160, W23571, W27156, W23572, W23573, W23576, W23578, W23537, W27205, W27204, W23531, W27199, W27198, W23533, W27193, W27186, W23545, W27183, W23554, W23556, W23557, W23840, W26875, W23843, W26872, W26871, W23848, W26865, W23839, W26856, W26855, W23862, W23864, W26851, W23865, W26846, W26896, W23804, W23807, W26905, W23809, W23820, W26897, W26892, W26889, W23832, W26880, W23934, W23913, W23916, W23919, W23925, W23929, W23912, W26791, W26790, W26789, W23947, W26773, W23957, W26843, W26842, W23871, W23879, W23882, W23803, W26826, W23891, W23892, W23896, W23901, W23905, W23908, W23911, W26982, W23737, W26988, W26985, W23740, W23730, W26981, W23743, W26979, W23744, W26976, W23749, W23751, W23753, W23714, W27017, W23706, W27015, W23708, W27011, W27009, W27008, W23713, W23715, W27003, W27002, W26998, W23725, W23728, W23782, W23784, W26933, W23788, W23781, W26926, W26924, W26923, W23791, W26919, W23794, W23801, W23754, W26965, W26958, W26957, W23763, W23764, W23766, W23769, W23770, W26946, W23772, W23776, W25673, W25011, W25682, W25013, W25680, W25679, W25678, W25677, W25676, W25674, W25685, W25021, W25023, W25666, W25032, W24985, W24988, W25708, W24989, W24990, W24994, W25702, W25654, W24995, W25695, W25004, W25692, W25689, W25688, W25008, W25610, W25066, W25070, W25618, W25617, W25073, W25074, W25078, W25623, W25608, W25081, W25602, W25086, W25639, W25653, W25652, W25651, W25646, W25049, W25715, W25638, W25052, W25055, W25060, W25624, W24900, W25795, W25793, W25792, W24912, W24916, W25779, W24921, W25776, W24924, W25774, W24926, W24875, W25831, W25829, W24870, W24872, W25826, W24873, W25818, W24883, W25806, W25800, W25740, W25739, W24960, W24963, W25730, W24952, W25727, W25723, W24975, W25718, W25717, W24930, W24932, W24934, W24937, W25598, W24941, W25754, W24943, W25749, W24950, W25745, W25420, W25431, W25430, W25428, W25260, W25261, W25262, W25435, W25263, W25418, W25268, W25409, W25452, W25228, W25466, W25462, W25461, W25458, W25455, W25454, W25449, W25448, W25446, W25245, W25246, W25249, W25437, W25319, W25364, W25359, W25331, W25355, W25334, W25349, W25341, W25345, W25344, W25286, W25403, W25277, W25281, W25225, W25292, W25294, W25388, W25385, W25304, W25375, W25134, W25127, W25130, W25131, W25557, W25556, W25555, W25554, W25119, W25136, W25137, W25139, W25142, W25543, W25542, W25146, W25539, W25583, W25090, W25596, W25092, W25592, W25590, W25589, W25588, W25579, W25577, W25108, W25110, W25111, W25116, W25497, W25199, W25494, W25492, W25202, W25489, W25205, W25208, W25482, W25480, W25212, W25213, W25476, W25475, W25473, W25219, W25151, W25158, W25531, W25160, W25168, W25170, W25523, W24864, W25520, W25517, W25179, W25182, W24571, W24582, W24583, W26154, W24594, W26131, W24598, W26129, W26127, W26126, W26180, W26179, W26178, W24549, W26175, W24553, W24558, W24559, W24560, W26166, W26164, W24570, W24648, W26095, W26094, W24634, W24636, W24641, W24642, W24643, W24644, W26084, W24650, W24654, W24655, W26074, W24660, W24662, W24664, W24668, W26112, W26122, W24605, W26118, W24609, W26116, W24626, W26105, W24629, W24632, W26097, W24487, W24478, W26260, W24480, W24482, W26256, W24484, W24485, W26253, W24473, W26251, W26247, W24492, W26243, W26281, W24452, W26292, W26290, W26288, W24458, W24461, W26239, W24466, W26278, W26277, W26276, W24469, W26272, W26270, W26269, W24530, W24523, W24524, W26206, W26204, W24526, W26200, W24529, W26198, W26211, W24531, W24532, W24534, W24540, W24546, W26183, W24496, W24497, W26232, W26228, W26227, W24509, W24510, W24670, W26221, W24513, W26219, W26216, W24515, W24517, W25930, W24782, W24784, W24786, W25923, W25921, W25919, W24781, W24799, W25906, W24801, W24802, W25902, W25898, W24770, W24759, W24760, W25954, W25951, W24764, W24765, W25894, W25944, W25943, W24771, W24773, W24774, W25936, W25932, W24850, W24842, W24846, W25859, W25855, W25854, W25851, W25849, W25847, W24857, W24861, W25842, W25841, W25838, W25837, W25891, W25888, W25886, W25885, W24821, W24830, W24833, W24834, W25870, W25869, W25868, W26039, W26038, W26037, W26034, W24694, W24695, W24696, W26026, W24702, W26024, W24703, W26022, W24704, W26019, W26017, W26056, W26066, W24671, W24672, W24673, W26062, W26059, W24710, W24678, W24680, W26050, W26048, W26047, W26045, W24751, W25981, W24739, W24740, W25978, W25976, W25975, W24742, W24744, W24735, W24752, W24755, W25964, W25961, W25960, W25959, W24724, W24711, W26013, W26012, W24712, W24717, W26004, W26003, W24726, W25995, W24728, W25992, W25989, W25988, W25985, W25984, W22243, W22225, W28530, W28526, W28525, W22233, W22235, W28521, W22250, W22253, W22256, W28506, W28504, W22212, W22198, W22203, W22204, W22206, W28555, W28554, W28553, W28551, W22260, W22213, W22214, W28544, W28543, W22218, W28541, W28539, W22220, W22292, W22293, W22294, W28466, W22297, W28463, W28462, W28461, W22302, W22307, W22311, W28447, W28445, W22276, W28501, W22261, W28497, W22265, W22269, W28494, W28488, W22197, W22279, W22282, W28481, W22284, W22287, W28475, W28634, W22126, W28647, W28644, W22132, W22134, W28637, W22135, W28650, W22154, W22155, W22156, W22157, W22158, W28615, W28683, W22093, W28671, W22103, W28666, W22107, W22160, W22108, W22109, W22113, W22114, W28655, W22116, W28653, W22123, W28573, W28583, W22186, W22187, W22188, W28578, W28577, W22190, W28574, W28585, W22192, W22193, W22194, W28568, W28567, W22195, W28563, W28613, W28612, W28611, W28608, W28607, W22163, W28604, W22315, W22172, W22174, W22175, W28596, W22180, W28278, W22439, W28285, W28284, W22442, W28280, W22445, W28289, W22449, W22452, W22454, W22457, W22468, W28261, W28319, W22417, W22424, W22478, W28300, W28299, W28298, W22433, W28296, W28291, W28220, W28234, W22505, W28228, W22515, W22516, W22519, W28235, W22525, W28217, W28215, W22532, W22538, W22539, W28206, W28248, W28257, W28256, W22482, W22483, W28252, W28250, W28247, W22487, W22488, W22493, W22496, W28236, W28400, W22355, W28398, W22356, W28395, W28393, W28391, W22364, W28386, W28382, W22372, W28377, W28420, W28441, W28438, W22321, W28429, W22329, W22332, W22374, W28419, W28416, W22341, W28413, W22342, W22346, W22347, W22352, W22396, W28342, W22397, W28339, W22399, W22400, W28330, W22407, W28324, W22383, W28374, W22376, W22377, W22381, W28365, W28363, W22088, W28361, W22384, W22386, W22387, W28355, W28354, W21775, W21776, W21778, W21780, W29012, W21788, W29005, W21791, W29001, W29000, W28997, W21795, W28995, W21764, W29045, W21758, W29043, W29042, W29040, W29039, W21800, W21765, W21766, W29027, W21770, W21771, W21773, W28961, W28960, W21833, W21835, W21838, W21840, W21845, W28945, W28944, W28938, W21853, W28989, W21801, W21802, W21805, W21810, W21811, W21754, W28974, W21827, W28965, W28964, W21652, W21645, W29147, W29146, W21646, W29144, W21648, W29151, W29138, W21656, W21657, W29134, W21658, W29131, W21664, W21666, W21627, W21606, W21608, W29175, W29173, W21614, W29171, W21620, W21668, W21628, W21630, W29162, W29158, W21635, W29156, W21640, W21737, W21717, W29082, W21720, W21721, W21724, W21716, W21741, W21745, W29056, W21747, W29053, W29052, W29050, W21698, W21674, W21682, W21688, W29110, W29107, W28935, W29098, W21710, W29090, W21715, W29087, W22019, W28776, W22014, W28769, W22018, W22006, W28752, W22029, W28749, W22035, W22039, W22041, W28795, W21968, W28811, W28807, W28806, W28803, W21983, W21987, W21988, W28743, W21993, W28792, W22002, W28784, W22003, W28781, W28712, W28711, W22063, W28709, W22074, W28700, W28699, W28697, W28695, W28694, W22078, W22079, W28685, W28730, W22043, W22044, W28738, W28734, W28814, W28727, W28725, W28723, W28721, W22053, W28718, W21880, W28905, W21884, W28896, W28909, W21893, W28889, W28888, W28884, W21903, W21904, W28879, W21905, W21862, W28934, W28933, W21854, W28930, W21855, W21856, W21907, W28921, W28920, W21866, W21871, W21873, W28828, W28841, W21940, W28837, W21945, W21948, W21950, W28846, W28827, W21954, W21955, W28818, W21967, W28815, W28862, W28874, W28873, W28872, W21910, W28869, W21911, W21915, W22544, W21918, W21919, W21924, W21927, W21928, W28849, W21930, W23160, W23145, W27585, W23157, W23158, W23159, W27577, W23163, W27573, W27572, W27570, W27567, W27566, W23167, W23112, W27629, W27628, W23104, W27626, W23106, W27624, W23108, W23109, W27618, W27563, W27613, W27610, W27609, W27599, W27595, W27594, W23223, W27531, W23206, W27526, W23214, W23216, W23222, W23229, W27514, W27512, W23232, W23233, W23170, W23173, W27557, W27556, W27555, W27630, W23178, W23179, W27546, W27543, W23188, W23192, W27535, W27703, W27715, W27714, W27712, W23028, W27704, W27719, W23039, W23040, W23041, W27692, W23052, W23054, W27732, W23000, W23001, W27741, W27738, W27737, W23009, W23012, W27684, W23016, W27729, W23018, W27727, W23020, W27723, W23075, W23076, W27657, W23077, W23080, W27649, W23082, W23074, W23086, W23090, W23095, W23097, W23099, W27632, W23103, W27682, W23059, W23061, W23062, W27505, W23064, W27669, W23066, W27667, W27663, W23070, W23072, W23388, W23390, W23394, W23396, W23397, W27349, W27363, W23403, W23406, W23408, W27339, W27337, W27336, W27334, W23349, W27390, W27388, W23362, W27380, W27333, W27376, W27375, W23370, W27371, W27369, W23375, W23385, W27286, W23446, W27295, W23451, W23452, W23453, W23454, W23460, W23461, W23464, W27278, W27277, W27275, W27321, W23413, W27331, W23414, W23416, W23417, W27324, W27323, W23345, W27319, W23426, W27313, W27311, W23440, W27479, W23265, W23266, W23269, W27465, W27462, W27460, W23272, W27455, W27492, W27504, W27501, W27499, W27497, W23246, W23248, W27494, W23250, W27489, W27488, W27487, W23251, W27484, W23255, W27410, W27424, W23315, W23318, W23319, W23327, W27411, W27425, W27408, W27405, W27398, W23341, W23342, W23343, W27441, W23277, W27450, W27448, W23283, W23284, W23287, W22995, W23290, W27439, W23302, W23304, W23307, W23310, W22681, W22682, W28060, W28059, W22683, W22684, W22678, W22697, W22701, W28043, W28042, W28040, W22707, W28035, W22664, W28087, W22656, W22657, W28079, W22719, W28074, W28070, W22674, W28066, W22750, W22754, W27993, W27991, W27990, W22758, W27988, W27986, W27984, W22762, W22765, W27978, W22768, W28029, W28027, W22725, W28019, W22731, W22733, W28013, W28008, W22741, W22742, W28004, W22746, W28161, W22575, W22576, W28171, W22577, W22578, W22579, W22584, W22586, W22566, W28157, W22594, W28154, W22598, W28149, W22601, W28147, W28189, W28202, W22547, W22548, W28198, W28196, W22550, W22553, W22554, W28186, W22559, W28182, W22560, W22564, W22565, W22634, W22624, W28113, W28112, W22625, W22628, W22630, W22632, W22635, W28098, W22639, W22640, W22642, W22610, W22603, W28139, W22607, W28133, W22612, W28129, W28126, W22616, W28122, W22622, W22920, W27830, W22906, W22907, W22913, W22914, W27819, W27818, W22919, W27832, W22923, W22924, W22926, W27809, W27804, W22933, W27802, W27847, W22877, W22882, W22883, W22889, W27852, W22934, W22895, W22899, W27842, W27841, W27837, W27834, W27833, W22979, W22963, W22966, W22967, W22968, W27763, W22973, W22974, W22976, W22962, W22984, W22988, W22989, W22990, W22992, W22994, W22955, W27797, W27796, W27793, W22948, W22949, W22953, W27785, W27778, W22959, W22960, W22961, W27773, W27772, W22798, W22799, W22800, W22810, W22812, W27931, W27930, W22813, W22795, W22816, W22819, W22821, W22823, W27916, W27914, W22829, W22772, W27969, W27964, W27963, W22779, W22830, W22788, W22789, W22790, W27952, W27948, W27946, W27945, W27875, W27884, W22852, W27882, W22854, W27879, W27878, W22855, W22851, W22860, W27870, W22866, W22868, W27865, W22873, W22839, W27910, W27907, W22835, W22836, W27901, W17911, W27896, W22843, W22845, W22848, W22849, W27887, W27886, W38143, W12677, W12679, W38151, W38148, W12680, W38137, W38136, W38133, W38130, W12663, W12643, W38183, W12648, W38179, W12654, W38174, W12660, W12665, W12669, W38162, W38156, W12743, W12730, W38092, W38090, W12732, W12735, W38085, W12736, W12742, W12729, W12744, W12750, W12752, W12753, W12755, W12702, W12688, W12690, W38124, W12698, W38116, W38115, W12700, W12642, W38111, W12709, W38108, W12713, W12720, W12544, W38281, W12548, W12562, W12563, W38287, W12570, W38259, W12571, W38256, W12572, W12573, W12521, W38311, W12524, W12527, W12534, W12537, W38294, W12539, W12540, W12542, W12633, W12620, W12622, W12623, W38207, W38206, W12625, W38203, W12630, W12634, W12636, W12637, W38195, W38191, W12641, W12592, W12581, W12583, W38236, W12758, W12593, W12602, W12607, W12608, W12613, W38215, W12617, W12932, W12913, W12914, W12915, W12921, W37898, W12927, W12928, W37890, W12935, W37888, W37883, W12939, W12940, W12897, W37930, W12900, W37928, W37925, W12945, W12905, W37919, W12906, W12907, W12908, W37910, W12995, W12983, W37850, W12984, W12992, W12999, W13003, W13005, W13012, W37877, W12949, W37873, W37872, W12964, W12966, W37935, W37863, W12969, W37861, W12970, W12973, W37857, W12976, W12816, W12798, W12809, W38018, W12812, W38014, W12794, W38011, W12822, W12824, W12825, W38060, W12764, W12768, W12773, W12775, W12778, W12780, W37998, W12783, W38036, W12788, W38031, W12792, W38029, W12881, W12864, W12868, W12871, W37960, W12874, W37954, W12880, W12857, W37950, W12885, W37945, W12886, W12889, W37993, W37991, W12837, W12839, W12842, W12843, W38315, W37982, W37979, W12850, W37976, W12852, W12853, W37971, W38632, W12229, W38629, W12233, W12236, W12241, W12228, W12245, W12249, W38605, W12205, W38656, W12206, W12251, W12207, W38646, W12223, W38638, W38637, W12305, W12290, W38562, W12297, W38557, W38555, W12302, W12303, W12306, W12307, W38542, W12313, W38539, W12256, W12257, W12268, W38592, W12269, W12271, W38587, W12203, W38582, W38581, W38576, W38572, W12283, W12106, W38756, W12094, W12095, W12098, W38750, W12099, W38746, W12111, W12112, W12119, W12121, W38728, W12076, W12070, W38781, W12074, W12075, W38774, W12129, W12085, W12086, W12087, W12089, W38762, W12090, W38694, W12170, W12173, W38689, W12175, W12180, W12181, W12163, W12191, W12194, W38672, W12195, W12197, W12199, W12142, W12130, W12131, W12132, W12133, W38721, W12134, W12135, W12136, W12149, W12150, W12151, W38711, W12152, W12155, W12156, W38704, W12162, W38406, W38403, W12439, W12443, W12444, W12433, W12449, W12450, W38386, W38436, W12407, W12411, W12414, W12416, W12420, W12453, W12423, W38421, W12426, W38417, W38415, W12430, W12432, W38411, W12499, W12483, W38350, W12484, W38348, W12485, W38345, W12491, W38343, W38354, W12501, W12507, W12513, W38370, W12458, W38378, W12460, W12461, W12463, W38371, W12466, W12468, W12471, W38362, W12474, W12479, W12347, W12351, W38505, W12353, W38502, W38512, W12357, W38495, W12358, W12359, W38490, W12326, W12315, W12316, W38535, W12320, W12322, W38529, W12323, W12324, W12327, W12330, W12331, W12342, W12379, W12381, W12385, W12386, W38466, W12392, W12393, W12395, W12397, W38442, W12368, W38488, W38487, W12361, W12362, W38482, W12363, W12365, W13013, W38475, W12369, W12374, W12377, W38469, W38468, W13686, W13675, W37156, W13677, W13679, W13680, W13688, W13696, W13697, W37136, W13700, W13701, W37128, W13641, W13642, W37188, W37187, W13651, W13654, W13657, W13660, W37170, W13666, W13673, W37161, W13734, W13738, W37096, W37090, W13744, W13745, W13748, W13749, W13752, W37081, W37080, W13754, W13755, W13709, W13710, W13716, W13719, W13720, W13721, W13724, W13640, W13728, W37110, W37109, W37107, W13729, W13542, W37281, W13548, W13566, W37267, W13574, W37262, W13576, W13578, W13580, W13530, W13518, W13521, W37312, W13523, W13526, W13528, W13535, W13536, W13539, W37219, W37217, W13619, W13623, W37212, W37210, W13630, W13631, W13617, W13633, W37199, W37196, W13637, W37251, W13587, W37248, W13589, W13594, W13599, W37076, W13604, W13606, W13610, W37226, W37222, W36941, W13881, W13883, W13887, W13888, W13890, W13892, W36929, W13897, W36921, W36952, W36965, W13871, W36962, W36956, W13876, W36953, W36950, W13878, W36945, W36944, W13944, W13930, W13939, W36878, W36877, W13927, W36873, W36870, W36869, W13948, W36867, W13949, W36861, W13905, W13907, W36914, W36910, W13911, W13913, W13869, W13914, W36903, W36900, W13916, W13797, W13781, W13783, W13785, W13788, W13790, W13780, W37036, W13798, W13802, W13804, W37029, W37028, W13760, W37070, W13763, W13764, W13765, W13766, W37027, W37063, W13768, W13773, W37055, W13775, W36999, W13837, W36996, W13839, W13841, W13836, W36983, W36982, W13852, W36978, W13854, W36975, W13858, W37015, W13805, W13807, W13808, W13809, W37021, W37020, W13810, W13815, W13817, W37012, W37011, W13822, W13825, W37005, W13833, W13834, W13162, W13163, W13164, W13169, W13172, W37653, W13175, W37648, W37645, W37643, W13183, W13139, W13140, W13142, W13145, W13186, W13151, W13153, W13158, W13159, W13160, W13254, W37601, W13231, W37599, W13239, W13247, W37590, W13253, W37603, W37583, W37582, W37577, W37575, W37570, W13271, W13212, W37638, W37637, W13191, W37620, W13214, W13218, W13221, W37609, W13226, W37607, W37783, W37781, W13060, W13063, W13066, W13073, W13056, W37763, W37761, W37758, W13078, W37755, W37812, W13016, W13018, W13020, W37815, W13023, W13034, W13036, W13037, W13045, W13051, W13119, W13113, W37722, W37721, W13115, W13121, W13122, W37704, W13126, W37700, W13130, W13084, W13087, W13089, W13093, W13094, W13275, W37739, W13097, W37735, W13103, W13106, W13109, W13110, W37411, W37409, W37408, W37403, W13441, W37395, W37393, W13431, W13454, W13455, W13458, W13460, W37380, W13464, W13395, W13399, W13403, W37439, W13405, W37434, W37376, W37431, W37430, W13421, W13422, W37421, W13428, W37413, W37333, W13492, W13497, W13498, W13503, W37332, W37331, W37330, W37329, W13506, W13509, W13513, W37359, W13466, W37374, W13471, W13477, W13479, W37447, W37355, W13482, W13483, W13485, W37350, W37519, W37533, W13313, W13317, W13324, W37522, W37516, W13328, W13337, W37507, W13338, W13276, W13279, W13284, W13295, W13296, W13297, W37504, W13298, W37546, W13301, W13302, W13309, W37538, W13382, W37476, W37475, W13362, W13367, W13371, W13375, W13379, W37460, W13383, W13384, W13387, W13390, W13392, W13339, W13340, W37500, W13345, W13346, W37493, W13349, W13350, W37489, W37488, W37487, W13355, W10829, W10821, W10823, W10825, W10826, W10827, W10828, W10830, W10837, W40031, W10844, W10845, W10846, W40082, W10789, W10793, W10798, W10799, W10800, W40068, W40065, W10805, W40024, W10807, W10809, W10810, W10812, W10813, W40054, W10815, W10874, W10881, W39987, W10883, W39983, W10888, W10891, W10893, W10912, W40023, W10848, W10852, W10854, W10855, W10858, W10860, W40001, W10866, W10867, W10869, W40178, W40176, W40175, W10693, W10698, W40169, W10703, W10706, W10712, W10714, W10715, W40202, W10655, W10662, W10669, W40147, W10671, W10677, W40185, W40184, W10766, W10750, W40114, W40111, W10756, W10770, W10774, W10775, W10776, W40086, W10780, W10732, W10727, W10728, W40137, W39955, W10734, W10737, W10741, W40128, W11071, W39810, W11060, W11065, W11066, W39799, W11067, W11075, W11078, W11084, W39788, W39786, W11030, W11016, W11020, W11025, W39831, W11027, W11037, W39819, W11042, W11046, W11047, W11049, W11117, W39752, W39748, W11120, W11116, W39745, W11121, W11122, W11124, W11126, W11127, W11110, W11092, W11093, W11094, W11095, W11098, W11104, W11107, W11108, W39767, W39766, W39765, W11113, W11115, W39757, W10936, W39918, W10941, W10943, W10927, W39914, W39909, W10948, W39906, W10949, W10953, W10954, W10918, W10913, W10914, W39948, W39946, W10959, W39942, W10921, W10925, W39934, W39933, W10926, W11007, W11001, W11003, W39858, W11000, W39854, W39848, W11013, W39897, W10961, W10969, W10970, W39890, W10974, W10977, W10646, W10980, W10983, W39879, W10990, W10994, W39870, W10351, W10329, W40552, W40550, W10341, W10342, W10345, W10350, W10327, W40538, W40536, W10356, W10363, W40529, W10371, W40524, W10376, W40566, W10306, W10307, W10310, W10311, W40570, W10313, W10314, W40521, W10320, W10322, W40559, W10325, W10326, W40556, W10414, W10398, W40488, W10405, W10406, W10408, W10411, W40474, W10418, W10420, W10421, W10425, W40466, W10426, W40510, W40502, W10303, W10391, W10392, W10393, W10394, W10395, W10397, W10228, W10218, W10219, W10220, W10227, W40649, W10229, W40647, W10231, W40643, W10233, W10234, W10201, W10188, W10193, W10195, W10196, W10198, W40679, W10236, W40674, W10205, W10206, W40670, W10210, W40664, W10278, W10280, W40594, W10289, W10273, W10291, W10296, W10297, W10300, W10302, W10255, W10238, W10239, W10240, W10248, W40626, W40625, W10427, W10261, W10262, W10264, W10267, W10268, W10572, W10566, W40311, W40310, W10568, W40307, W40305, W10569, W40314, W40299, W10575, W10579, W10581, W10532, W10534, W40340, W10539, W10541, W10542, W10546, W40333, W10548, W10557, W40320, W10558, W10559, W10622, W40243, W40241, W40240, W10635, W10637, W10640, W40226, W10645, W10595, W10582, W40286, W40284, W10587, W10589, W10594, W10530, W40271, W10597, W40267, W10604, W40262, W40260, W10607, W10463, W10448, W40431, W10455, W40423, W10464, W10471, W10472, W10473, W10428, W10430, W10431, W10433, W40450, W10436, W10438, W10439, W40440, W10521, W40374, W10517, W40364, W10518, W10519, W10510, W10522, W10523, W10527, W10528, W40354, W40349, W10493, W40404, W10484, W10492, W40392, W10495, W10496, W10501, W10509, W11750, W11737, W11739, W11740, W11746, W11748, W11755, W11756, W11760, W39094, W39092, W11762, W11763, W11718, W11703, W11708, W39144, W11715, W11717, W11765, W11721, W11723, W11725, W11726, W11727, W11731, W11735, W11841, W11811, W39049, W11821, W11824, W39040, W39038, W11834, W39052, W11843, W39028, W11845, W39023, W11852, W11853, W11791, W11774, W39079, W11778, W11779, W11785, W11787, W11702, W11792, W11793, W39061, W11802, W11803, W11806, W11614, W11603, W11606, W11612, W11613, W39251, W39229, W11617, W11622, W11625, W11627, W11588, W39276, W39275, W11573, W11575, W11583, W11585, W11587, W11589, W11591, W11593, W39258, W11595, W11596, W11671, W11676, W11677, W11679, W11682, W11687, W39183, W11689, W11695, W11698, W11700, W11634, W39206, W11636, W11637, W11643, W11648, W11855, W11652, W11657, W11658, W11665, W11668, W12007, W11993, W38868, W12000, W38862, W12004, W12005, W11992, W12008, W12014, W12016, W12021, W38843, W11981, W11972, W11973, W11975, W11978, W11979, W12027, W11982, W38882, W11987, W11989, W11990, W38873, W12046, W38806, W12049, W12052, W12054, W38798, W38796, W12055, W12056, W12061, W12063, W38789, W12064, W12068, W12034, W38831, W12033, W38825, W11971, W12035, W38822, W12039, W38814, W11910, W11897, W38986, W11900, W11903, W38973, W11893, W38970, W38963, W11917, W38959, W38958, W11872, W11856, W11858, W11860, W39010, W11866, W11869, W38957, W11875, W11877, W11881, W38996, W38993, W11890, W11955, W38926, W11946, W38922, W11948, W38920, W38913, W11959, W11960, W11962, W11963, W11967, W11968, W11925, W11926, W11928, W11929, W38944, W11934, W11938, W11940, W38932, W11288, W11262, W11264, W11268, W11271, W11273, W11279, W11283, W11261, W11289, W11290, W11291, W39581, W11248, W11238, W39629, W11239, W11240, W11242, W11294, W39619, W11249, W11250, W39616, W11254, W11260, W11335, W11320, W11321, W39545, W11323, W39536, W11332, W11338, W11339, W39525, W11343, W11295, W11296, W11300, W11301, W11302, W11303, W11304, W39635, W11309, W11310, W11312, W11314, W11315, W39552, W11318, W11173, W11151, W39705, W11158, W11159, W11164, W11165, W11167, W39695, W11176, W11184, W11185, W11187, W11192, W11193, W11195, W39734, W11135, W11136, W39726, W11137, W39724, W11198, W39719, W11140, W11145, W11146, W11217, W39655, W11218, W11219, W11224, W39648, W11225, W11228, W11234, W39637, W11210, W11204, W11205, W11206, W11207, W11208, W11209, W11347, W39666, W11211, W11212, W11214, W11215, W11501, W11485, W11489, W39359, W11494, W11499, W39353, W11481, W39349, W11504, W11506, W11507, W11509, W11457, W11452, W39398, W39397, W39396, W11454, W11455, W39382, W11472, W11473, W11479, W11547, W11529, W11537, W11539, W11540, W39312, W11556, W39285, W11561, W11565, W11566, W39280, W11518, W11510, W39336, W39335, W11512, W11516, W11523, W11525, W11526, W39315, W11390, W11371, W11373, W11374, W11383, W39476, W11389, W11370, W11394, W39469, W11397, W11398, W39460, W39503, W11349, W39511, W11353, W11358, W39508, W11361, W11399, W11365, W11366, W11369, W11437, W39427, W39426, W39421, W11432, W11435, W39417, W11428, W11440, W11441, W11442, W11443, W11400, W11403, W11404, W11407, W39439, W11419, W11420, W11426, W39431, W16635, W16639, W34251, W16641, W16643, W16644, W16633, W16647, W16650, W16653, W16606, W16612, W16613, W16662, W34269, W16620, W34267, W16626, W16629, W34259, W34189, W34202, W16694, W34197, W34196, W16697, W16706, W34178, W16717, W16718, W16677, W16663, W16664, W16667, W34227, W16672, W16673, W16675, W34220, W34286, W16683, W34213, W16685, W16686, W16513, W34383, W16501, W34377, W16505, W16506, W34373, W34370, W16515, W34361, W34360, W16522, W16527, W16529, W34353, W16477, W16447, W34416, W16459, W16467, W16471, W16478, W16481, W16486, W16492, W16493, W16591, W16576, W16577, W16578, W34310, W16585, W34305, W34304, W16575, W34298, W16598, W16601, W16605, W16558, W16538, W16540, W16546, W16550, W34331, W16566, W34325, W16567, W16572, W16898, W34018, W16881, W16886, W34012, W16892, W34005, W34003, W16905, W16907, W16910, W33991, W33989, W16845, W34049, W16852, W16864, W16866, W16912, W16869, W16870, W16872, W16873, W16952, W16954, W33949, W16957, W16959, W16960, W16962, W16964, W16948, W33937, W16970, W16974, W33931, W33929, W33927, W33970, W16913, W16917, W16922, W33972, W33971, W34057, W33968, W16939, W16942, W16943, W16741, W34145, W34140, W16753, W34132, W16771, W34121, W16774, W16777, W34115, W34158, W16723, W16725, W16726, W16727, W16731, W34157, W16736, W34153, W16738, W34150, W34149, W16825, W16812, W16815, W16817, W16818, W34078, W16820, W34073, W16823, W16829, W16834, W34059, W16781, W16785, W34105, W34104, W16794, W16796, W16798, W16804, W34093, W34091, W34089, W16808, W16082, W16072, W34747, W34746, W34745, W16074, W16081, W16071, W34736, W16087, W16091, W34730, W34728, W16093, W34725, W16062, W34775, W16047, W16051, W16054, W34766, W34765, W16058, W16060, W34723, W16063, W16064, W16065, W16068, W34753, W16132, W34697, W16123, W16126, W16127, W16128, W34690, W16129, W34686, W34685, W16135, W16148, W34722, W34719, W16101, W16103, W34712, W34710, W34708, W16110, W16114, W16115, W16118, W16121, W16122, W15980, W34858, W15968, W15975, W15978, W15979, W15964, W15981, W15983, W15986, W15987, W15988, W34835, W15991, W34886, W15947, W15948, W15949, W34880, W34877, W15953, W15955, W34831, W34872, W34871, W15957, W15959, W34866, W15960, W34861, W34806, W34803, W34799, W16029, W34797, W34796, W16015, W16031, W34792, W34791, W34783, W16040, W16041, W34829, W15996, W15998, W16000, W34821, W16001, W16003, W16149, W16006, W34815, W16007, W16010, W16011, W16014, W34808, W16340, W16349, W34504, W34502, W16334, W34496, W16360, W16361, W16369, W34486, W16373, W34528, W16313, W16315, W16319, W16322, W16325, W34529, W16326, W16327, W16330, W34522, W16332, W16333, W34519, W16409, W34453, W16412, W16414, W16421, W34444, W16423, W16407, W16430, W16431, W34435, W34431, W34428, W16376, W34480, W16377, W16378, W34475, W16382, W16386, W16307, W16391, W16393, W16397, W16398, W16400, W16402, W16406, W16228, W16200, W16202, W16206, W16208, W16213, W34615, W34636, W16229, W16230, W34610, W16234, W34604, W34603, W16186, W16165, W34659, W16176, W16184, W16236, W16190, W16191, W16192, W16193, W34643, W16194, W34641, W34639, W34638, W16290, W16276, W16280, W16281, W16282, W16286, W16287, W16289, W16293, W16294, W34548, W16300, W16306, W16244, W34597, W16250, W16251, W16256, W16263, W16264, W16265, W34579, W16266, W16269, W16270, W17627, W33284, W17603, W33279, W17608, W17616, W17618, W17623, W33266, W17630, W17633, W17635, W33257, W17639, W17588, W33319, W33315, W17567, W17574, W17576, W33304, W17586, W33253, W33298, W17591, W17592, W17594, W17597, W17666, W17655, W33227, W33225, W17660, W17664, W17652, W33215, W17669, W33206, W17673, W33203, W17644, W33246, W33244, W17646, W17650, W33234, W33391, W17495, W33402, W33400, W33396, W33395, W17502, W17493, W17503, W33386, W33385, W33383, W17509, W17510, W33423, W33434, W33433, W33430, W17477, W17511, W17480, W33418, W33415, W17488, W33408, W17551, W17538, W17541, W33344, W17550, W17537, W33335, W17556, W17559, W17562, W33362, W33376, W17515, W33372, W17517, W17518, W17521, W17523, W33366, W17526, W17527, W17529, W33357, W17532, W17533, W33352, W17833, W33053, W33052, W17826, W17830, W33045, W17821, W17834, W17836, W33035, W33033, W33032, W33031, W33080, W33079, W33075, W33074, W17803, W17804, W33024, W17810, W17813, W33063, W17817, W17818, W17819, W33057, W17897, W17878, W32984, W32983, W17892, W32975, W17895, W32989, W17901, W32966, W17905, W17908, W33021, W17852, W17854, W33014, W33013, W17856, W33010, W33009, W17787, W17859, W17862, W33001, W17871, W32995, W32990, W17702, W17704, W17705, W33158, W17711, W33167, W17713, W17714, W33151, W17718, W17721, W17722, W17723, W33144, W33185, W33198, W17678, W33193, W33191, W33190, W17689, W33177, W17698, W33173, W17699, W17700, W33170, W33168, W33099, W17761, W17764, W17768, W33103, W33100, W17773, W33095, W17776, W17786, W33127, W33142, W33141, W33139, W17733, W17737, W17741, W17742, W17467, W17743, W17744, W33124, W17745, W17748, W17753, W17133, W33771, W17137, W33762, W17143, W33759, W17123, W33757, W17145, W17147, W17148, W33752, W33751, W33750, W17149, W17099, W17102, W33803, W17104, W33799, W17109, W17113, W33791, W17115, W17120, W33782, W33779, W17211, W17181, W17186, W33716, W33710, W33703, W33696, W17215, W17217, W33687, W33746, W33745, W17157, W33739, W33737, W17162, W33729, W17167, W17175, W17178, W17036, W17018, W17021, W17028, W33884, W33878, W33876, W17038, W17041, W17042, W33870, W33868, W17045, W33865, W17004, W33920, W33912, W33910, W33863, W17005, W33907, W17007, W17011, W17013, W17014, W33896, W17085, W33827, W17086, W17078, W17090, W33817, W17091, W17094, W17061, W17048, W17050, W33860, W33858, W17053, W17058, W33686, W33845, W17067, W17074, W33840, W17075, W33531, W33529, W33528, W17368, W17376, W33517, W33516, W33514, W33511, W17383, W17386, W33506, W17387, W33564, W17331, W33559, W17337, W17338, W33555, W17341, W17342, W17345, W17346, W17347, W33542, W17355, W17360, W33449, W17437, W17438, W17456, W17421, W17457, W33446, W17462, W17463, W33440, W17465, W17466, W33489, W33503, W33501, W17394, W17396, W17397, W17401, W33494, W33491, W33565, W17406, W17407, W17408, W33482, W17415, W17420, W33641, W17252, W33652, W17255, W17257, W33642, W33656, W17264, W17267, W33634, W17223, W17224, W17225, W33678, W17232, W17272, W17238, W33668, W17239, W17244, W17246, W33657, W33590, W33588, W17311, W33586, W17314, W17317, W17308, W17323, W17325, W17328, W33571, W33568, W17288, W17275, W17276, W17278, W17280, W33617, W17285, W17287, W15945, W33605, W33603, W33598, W33592, W14617, W36216, W14602, W14604, W14606, W14607, W36208, W36205, W14595, W14619, W14622, W14623, W14624, W14626, W14627, W36191, W14585, W36243, W14570, W14577, W36237, W14582, W14583, W14584, W14586, W14588, W14589, W14593, W36140, W36154, W14668, W14669, W36148, W14675, W36144, W36142, W36135, W14684, W36132, W14685, W36130, W14641, W14630, W36181, W14637, W36177, W36175, W36245, W14644, W14647, W14648, W14651, W14656, W14657, W36160, W14661, W14468, W36339, W36337, W36336, W14475, W14481, W36326, W14486, W14467, W36319, W36318, W36317, W14491, W14492, W14495, W36358, W14443, W14446, W14449, W36362, W14451, W14497, W36353, W36350, W36348, W14463, W14464, W14465, W14534, W14535, W36277, W36270, W14532, W14547, W14561, W14565, W14519, W14504, W14505, W14507, W14515, W36298, W36295, W14688, W14521, W14526, W14527, W14529, W14531, W35987, W35986, W35984, W35982, W14820, W35978, W14827, W35988, W14834, W14838, W35962, W35961, W14808, W36011, W14799, W14800, W14801, W14802, W14807, W14809, W14811, W35994, W14817, W14882, W14870, W14875, W14878, W14879, W14886, W14888, W35907, W35899, W35939, W14851, W14854, W35947, W35944, W35941, W14859, W14861, W14862, W14863, W14864, W14865, W14867, W36099, W14714, W14716, W14719, W36093, W36091, W14724, W14726, W14728, W14729, W36080, W14730, W14696, W14689, W14691, W36125, W36123, W14692, W14694, W36118, W14731, W14698, W14701, W14702, W14703, W14705, W36107, W14710, W14712, W14761, W14764, W36041, W14769, W14775, W14778, W14780, W14758, W14788, W14789, W14794, W36015, W36077, W36076, W14735, W14737, W14738, W14740, W14743, W36060, W14748, W14751, W14129, W14116, W14118, W36709, W36708, W14119, W14120, W36703, W14115, W36696, W14130, W14132, W14139, W14140, W14142, W36687, W36729, W14085, W14086, W36734, W14092, W36731, W14093, W36678, W14098, W36725, W14103, W36720, W14107, W36718, W14109, W14182, W14173, W36649, W14174, W14176, W36644, W14178, W14179, W14183, W14190, W14194, W14198, W14160, W36674, W36672, W14156, W14158, W14159, W36667, W14163, W36663, W14164, W14166, W14169, W14171, W36821, W13992, W36827, W13998, W13990, W13999, W14001, W14003, W14005, W36813, W36811, W36843, W36859, W13955, W13959, W13962, W13963, W13969, W13971, W13975, W14007, W36842, W13978, W13980, W13985, W13987, W14059, W36768, W14062, W14063, W14064, W14066, W36757, W14057, W36755, W14070, W14078, W14079, W14080, W36747, W14082, W14029, W36809, W36805, W14016, W14021, W36798, W36795, W14024, W14208, W36789, W14039, W14041, W14042, W14052, W14053, W36448, W14364, W14365, W14370, W14373, W36457, W36452, W14359, W36445, W36444, W36443, W36440, W14348, W14338, W14339, W36493, W14340, W14344, W14349, W14357, W14410, W14412, W14415, W36402, W36400, W14406, W36388, W36386, W36378, W14442, W14387, W14388, W36432, W14391, W36427, W14394, W36424, W14397, W14398, W14400, W14401, W36415, W14405, W14250, W14238, W14240, W14241, W36584, W14245, W36578, W14248, W14237, W14252, W14255, W14260, W14262, W14266, W36557, W14223, W36618, W14209, W36616, W36615, W14211, W14218, W36610, W14267, W14228, W14229, W14233, W14236, W14301, W14303, W36517, W14310, W14312, W14315, W14327, W14331, W14332, W36503, W14333, W14337, W36541, W36555, W14274, W14277, W14278, W14280, W36540, W14285, W14296, W36532, W36529, W14298, W15568, W15570, W35233, W15576, W15577, W35229, W35227, W15583, W15587, W35220, W35219, W15592, W35216, W15594, W15548, W35284, W15525, W15531, W35277, W15540, W35269, W15543, W15546, W15595, W15550, W15555, W15557, W15558, W35252, W15562, W35248, W15654, W15647, W35167, W15649, W15651, W15655, W15662, W35152, W35150, W15667, W15668, W35190, W35210, W15604, W35207, W15616, W35195, W15631, W15636, W15637, W35181, W15640, W35176, W15645, W15429, W35375, W35374, W15414, W15417, W15422, W15424, W15425, W35376, W15433, W35356, W35355, W15439, W35353, W35352, W35387, W15399, W15400, W35395, W15445, W15411, W35384, W35382, W35377, W35306, W35313, W35311, W35310, W15490, W15491, W15493, W15483, W35303, W15500, W15502, W15505, W15509, W15520, W15521, W15470, W15449, W15450, W15451, W15453, W35341, W15454, W15670, W35329, W15473, W35326, W15481, W15482, W35321, W34977, W34976, W15851, W34972, W34971, W15852, W15859, W15844, W34959, W15878, W15880, W15881, W34946, W15893, W34997, W15814, W15817, W15819, W15822, W15823, W15896, W34995, W34993, W15832, W15833, W34986, W34897, W15926, W34905, W15931, W34900, W15933, W15935, W15937, W15939, W15940, W15941, W34891, W15942, W15944, W15908, W15899, W34935, W15904, W15905, W34930, W15906, W15911, W15913, W15915, W15921, W15925, W34911, W15724, W15712, W35107, W15715, W15716, W15720, W15722, W35111, W15725, W15729, W15733, W15735, W15736, W15741, W15747, W35126, W15671, W35142, W15672, W15678, W15679, W15683, W15688, W15690, W15694, W15696, W15697, W15700, W15705, W35040, W15783, W15784, W35037, W35036, W15789, W15792, W15781, W15796, W35027, W35023, W35022, W35021, W15803, W15812, W35072, W15752, W15754, W15759, W15761, W15768, W15392, W15769, W15771, W15777, W35045, W35043, W35726, W15058, W15059, W15063, W15064, W15066, W15067, W35727, W15073, W35722, W15074, W15075, W15077, W15081, W15084, W15035, W15025, W35762, W15026, W15031, W15032, W15038, W15047, W15055, W35677, W15132, W15135, W15136, W15140, W35666, W15147, W15148, W15150, W35660, W15151, W35658, W15156, W35711, W35705, W35704, W15096, W15099, W15100, W15108, W35765, W15111, W15112, W35693, W15116, W35688, W35687, W15119, W15131, W35851, W14930, W14931, W35855, W14934, W14935, W35852, W14924, W14943, W14944, W35838, W35837, W35835, W14951, W14952, W35877, W14900, W14901, W35884, W14905, W14914, W35876, W35874, W14918, W14919, W14922, W15009, W35793, W14997, W35787, W15000, W15008, W35798, W15011, W35778, W15012, W35776, W15013, W15022, W35767, W14957, W14961, W14963, W14964, W14965, W35817, W14976, W14977, W35808, W14978, W35805, W35804, W14983, W14987, W35493, W35491, W35489, W15305, W15307, W15314, W35478, W35477, W15321, W15323, W15287, W15275, W15276, W15282, W15284, W35512, W15285, W15288, W15291, W15296, W15301, W15304, W15380, W15358, W15359, W35435, W15372, W35423, W15377, W15378, W15357, W35419, W15382, W15390, W35409, W35452, W15331, W15333, W35460, W15341, W15343, W35454, W35523, W15347, W35448, W15348, W15349, W35442, W15352, W15356, W35602, W15192, W15197, W15198, W35604, W35617, W35600, W15205, W15208, W15212, W15217, W15183, W15161, W15173, W15177, W15181, W35625, W15187, W35623, W15190, W35620, W15191, W15257, W15251, W35549, W35548, W15249, W15258, W15260, W15262, W35535, W15265, W15267, W35525, W15222, W15225, W15229, W15234, W35571, W35570, W15235, W15236, W15237, W15240, W15245, W15246;

  NOR2X1 G0 (.A1(W778), .A2(W3643), .ZN(W12294));
  NOR2X1 G1 (.A1(W782), .A2(W20181), .ZN(W38549));
  NOR2X1 G2 (.A1(I854), .A2(I1248), .ZN(O591));
  NOR2X1 G3 (.A1(W30007), .A2(W34844), .ZN(O9647));
  NOR2X1 G4 (.A1(W2360), .A2(W9846), .ZN(W21249));
  NOR2X1 G5 (.A1(W2777), .A2(W2360), .ZN(W12301));
  NOR2X1 G6 (.A1(W4028), .A2(W7314), .ZN(W12299));
  NOR2X1 G7 (.A1(W7580), .A2(W9865), .ZN(W12296));
  NOR2X1 G8 (.A1(W2849), .A2(I966), .ZN(W12295));
  NOR2X1 G9 (.A1(W35515), .A2(W15976), .ZN(O9645));
  NOR2X1 G10 (.A1(W13521), .A2(W16906), .ZN(W21253));
  NOR2X1 G11 (.A1(W10526), .A2(W3469), .ZN(W12292));
  NOR2X1 G12 (.A1(W10291), .A2(W939), .ZN(O9653));
  NOR2X1 G13 (.A1(W23544), .A2(W8970), .ZN(W29509));
  NOR2X1 G14 (.A1(W7388), .A2(W883), .ZN(W12289));
  NOR2X1 G15 (.A1(W2309), .A2(W2397), .ZN(W12288));
  NOR2X1 G16 (.A1(W24083), .A2(W20601), .ZN(O9655));
  NOR2X1 G17 (.A1(W12830), .A2(W1193), .ZN(W29506));
  NOR2X1 G18 (.A1(W3308), .A2(W15183), .ZN(O2192));
  NOR2X1 G19 (.A1(W3044), .A2(W5405), .ZN(W12325));
  NOR2X1 G20 (.A1(I828), .A2(W24532), .ZN(O9633));
  NOR2X1 G21 (.A1(W20439), .A2(W32182), .ZN(W38530));
  NOR2X1 G22 (.A1(I1265), .A2(W6401), .ZN(W12321));
  NOR2X1 G23 (.A1(I814), .A2(W18654), .ZN(W21243));
  NOR2X1 G24 (.A1(W2221), .A2(W9046), .ZN(O593));
  NOR2X1 G25 (.A1(W3068), .A2(W8639), .ZN(W38533));
  NOR2X1 G26 (.A1(W2084), .A2(W27541), .ZN(W29517));
  NOR2X1 G27 (.A1(W18493), .A2(I1140), .ZN(W29503));
  NOR2X1 G28 (.A1(W18365), .A2(W22326), .ZN(W38537));
  NOR2X1 G29 (.A1(W11391), .A2(W5144), .ZN(W12314));
  NOR2X1 G30 (.A1(W22995), .A2(W36211), .ZN(W38540));
  NOR2X1 G31 (.A1(W28933), .A2(W16952), .ZN(O4930));
  NOR2X1 G32 (.A1(W5412), .A2(W9775), .ZN(W12310));
  NOR2X1 G33 (.A1(W6), .A2(W11328), .ZN(W12309));
  NOR2X1 G34 (.A1(W1118), .A2(W11936), .ZN(W12308));
  NOR2X1 G35 (.A1(W16175), .A2(W8954), .ZN(W21266));
  NOR2X1 G36 (.A1(W4654), .A2(W18637), .ZN(W21264));
  NOR2X1 G37 (.A1(W9162), .A2(W8306), .ZN(W12263));
  NOR2X1 G38 (.A1(I121), .A2(I1640), .ZN(W12262));
  NOR2X1 G39 (.A1(W4058), .A2(W663), .ZN(W12261));
  NOR2X1 G40 (.A1(W252), .A2(W9512), .ZN(W12260));
  NOR2X1 G41 (.A1(W2273), .A2(W17779), .ZN(O9672));
  NOR2X1 G42 (.A1(W5831), .A2(W28162), .ZN(W38599));
  NOR2X1 G43 (.A1(W15239), .A2(W560), .ZN(W38600));
  NOR2X1 G44 (.A1(W25362), .A2(W1067), .ZN(W38595));
  NOR2X1 G45 (.A1(W536), .A2(W16762), .ZN(O2196));
  NOR2X1 G46 (.A1(W9337), .A2(W10486), .ZN(W12253));
  NOR2X1 G47 (.A1(W12605), .A2(W34810), .ZN(O9674));
  NOR2X1 G48 (.A1(W8521), .A2(W6171), .ZN(W29496));
  NOR2X1 G49 (.A1(W15741), .A2(W211), .ZN(W21269));
  NOR2X1 G50 (.A1(W27499), .A2(W5520), .ZN(W29495));
  NOR2X1 G51 (.A1(W15284), .A2(W14614), .ZN(W38609));
  NOR2X1 G52 (.A1(W35134), .A2(W18522), .ZN(O9680));
  NOR2X1 G53 (.A1(W8863), .A2(W8965), .ZN(W12274));
  NOR2X1 G54 (.A1(W19474), .A2(W32420), .ZN(O9660));
  NOR2X1 G55 (.A1(W25859), .A2(W11030), .ZN(W29500));
  NOR2X1 G56 (.A1(W26847), .A2(W18466), .ZN(W38574));
  NOR2X1 G57 (.A1(W1731), .A2(W26664), .ZN(O9663));
  NOR2X1 G58 (.A1(W38562), .A2(W5045), .ZN(W38579));
  NOR2X1 G59 (.A1(W7505), .A2(W6965), .ZN(W12277));
  NOR2X1 G60 (.A1(W8169), .A2(W1723), .ZN(O588));
  NOR2X1 G61 (.A1(W11555), .A2(W20649), .ZN(W38580));
  NOR2X1 G62 (.A1(W1271), .A2(W78), .ZN(O9631));
  NOR2X1 G63 (.A1(W31724), .A2(I1505), .ZN(W38585));
  NOR2X1 G64 (.A1(W25755), .A2(W14255), .ZN(W29499));
  NOR2X1 G65 (.A1(W26586), .A2(W30094), .ZN(O9669));
  NOR2X1 G66 (.A1(W10858), .A2(W12091), .ZN(O2195));
  NOR2X1 G67 (.A1(W11216), .A2(W6311), .ZN(W38591));
  NOR2X1 G68 (.A1(W18537), .A2(W10673), .ZN(W21262));
  NOR2X1 G69 (.A1(W5841), .A2(W10528), .ZN(W12266));
  NOR2X1 G70 (.A1(W12793), .A2(W22598), .ZN(W38471));
  NOR2X1 G71 (.A1(W8076), .A2(I1001), .ZN(O9589));
  NOR2X1 G72 (.A1(W10318), .A2(W13417), .ZN(O2187));
  NOR2X1 G73 (.A1(W5685), .A2(W11942), .ZN(W29537));
  NOR2X1 G74 (.A1(W15365), .A2(W18474), .ZN(O2189));
  NOR2X1 G75 (.A1(W11907), .A2(I906), .ZN(W12378));
  NOR2X1 G76 (.A1(W3805), .A2(W19801), .ZN(W21229));
  NOR2X1 G77 (.A1(I186), .A2(I1256), .ZN(W12376));
  NOR2X1 G78 (.A1(W12235), .A2(W7083), .ZN(W12375));
  NOR2X1 G79 (.A1(W33186), .A2(W18719), .ZN(O9587));
  NOR2X1 G80 (.A1(W2574), .A2(W12252), .ZN(W12373));
  NOR2X1 G81 (.A1(W10994), .A2(W6616), .ZN(W12372));
  NOR2X1 G82 (.A1(I1873), .A2(W7893), .ZN(W12371));
  NOR2X1 G83 (.A1(W38288), .A2(W36433), .ZN(O9597));
  NOR2X1 G84 (.A1(W4619), .A2(W38206), .ZN(W38474));
  NOR2X1 G85 (.A1(W7348), .A2(W9121), .ZN(W38477));
  NOR2X1 G86 (.A1(W25070), .A2(W2944), .ZN(O4943));
  NOR2X1 G87 (.A1(W2307), .A2(W10418), .ZN(W12366));
  NOR2X1 G88 (.A1(W10436), .A2(W1338), .ZN(W12391));
  NOR2X1 G89 (.A1(W15724), .A2(W25538), .ZN(O9575));
  NOR2X1 G90 (.A1(W4191), .A2(W314), .ZN(W12398));
  NOR2X1 G91 (.A1(W12374), .A2(I1382), .ZN(O9578));
  NOR2X1 G92 (.A1(W10934), .A2(W29063), .ZN(W38444));
  NOR2X1 G93 (.A1(W10619), .A2(W9078), .ZN(W21220));
  NOR2X1 G94 (.A1(W2295), .A2(W5854), .ZN(W12394));
  NOR2X1 G95 (.A1(W2929), .A2(W22816), .ZN(O9580));
  NOR2X1 G96 (.A1(W12677), .A2(W14542), .ZN(W29543));
  NOR2X1 G97 (.A1(W8966), .A2(W24001), .ZN(O4942));
  NOR2X1 G98 (.A1(W7939), .A2(W8619), .ZN(W12390));
  NOR2X1 G99 (.A1(W9069), .A2(W22557), .ZN(O9583));
  NOR2X1 G100 (.A1(W20321), .A2(W26909), .ZN(W29541));
  NOR2X1 G101 (.A1(W20836), .A2(W2367), .ZN(W29540));
  NOR2X1 G102 (.A1(I405), .A2(W15011), .ZN(W29539));
  NOR2X1 G103 (.A1(W547), .A2(W8828), .ZN(O4944));
  NOR2X1 G104 (.A1(W3601), .A2(W1580), .ZN(W12384));
  NOR2X1 G105 (.A1(W1934), .A2(I303), .ZN(W12335));
  NOR2X1 G106 (.A1(W10781), .A2(W2547), .ZN(O595));
  NOR2X1 G107 (.A1(W10031), .A2(W3643), .ZN(W12343));
  NOR2X1 G108 (.A1(W1523), .A2(W3776), .ZN(W12341));
  NOR2X1 G109 (.A1(I446), .A2(W6824), .ZN(W12340));
  NOR2X1 G110 (.A1(W5065), .A2(W11620), .ZN(W12339));
  NOR2X1 G111 (.A1(W12214), .A2(W1161), .ZN(W12338));
  NOR2X1 G112 (.A1(W35551), .A2(W36111), .ZN(O9625));
  NOR2X1 G113 (.A1(W7994), .A2(W3115), .ZN(O594));
  NOR2X1 G114 (.A1(W10165), .A2(W1253), .ZN(W12345));
  NOR2X1 G115 (.A1(W4209), .A2(W5418), .ZN(W12334));
  NOR2X1 G116 (.A1(W16430), .A2(W23274), .ZN(W29525));
  NOR2X1 G117 (.A1(W6372), .A2(W8562), .ZN(W12332));
  NOR2X1 G118 (.A1(W15854), .A2(W24685), .ZN(O4935));
  NOR2X1 G119 (.A1(W23847), .A2(W21456), .ZN(O9629));
  NOR2X1 G120 (.A1(W9173), .A2(W3855), .ZN(W12329));
  NOR2X1 G121 (.A1(W13094), .A2(W27005), .ZN(W38524));
  NOR2X1 G122 (.A1(W21859), .A2(W12604), .ZN(O4932));
  NOR2X1 G123 (.A1(W11389), .A2(W4021), .ZN(W12354));
  NOR2X1 G124 (.A1(W763), .A2(W3479), .ZN(W12364));
  NOR2X1 G125 (.A1(W35486), .A2(W29881), .ZN(O9601));
  NOR2X1 G126 (.A1(W23883), .A2(W18827), .ZN(O9604));
  NOR2X1 G127 (.A1(W3330), .A2(W9883), .ZN(W21234));
  NOR2X1 G128 (.A1(W30709), .A2(W14691), .ZN(W38493));
  NOR2X1 G129 (.A1(W2088), .A2(W2213), .ZN(O9610));
  NOR2X1 G130 (.A1(W7598), .A2(I974), .ZN(W12356));
  NOR2X1 G131 (.A1(W20857), .A2(W15975), .ZN(O9615));
  NOR2X1 G132 (.A1(W10604), .A2(W28508), .ZN(W29490));
  NOR2X1 G133 (.A1(W34104), .A2(W32046), .ZN(W38504));
  NOR2X1 G134 (.A1(W9886), .A2(W3187), .ZN(O4938));
  NOR2X1 G135 (.A1(W21954), .A2(W3571), .ZN(W38508));
  NOR2X1 G136 (.A1(W11627), .A2(W2782), .ZN(W12350));
  NOR2X1 G137 (.A1(W9040), .A2(W16960), .ZN(W21236));
  NOR2X1 G138 (.A1(W1746), .A2(I1526), .ZN(W12348));
  NOR2X1 G139 (.A1(W11646), .A2(W32333), .ZN(W38511));
  NOR2X1 G140 (.A1(W6890), .A2(W1656), .ZN(O2210));
  NOR2X1 G141 (.A1(W7134), .A2(W2249), .ZN(W12148));
  NOR2X1 G142 (.A1(W9918), .A2(W11932), .ZN(W12147));
  NOR2X1 G143 (.A1(W11488), .A2(W2338), .ZN(W12146));
  NOR2X1 G144 (.A1(W24157), .A2(W10767), .ZN(O4907));
  NOR2X1 G145 (.A1(W710), .A2(W8012), .ZN(W12144));
  NOR2X1 G146 (.A1(W11780), .A2(W319), .ZN(W12143));
  NOR2X1 G147 (.A1(W11949), .A2(W8119), .ZN(W12141));
  NOR2X1 G148 (.A1(W5577), .A2(W2971), .ZN(W12140));
  NOR2X1 G149 (.A1(W33433), .A2(W6175), .ZN(W38714));
  NOR2X1 G150 (.A1(W1168), .A2(W706), .ZN(W12138));
  NOR2X1 G151 (.A1(W3905), .A2(W10626), .ZN(W12137));
  NOR2X1 G152 (.A1(W13896), .A2(W3345), .ZN(O2211));
  NOR2X1 G153 (.A1(W36080), .A2(W25809), .ZN(O9748));
  NOR2X1 G154 (.A1(W9811), .A2(W13291), .ZN(O4904));
  NOR2X1 G155 (.A1(W17576), .A2(W38469), .ZN(W38722));
  NOR2X1 G156 (.A1(W15235), .A2(W12774), .ZN(W21310));
  NOR2X1 G157 (.A1(W33203), .A2(W34828), .ZN(O9751));
  NOR2X1 G158 (.A1(W17611), .A2(W29211), .ZN(O4909));
  NOR2X1 G159 (.A1(W17106), .A2(W28318), .ZN(O9734));
  NOR2X1 G160 (.A1(W11076), .A2(W6475), .ZN(O9735));
  NOR2X1 G161 (.A1(W10139), .A2(W3118), .ZN(W12165));
  NOR2X1 G162 (.A1(W15967), .A2(W11817), .ZN(O2205));
  NOR2X1 G163 (.A1(W26017), .A2(W28993), .ZN(W29469));
  NOR2X1 G164 (.A1(W14781), .A2(W20191), .ZN(W21297));
  NOR2X1 G165 (.A1(I1591), .A2(W3007), .ZN(W21298));
  NOR2X1 G166 (.A1(W6335), .A2(W10227), .ZN(O572));
  NOR2X1 G167 (.A1(W23192), .A2(W3543), .ZN(O9752));
  NOR2X1 G168 (.A1(W12052), .A2(W7525), .ZN(W12157));
  NOR2X1 G169 (.A1(W15187), .A2(W26450), .ZN(W29466));
  NOR2X1 G170 (.A1(W24180), .A2(W6755), .ZN(O4908));
  NOR2X1 G171 (.A1(W20043), .A2(W4232), .ZN(W21303));
  NOR2X1 G172 (.A1(W17841), .A2(W11409), .ZN(O9742));
  NOR2X1 G173 (.A1(W1180), .A2(W15162), .ZN(O2207));
  NOR2X1 G174 (.A1(W578), .A2(W25899), .ZN(O9744));
  NOR2X1 G175 (.A1(W8353), .A2(W9482), .ZN(W12101));
  NOR2X1 G176 (.A1(W32870), .A2(W31473), .ZN(O9762));
  NOR2X1 G177 (.A1(W8218), .A2(W2076), .ZN(W12109));
  NOR2X1 G178 (.A1(W11575), .A2(W9833), .ZN(W12108));
  NOR2X1 G179 (.A1(W533), .A2(W22508), .ZN(O9763));
  NOR2X1 G180 (.A1(W18317), .A2(W19597), .ZN(O9764));
  NOR2X1 G181 (.A1(W10769), .A2(W379), .ZN(W12105));
  NOR2X1 G182 (.A1(W15650), .A2(W8956), .ZN(W38745));
  NOR2X1 G183 (.A1(W11270), .A2(W12872), .ZN(W29452));
  NOR2X1 G184 (.A1(W24733), .A2(W6874), .ZN(W38739));
  NOR2X1 G185 (.A1(W26875), .A2(W9389), .ZN(W29451));
  NOR2X1 G186 (.A1(W10012), .A2(W16718), .ZN(W29450));
  NOR2X1 G187 (.A1(W25036), .A2(W4848), .ZN(O4897));
  NOR2X1 G188 (.A1(W7561), .A2(W9546), .ZN(W12096));
  NOR2X1 G189 (.A1(W14566), .A2(W38346), .ZN(O9768));
  NOR2X1 G190 (.A1(W35623), .A2(W26461), .ZN(W38757));
  NOR2X1 G191 (.A1(W8960), .A2(W2289), .ZN(W12092));
  NOR2X1 G192 (.A1(W7687), .A2(W7881), .ZN(W29444));
  NOR2X1 G193 (.A1(W2480), .A2(I713), .ZN(O568));
  NOR2X1 G194 (.A1(W18083), .A2(W2300), .ZN(O4902));
  NOR2X1 G195 (.A1(W7859), .A2(W25769), .ZN(W38729));
  NOR2X1 G196 (.A1(W25590), .A2(W36628), .ZN(O9754));
  NOR2X1 G197 (.A1(W11167), .A2(W2403), .ZN(W12126));
  NOR2X1 G198 (.A1(W8612), .A2(W4695), .ZN(W12125));
  NOR2X1 G199 (.A1(W6372), .A2(W7986), .ZN(O569));
  NOR2X1 G200 (.A1(W10840), .A2(W5402), .ZN(W12123));
  NOR2X1 G201 (.A1(W10965), .A2(W12728), .ZN(W29455));
  NOR2X1 G202 (.A1(W1730), .A2(W8361), .ZN(W12168));
  NOR2X1 G203 (.A1(W31247), .A2(W31803), .ZN(O9757));
  NOR2X1 G204 (.A1(W19534), .A2(W24050), .ZN(O9760));
  NOR2X1 G205 (.A1(W3836), .A2(W6124), .ZN(W12116));
  NOR2X1 G206 (.A1(I1620), .A2(W9129), .ZN(W12115));
  NOR2X1 G207 (.A1(W2169), .A2(W9707), .ZN(W12114));
  NOR2X1 G208 (.A1(I361), .A2(I1176), .ZN(W12113));
  NOR2X1 G209 (.A1(W28991), .A2(W4301), .ZN(W38738));
  NOR2X1 G210 (.A1(W5356), .A2(W5313), .ZN(W12218));
  NOR2X1 G211 (.A1(W7399), .A2(I592), .ZN(W21278));
  NOR2X1 G212 (.A1(W24367), .A2(W29763), .ZN(O9695));
  NOR2X1 G213 (.A1(W6441), .A2(W6333), .ZN(W29485));
  NOR2X1 G214 (.A1(W7755), .A2(W17184), .ZN(O2201));
  NOR2X1 G215 (.A1(W36811), .A2(W11119), .ZN(W38644));
  NOR2X1 G216 (.A1(W9812), .A2(W21957), .ZN(W29484));
  NOR2X1 G217 (.A1(W5076), .A2(W4245), .ZN(W12220));
  NOR2X1 G218 (.A1(W26364), .A2(W34863), .ZN(O9702));
  NOR2X1 G219 (.A1(W37543), .A2(W4934), .ZN(W38634));
  NOR2X1 G220 (.A1(W5542), .A2(W10049), .ZN(W12217));
  NOR2X1 G221 (.A1(W1652), .A2(W38632), .ZN(O9703));
  NOR2X1 G222 (.A1(W4581), .A2(W8330), .ZN(W12215));
  NOR2X1 G223 (.A1(W5395), .A2(W7162), .ZN(W12214));
  NOR2X1 G224 (.A1(W5029), .A2(W5796), .ZN(W12213));
  NOR2X1 G225 (.A1(W22073), .A2(W19613), .ZN(W38650));
  NOR2X1 G226 (.A1(W630), .A2(W7987), .ZN(O9704));
  NOR2X1 G227 (.A1(W5389), .A2(W7947), .ZN(W12210));
  NOR2X1 G228 (.A1(W25212), .A2(W31907), .ZN(W38627));
  NOR2X1 G229 (.A1(W25623), .A2(W21715), .ZN(W38614));
  NOR2X1 G230 (.A1(W6378), .A2(W1789), .ZN(W12243));
  NOR2X1 G231 (.A1(W7854), .A2(W11428), .ZN(O2199));
  NOR2X1 G232 (.A1(W10496), .A2(W18463), .ZN(O2200));
  NOR2X1 G233 (.A1(W10675), .A2(I1143), .ZN(O583));
  NOR2X1 G234 (.A1(W3486), .A2(W7793), .ZN(W12238));
  NOR2X1 G235 (.A1(W29987), .A2(W9434), .ZN(W38623));
  NOR2X1 G236 (.A1(W15872), .A2(W4769), .ZN(W21276));
  NOR2X1 G237 (.A1(W3433), .A2(W10413), .ZN(O579));
  NOR2X1 G238 (.A1(W376), .A2(W12157), .ZN(W12234));
  NOR2X1 G239 (.A1(I1266), .A2(W27447), .ZN(O9691));
  NOR2X1 G240 (.A1(W6235), .A2(W3763), .ZN(W12232));
  NOR2X1 G241 (.A1(W4181), .A2(W826), .ZN(W12231));
  NOR2X1 G242 (.A1(W35939), .A2(W14413), .ZN(O9692));
  NOR2X1 G243 (.A1(W21018), .A2(W17819), .ZN(W29487));
  NOR2X1 G244 (.A1(W11470), .A2(W5900), .ZN(O9693));
  NOR2X1 G245 (.A1(W27793), .A2(W33263), .ZN(O9727));
  NOR2X1 G246 (.A1(W30454), .A2(W7473), .ZN(W38678));
  NOR2X1 G247 (.A1(W20294), .A2(W36678), .ZN(O9723));
  NOR2X1 G248 (.A1(I1260), .A2(W1941), .ZN(W12187));
  NOR2X1 G249 (.A1(W9428), .A2(W5417), .ZN(W12186));
  NOR2X1 G250 (.A1(W27892), .A2(W25304), .ZN(O4917));
  NOR2X1 G251 (.A1(W8049), .A2(W5320), .ZN(W12182));
  NOR2X1 G252 (.A1(W15853), .A2(W14626), .ZN(W21290));
  NOR2X1 G253 (.A1(W6038), .A2(W175), .ZN(O9726));
  NOR2X1 G254 (.A1(W2931), .A2(W2983), .ZN(W12190));
  NOR2X1 G255 (.A1(W110), .A2(W9832), .ZN(W12178));
  NOR2X1 G256 (.A1(W26283), .A2(W7793), .ZN(O4914));
  NOR2X1 G257 (.A1(W21203), .A2(W15818), .ZN(W38688));
  NOR2X1 G258 (.A1(W9476), .A2(W9591), .ZN(O9730));
  NOR2X1 G259 (.A1(W31774), .A2(W32085), .ZN(O9732));
  NOR2X1 G260 (.A1(W10135), .A2(W8284), .ZN(W12172));
  NOR2X1 G261 (.A1(W8255), .A2(W11792), .ZN(W12171));
  NOR2X1 G262 (.A1(W32390), .A2(W26141), .ZN(O9733));
  NOR2X1 G263 (.A1(W17874), .A2(W34971), .ZN(O9717));
  NOR2X1 G264 (.A1(W6195), .A2(I1473), .ZN(W12208));
  NOR2X1 G265 (.A1(I405), .A2(W2118), .ZN(O9705));
  NOR2X1 G266 (.A1(W4967), .A2(W27005), .ZN(O9708));
  NOR2X1 G267 (.A1(W11569), .A2(W14711), .ZN(O9713));
  NOR2X1 G268 (.A1(W31021), .A2(W15040), .ZN(W38663));
  NOR2X1 G269 (.A1(W1779), .A2(W329), .ZN(W38664));
  NOR2X1 G270 (.A1(W31965), .A2(W24028), .ZN(O9715));
  NOR2X1 G271 (.A1(W9020), .A2(I858), .ZN(W12201));
  NOR2X1 G272 (.A1(W2543), .A2(W8434), .ZN(W12400));
  NOR2X1 G273 (.A1(W18185), .A2(W9859), .ZN(W38669));
  NOR2X1 G274 (.A1(W16723), .A2(W385), .ZN(W21283));
  NOR2X1 G275 (.A1(W11894), .A2(W563), .ZN(W12196));
  NOR2X1 G276 (.A1(W6257), .A2(W20189), .ZN(W21284));
  NOR2X1 G277 (.A1(W14841), .A2(W37781), .ZN(O9720));
  NOR2X1 G278 (.A1(W9896), .A2(W30258), .ZN(W38674));
  NOR2X1 G279 (.A1(W16695), .A2(W20325), .ZN(W21286));
  NOR2X1 G280 (.A1(W8700), .A2(I1001), .ZN(W21149));
  NOR2X1 G281 (.A1(W14724), .A2(W4593), .ZN(O4977));
  NOR2X1 G282 (.A1(W4419), .A2(W5060), .ZN(W12615));
  NOR2X1 G283 (.A1(W10317), .A2(W2928), .ZN(W12614));
  NOR2X1 G284 (.A1(W470), .A2(W10355), .ZN(W21145));
  NOR2X1 G285 (.A1(W22327), .A2(W1851), .ZN(W38218));
  NOR2X1 G286 (.A1(W6113), .A2(W9909), .ZN(W12610));
  NOR2X1 G287 (.A1(W6208), .A2(W4913), .ZN(W29616));
  NOR2X1 G288 (.A1(W29452), .A2(W37895), .ZN(O9443));
  NOR2X1 G289 (.A1(W19468), .A2(W20805), .ZN(W29620));
  NOR2X1 G290 (.A1(W5439), .A2(W31291), .ZN(O9444));
  NOR2X1 G291 (.A1(W4255), .A2(W5901), .ZN(W12604));
  NOR2X1 G292 (.A1(W17078), .A2(I135), .ZN(W38225));
  NOR2X1 G293 (.A1(W3398), .A2(W10704), .ZN(W21150));
  NOR2X1 G294 (.A1(W34480), .A2(W32280), .ZN(O9445));
  NOR2X1 G295 (.A1(W19461), .A2(W14143), .ZN(O9447));
  NOR2X1 G296 (.A1(W9577), .A2(I1121), .ZN(W12598));
  NOR2X1 G297 (.A1(W9036), .A2(W3323), .ZN(O620));
  NOR2X1 G298 (.A1(W9013), .A2(I811), .ZN(W38205));
  NOR2X1 G299 (.A1(W1276), .A2(W15917), .ZN(O9431));
  NOR2X1 G300 (.A1(I255), .A2(W21255), .ZN(O4978));
  NOR2X1 G301 (.A1(W2992), .A2(W2363), .ZN(W12631));
  NOR2X1 G302 (.A1(W6085), .A2(W2265), .ZN(W21141));
  NOR2X1 G303 (.A1(W5027), .A2(W10953), .ZN(W12629));
  NOR2X1 G304 (.A1(W6521), .A2(W7764), .ZN(W12628));
  NOR2X1 G305 (.A1(W18548), .A2(W28611), .ZN(O9434));
  NOR2X1 G306 (.A1(W6030), .A2(I528), .ZN(W12626));
  NOR2X1 G307 (.A1(W24910), .A2(W979), .ZN(O4973));
  NOR2X1 G308 (.A1(W4892), .A2(W10064), .ZN(O624));
  NOR2X1 G309 (.A1(W23838), .A2(W5362), .ZN(W29622));
  NOR2X1 G310 (.A1(W29998), .A2(W11273), .ZN(O9436));
  NOR2X1 G311 (.A1(I873), .A2(W2378), .ZN(W12621));
  NOR2X1 G312 (.A1(W5197), .A2(W32629), .ZN(O9437));
  NOR2X1 G313 (.A1(W17790), .A2(W34684), .ZN(O9438));
  NOR2X1 G314 (.A1(W10689), .A2(I562), .ZN(W12618));
  NOR2X1 G315 (.A1(W5255), .A2(W12009), .ZN(O614));
  NOR2X1 G316 (.A1(W28096), .A2(I1003), .ZN(W38251));
  NOR2X1 G317 (.A1(W37006), .A2(W4218), .ZN(W38252));
  NOR2X1 G318 (.A1(W2610), .A2(I1622), .ZN(W21158));
  NOR2X1 G319 (.A1(W20808), .A2(W16149), .ZN(O9464));
  NOR2X1 G320 (.A1(W18493), .A2(I995), .ZN(W38258));
  NOR2X1 G321 (.A1(W13817), .A2(W22153), .ZN(W38260));
  NOR2X1 G322 (.A1(W28015), .A2(W34812), .ZN(O9466));
  NOR2X1 G323 (.A1(W4485), .A2(W3120), .ZN(W21159));
  NOR2X1 G324 (.A1(W37810), .A2(W11697), .ZN(O9462));
  NOR2X1 G325 (.A1(W2889), .A2(W1022), .ZN(W12566));
  NOR2X1 G326 (.A1(W5903), .A2(W145), .ZN(W21160));
  NOR2X1 G327 (.A1(I353), .A2(W13190), .ZN(W38265));
  NOR2X1 G328 (.A1(W29015), .A2(W7200), .ZN(O9469));
  NOR2X1 G329 (.A1(W9058), .A2(W16654), .ZN(W38267));
  NOR2X1 G330 (.A1(W16173), .A2(W26994), .ZN(O9470));
  NOR2X1 G331 (.A1(W4392), .A2(W12421), .ZN(O9471));
  NOR2X1 G332 (.A1(W10278), .A2(W9017), .ZN(W12559));
  NOR2X1 G333 (.A1(W5140), .A2(I1934), .ZN(W12587));
  NOR2X1 G334 (.A1(W13458), .A2(W24227), .ZN(W38231));
  NOR2X1 G335 (.A1(W11069), .A2(I915), .ZN(W12594));
  NOR2X1 G336 (.A1(W24870), .A2(W21486), .ZN(O9449));
  NOR2X1 G337 (.A1(W7197), .A2(W7470), .ZN(W29612));
  NOR2X1 G338 (.A1(W4281), .A2(W10674), .ZN(W12591));
  NOR2X1 G339 (.A1(W29466), .A2(W10947), .ZN(O9452));
  NOR2X1 G340 (.A1(W695), .A2(I812), .ZN(W12589));
  NOR2X1 G341 (.A1(W14735), .A2(W10710), .ZN(O9453));
  NOR2X1 G342 (.A1(W8596), .A2(W32771), .ZN(W38199));
  NOR2X1 G343 (.A1(W17235), .A2(W14375), .ZN(W29611));
  NOR2X1 G344 (.A1(W12268), .A2(W30479), .ZN(W38240));
  NOR2X1 G345 (.A1(I895), .A2(W2060), .ZN(W12584));
  NOR2X1 G346 (.A1(W22956), .A2(W30276), .ZN(W38241));
  NOR2X1 G347 (.A1(W16630), .A2(W1569), .ZN(O9457));
  NOR2X1 G348 (.A1(I315), .A2(W35459), .ZN(O9458));
  NOR2X1 G349 (.A1(W1162), .A2(W2824), .ZN(W12578));
  NOR2X1 G350 (.A1(W4866), .A2(W13297), .ZN(W38135));
  NOR2X1 G351 (.A1(W16745), .A2(W32266), .ZN(O9389));
  NOR2X1 G352 (.A1(W17878), .A2(W6115), .ZN(W38123));
  NOR2X1 G353 (.A1(W11922), .A2(W11008), .ZN(W12692));
  NOR2X1 G354 (.A1(W27179), .A2(W37071), .ZN(O9390));
  NOR2X1 G355 (.A1(W28012), .A2(W8818), .ZN(O4986));
  NOR2X1 G356 (.A1(W2187), .A2(W31624), .ZN(O9392));
  NOR2X1 G357 (.A1(W7791), .A2(W5660), .ZN(W12687));
  NOR2X1 G358 (.A1(W29526), .A2(W24083), .ZN(W38132));
  NOR2X1 G359 (.A1(W10508), .A2(I388), .ZN(W12695));
  NOR2X1 G360 (.A1(W29261), .A2(W2927), .ZN(W38139));
  NOR2X1 G361 (.A1(W11788), .A2(W7549), .ZN(W12683));
  NOR2X1 G362 (.A1(W25795), .A2(W29612), .ZN(O4985));
  NOR2X1 G363 (.A1(W11246), .A2(W14421), .ZN(O9399));
  NOR2X1 G364 (.A1(W31293), .A2(W30692), .ZN(W38152));
  NOR2X1 G365 (.A1(W2106), .A2(W1332), .ZN(O633));
  NOR2X1 G366 (.A1(W5778), .A2(W24086), .ZN(W29641));
  NOR2X1 G367 (.A1(W22793), .A2(W33024), .ZN(O9407));
  NOR2X1 G368 (.A1(W6363), .A2(W3275), .ZN(W12704));
  NOR2X1 G369 (.A1(W9675), .A2(W17269), .ZN(O9379));
  NOR2X1 G370 (.A1(W4931), .A2(W6090), .ZN(W12711));
  NOR2X1 G371 (.A1(W6828), .A2(W4886), .ZN(W12710));
  NOR2X1 G372 (.A1(I1927), .A2(I443), .ZN(W21117));
  NOR2X1 G373 (.A1(W1405), .A2(W26558), .ZN(W38110));
  NOR2X1 G374 (.A1(W22620), .A2(W34106), .ZN(O9381));
  NOR2X1 G375 (.A1(W2623), .A2(W11133), .ZN(W12706));
  NOR2X1 G376 (.A1(W9742), .A2(W565), .ZN(W12705));
  NOR2X1 G377 (.A1(W12560), .A2(W5193), .ZN(W12675));
  NOR2X1 G378 (.A1(W3829), .A2(W11327), .ZN(W12703));
  NOR2X1 G379 (.A1(W9616), .A2(W5655), .ZN(O9382));
  NOR2X1 G380 (.A1(W2878), .A2(W10216), .ZN(W12701));
  NOR2X1 G381 (.A1(W3733), .A2(W11996), .ZN(W21118));
  NOR2X1 G382 (.A1(W4056), .A2(W3362), .ZN(W12699));
  NOR2X1 G383 (.A1(W20167), .A2(W29779), .ZN(O9387));
  NOR2X1 G384 (.A1(W956), .A2(W26263), .ZN(W29647));
  NOR2X1 G385 (.A1(I531), .A2(I1748), .ZN(O4980));
  NOR2X1 G386 (.A1(W10420), .A2(W8661), .ZN(W12653));
  NOR2X1 G387 (.A1(I549), .A2(W17402), .ZN(W38177));
  NOR2X1 G388 (.A1(W37815), .A2(W4665), .ZN(W38180));
  NOR2X1 G389 (.A1(W8383), .A2(W172), .ZN(O4982));
  NOR2X1 G390 (.A1(W4364), .A2(W1018), .ZN(W12649));
  NOR2X1 G391 (.A1(W19232), .A2(W16231), .ZN(O9422));
  NOR2X1 G392 (.A1(W1415), .A2(W10056), .ZN(W12647));
  NOR2X1 G393 (.A1(W15504), .A2(W7244), .ZN(O2156));
  NOR2X1 G394 (.A1(W33041), .A2(W27267), .ZN(O9420));
  NOR2X1 G395 (.A1(W12912), .A2(W28302), .ZN(W29626));
  NOR2X1 G396 (.A1(W8704), .A2(W28578), .ZN(O9425));
  NOR2X1 G397 (.A1(W9049), .A2(W3260), .ZN(W12640));
  NOR2X1 G398 (.A1(W8485), .A2(W4170), .ZN(O2158));
  NOR2X1 G399 (.A1(W24353), .A2(W32778), .ZN(O9428));
  NOR2X1 G400 (.A1(W2514), .A2(W4014), .ZN(W29624));
  NOR2X1 G401 (.A1(W17743), .A2(W17717), .ZN(W38197));
  NOR2X1 G402 (.A1(W293), .A2(W12164), .ZN(O9430));
  NOR2X1 G403 (.A1(W24676), .A2(W35070), .ZN(O9416));
  NOR2X1 G404 (.A1(W4143), .A2(W1677), .ZN(W12674));
  NOR2X1 G405 (.A1(W4592), .A2(W6682), .ZN(W12673));
  NOR2X1 G406 (.A1(W36011), .A2(W26607), .ZN(W38157));
  NOR2X1 G407 (.A1(W9836), .A2(W20152), .ZN(W29640));
  NOR2X1 G408 (.A1(W4084), .A2(I1045), .ZN(O9412));
  NOR2X1 G409 (.A1(W16576), .A2(W4214), .ZN(O9413));
  NOR2X1 G410 (.A1(W26376), .A2(W11315), .ZN(O9414));
  NOR2X1 G411 (.A1(W6197), .A2(W9195), .ZN(W12666));
  NOR2X1 G412 (.A1(W19817), .A2(W27421), .ZN(W38270));
  NOR2X1 G413 (.A1(W8023), .A2(W3284), .ZN(O629));
  NOR2X1 G414 (.A1(W1782), .A2(W2824), .ZN(W12662));
  NOR2X1 G415 (.A1(W35348), .A2(W2093), .ZN(W38170));
  NOR2X1 G416 (.A1(W18661), .A2(W20176), .ZN(W21129));
  NOR2X1 G417 (.A1(W9769), .A2(W1615), .ZN(W12658));
  NOR2X1 G418 (.A1(W3196), .A2(W9816), .ZN(O9419));
  NOR2X1 G419 (.A1(W4969), .A2(W3331), .ZN(W12655));
  NOR2X1 G420 (.A1(W3568), .A2(W7201), .ZN(W12448));
  NOR2X1 G421 (.A1(W1037), .A2(W13284), .ZN(O4952));
  NOR2X1 G422 (.A1(W3575), .A2(I825), .ZN(O4951));
  NOR2X1 G423 (.A1(W12650), .A2(W20086), .ZN(W38382));
  NOR2X1 G424 (.A1(W12038), .A2(W9781), .ZN(W12455));
  NOR2X1 G425 (.A1(W7791), .A2(W14443), .ZN(W29561));
  NOR2X1 G426 (.A1(W9127), .A2(I1671), .ZN(W12452));
  NOR2X1 G427 (.A1(W12674), .A2(W10231), .ZN(O9540));
  NOR2X1 G428 (.A1(W22186), .A2(W27809), .ZN(O9542));
  NOR2X1 G429 (.A1(I60), .A2(W1106), .ZN(O9533));
  NOR2X1 G430 (.A1(W20101), .A2(W4277), .ZN(W21203));
  NOR2X1 G431 (.A1(W4209), .A2(W9502), .ZN(W12446));
  NOR2X1 G432 (.A1(W2567), .A2(W7826), .ZN(W12445));
  NOR2X1 G433 (.A1(W14123), .A2(W16889), .ZN(O2181));
  NOR2X1 G434 (.A1(W27318), .A2(W32125), .ZN(W38398));
  NOR2X1 G435 (.A1(W1938), .A2(W2706), .ZN(W12442));
  NOR2X1 G436 (.A1(W3543), .A2(I1414), .ZN(W12440));
  NOR2X1 G437 (.A1(W5640), .A2(W10280), .ZN(O4949));
  NOR2X1 G438 (.A1(W25473), .A2(W22282), .ZN(O9529));
  NOR2X1 G439 (.A1(W29688), .A2(W13060), .ZN(W38360));
  NOR2X1 G440 (.A1(W33598), .A2(W17851), .ZN(W38361));
  NOR2X1 G441 (.A1(W6412), .A2(W6134), .ZN(W12473));
  NOR2X1 G442 (.A1(W5754), .A2(W8706), .ZN(W12472));
  NOR2X1 G443 (.A1(W13132), .A2(W2744), .ZN(O4954));
  NOR2X1 G444 (.A1(W160), .A2(W19159), .ZN(O9526));
  NOR2X1 G445 (.A1(W8449), .A2(W9840), .ZN(W12469));
  NOR2X1 G446 (.A1(I1663), .A2(W35423), .ZN(O9528));
  NOR2X1 G447 (.A1(W7452), .A2(W11604), .ZN(W12438));
  NOR2X1 G448 (.A1(W9886), .A2(W8136), .ZN(W38369));
  NOR2X1 G449 (.A1(W276), .A2(W8420), .ZN(W12465));
  NOR2X1 G450 (.A1(W4735), .A2(I1779), .ZN(O603));
  NOR2X1 G451 (.A1(W13411), .A2(W2824), .ZN(W21196));
  NOR2X1 G452 (.A1(W23176), .A2(W16216), .ZN(W38374));
  NOR2X1 G453 (.A1(W34863), .A2(W20515), .ZN(W38375));
  NOR2X1 G454 (.A1(W14344), .A2(W357), .ZN(O2180));
  NOR2X1 G455 (.A1(W7120), .A2(W4784), .ZN(W12410));
  NOR2X1 G456 (.A1(W11628), .A2(W10203), .ZN(W12419));
  NOR2X1 G457 (.A1(W10047), .A2(W5247), .ZN(W12418));
  NOR2X1 G458 (.A1(W8834), .A2(I496), .ZN(W12417));
  NOR2X1 G459 (.A1(W8038), .A2(W7692), .ZN(W12415));
  NOR2X1 G460 (.A1(W16386), .A2(W9144), .ZN(W21216));
  NOR2X1 G461 (.A1(W12254), .A2(W12083), .ZN(W12413));
  NOR2X1 G462 (.A1(W7071), .A2(W25937), .ZN(O9567));
  NOR2X1 G463 (.A1(W37281), .A2(W25063), .ZN(O9568));
  NOR2X1 G464 (.A1(W5450), .A2(W6848), .ZN(W21214));
  NOR2X1 G465 (.A1(W9247), .A2(W8224), .ZN(O599));
  NOR2X1 G466 (.A1(W9582), .A2(I1090), .ZN(W12408));
  NOR2X1 G467 (.A1(W14020), .A2(W6323), .ZN(O9570));
  NOR2X1 G468 (.A1(W19873), .A2(W8089), .ZN(O9572));
  NOR2X1 G469 (.A1(W13588), .A2(W12028), .ZN(O4946));
  NOR2X1 G470 (.A1(W7551), .A2(W6614), .ZN(W21218));
  NOR2X1 G471 (.A1(W7443), .A2(W10175), .ZN(W12403));
  NOR2X1 G472 (.A1(I1455), .A2(W180), .ZN(O598));
  NOR2X1 G473 (.A1(W28698), .A2(W28328), .ZN(O9558));
  NOR2X1 G474 (.A1(W29180), .A2(W32494), .ZN(O9550));
  NOR2X1 G475 (.A1(W3348), .A2(W356), .ZN(W12436));
  NOR2X1 G476 (.A1(W1368), .A2(W164), .ZN(W12435));
  NOR2X1 G477 (.A1(W2336), .A2(W11605), .ZN(O4948));
  NOR2X1 G478 (.A1(W17699), .A2(W17702), .ZN(O9556));
  NOR2X1 G479 (.A1(W21404), .A2(W23033), .ZN(W29553));
  NOR2X1 G480 (.A1(W3554), .A2(I1709), .ZN(W12431));
  NOR2X1 G481 (.A1(W1365), .A2(W7451), .ZN(W12429));
  NOR2X1 G482 (.A1(W8790), .A2(W7256), .ZN(W29567));
  NOR2X1 G483 (.A1(W11656), .A2(W2165), .ZN(W29550));
  NOR2X1 G484 (.A1(W3586), .A2(W10583), .ZN(W21211));
  NOR2X1 G485 (.A1(W11441), .A2(W491), .ZN(W12425));
  NOR2X1 G486 (.A1(I1282), .A2(W3985), .ZN(W21212));
  NOR2X1 G487 (.A1(W34794), .A2(W24535), .ZN(O9561));
  NOR2X1 G488 (.A1(W11437), .A2(W12927), .ZN(W29548));
  NOR2X1 G489 (.A1(W1323), .A2(W1759), .ZN(W12421));
  NOR2X1 G490 (.A1(W11070), .A2(W1430), .ZN(W12529));
  NOR2X1 G491 (.A1(W21993), .A2(W5170), .ZN(W29596));
  NOR2X1 G492 (.A1(W20462), .A2(W13398), .ZN(W29594));
  NOR2X1 G493 (.A1(W8862), .A2(W3969), .ZN(O608));
  NOR2X1 G494 (.A1(W5953), .A2(W13651), .ZN(O2170));
  NOR2X1 G495 (.A1(W12141), .A2(W37710), .ZN(W38300));
  NOR2X1 G496 (.A1(W14104), .A2(W3995), .ZN(O4961));
  NOR2X1 G497 (.A1(W1728), .A2(W1136), .ZN(W12531));
  NOR2X1 G498 (.A1(W4918), .A2(W2687), .ZN(W12530));
  NOR2X1 G499 (.A1(W32866), .A2(I1488), .ZN(O9483));
  NOR2X1 G500 (.A1(W6490), .A2(W18171), .ZN(W21174));
  NOR2X1 G501 (.A1(W12356), .A2(W10964), .ZN(W38305));
  NOR2X1 G502 (.A1(W23188), .A2(W32904), .ZN(W38308));
  NOR2X1 G503 (.A1(W9170), .A2(W7647), .ZN(W12525));
  NOR2X1 G504 (.A1(W37147), .A2(W11330), .ZN(O9496));
  NOR2X1 G505 (.A1(W262), .A2(W6282), .ZN(O607));
  NOR2X1 G506 (.A1(W16907), .A2(W17583), .ZN(W38310));
  NOR2X1 G507 (.A1(W13907), .A2(W9239), .ZN(W21175));
  NOR2X1 G508 (.A1(W5271), .A2(W16385), .ZN(W21164));
  NOR2X1 G509 (.A1(W5924), .A2(W11085), .ZN(O611));
  NOR2X1 G510 (.A1(W7129), .A2(W9588), .ZN(W12555));
  NOR2X1 G511 (.A1(W15751), .A2(W16401), .ZN(W38272));
  NOR2X1 G512 (.A1(W18116), .A2(W26532), .ZN(O9472));
  NOR2X1 G513 (.A1(W19167), .A2(W34356), .ZN(W38275));
  NOR2X1 G514 (.A1(W2330), .A2(I776), .ZN(O4966));
  NOR2X1 G515 (.A1(W4178), .A2(W15322), .ZN(O2166));
  NOR2X1 G516 (.A1(I1289), .A2(W5394), .ZN(O9475));
  NOR2X1 G517 (.A1(W9012), .A2(W36427), .ZN(O9499));
  NOR2X1 G518 (.A1(I777), .A2(I1900), .ZN(W12547));
  NOR2X1 G519 (.A1(W8547), .A2(W23644), .ZN(W29601));
  NOR2X1 G520 (.A1(W1386), .A2(W842), .ZN(W12545));
  NOR2X1 G521 (.A1(W5944), .A2(W2337), .ZN(W29600));
  NOR2X1 G522 (.A1(W898), .A2(W15516), .ZN(O9479));
  NOR2X1 G523 (.A1(W7592), .A2(W7400), .ZN(O4965));
  NOR2X1 G524 (.A1(I39), .A2(I984), .ZN(W12541));
  NOR2X1 G525 (.A1(W3159), .A2(W11171), .ZN(W12486));
  NOR2X1 G526 (.A1(W11021), .A2(I876), .ZN(W12495));
  NOR2X1 G527 (.A1(W10495), .A2(W5902), .ZN(W12494));
  NOR2X1 G528 (.A1(W4343), .A2(W2356), .ZN(W29574));
  NOR2X1 G529 (.A1(W4875), .A2(W6233), .ZN(W12492));
  NOR2X1 G530 (.A1(W3583), .A2(W675), .ZN(O2174));
  NOR2X1 G531 (.A1(W4391), .A2(I986), .ZN(W12490));
  NOR2X1 G532 (.A1(W10634), .A2(W3368), .ZN(W12488));
  NOR2X1 G533 (.A1(W1852), .A2(W9434), .ZN(O604));
  NOR2X1 G534 (.A1(W15697), .A2(W20195), .ZN(W29577));
  NOR2X1 G535 (.A1(W4048), .A2(W28485), .ZN(O9519));
  NOR2X1 G536 (.A1(W1428), .A2(W906), .ZN(O2175));
  NOR2X1 G537 (.A1(W29180), .A2(W15167), .ZN(O4956));
  NOR2X1 G538 (.A1(W15878), .A2(W2808), .ZN(O2177));
  NOR2X1 G539 (.A1(W8144), .A2(W12037), .ZN(W12481));
  NOR2X1 G540 (.A1(W983), .A2(W4100), .ZN(W21191));
  NOR2X1 G541 (.A1(W3343), .A2(W2841), .ZN(O9520));
  NOR2X1 G542 (.A1(W16627), .A2(W7928), .ZN(W29569));
  NOR2X1 G543 (.A1(W15795), .A2(W20386), .ZN(W38329));
  NOR2X1 G544 (.A1(W6918), .A2(W1311), .ZN(O606));
  NOR2X1 G545 (.A1(W10806), .A2(W4973), .ZN(W12517));
  NOR2X1 G546 (.A1(W11340), .A2(I1005), .ZN(W12516));
  NOR2X1 G547 (.A1(W3434), .A2(W8699), .ZN(W12514));
  NOR2X1 G548 (.A1(W2481), .A2(W28300), .ZN(O9503));
  NOR2X1 G549 (.A1(W11423), .A2(W10159), .ZN(O4959));
  NOR2X1 G550 (.A1(W24358), .A2(W30718), .ZN(W38321));
  NOR2X1 G551 (.A1(W27417), .A2(W15250), .ZN(W38323));
  NOR2X1 G552 (.A1(W21062), .A2(W3363), .ZN(O9773));
  NOR2X1 G553 (.A1(W995), .A2(W2684), .ZN(O9511));
  NOR2X1 G554 (.A1(W9972), .A2(W37012), .ZN(O9512));
  NOR2X1 G555 (.A1(W21693), .A2(W27784), .ZN(O9513));
  NOR2X1 G556 (.A1(I1048), .A2(W3856), .ZN(W12500));
  NOR2X1 G557 (.A1(W30600), .A2(W13992), .ZN(W38337));
  NOR2X1 G558 (.A1(W31830), .A2(W5598), .ZN(W38338));
  NOR2X1 G559 (.A1(W2159), .A2(W8997), .ZN(O9516));
  NOR2X1 G560 (.A1(W8806), .A2(W28878), .ZN(O4823));
  NOR2X1 G561 (.A1(W1596), .A2(W35851), .ZN(O10029));
  NOR2X1 G562 (.A1(W21093), .A2(W27183), .ZN(W29308));
  NOR2X1 G563 (.A1(W6178), .A2(W8737), .ZN(W11675));
  NOR2X1 G564 (.A1(W2722), .A2(W17558), .ZN(O2252));
  NOR2X1 G565 (.A1(W11361), .A2(W6543), .ZN(O530));
  NOR2X1 G566 (.A1(W8448), .A2(W38082), .ZN(O10031));
  NOR2X1 G567 (.A1(W6145), .A2(W12001), .ZN(O10032));
  NOR2X1 G568 (.A1(W1331), .A2(W28459), .ZN(O4824));
  NOR2X1 G569 (.A1(W10583), .A2(W6302), .ZN(W11678));
  NOR2X1 G570 (.A1(W9524), .A2(W32078), .ZN(W39184));
  NOR2X1 G571 (.A1(W38979), .A2(W36191), .ZN(O10035));
  NOR2X1 G572 (.A1(W3598), .A2(W2656), .ZN(W11666));
  NOR2X1 G573 (.A1(W27314), .A2(W11056), .ZN(W39186));
  NOR2X1 G574 (.A1(W11172), .A2(W9996), .ZN(O10036));
  NOR2X1 G575 (.A1(I1300), .A2(I339), .ZN(W11663));
  NOR2X1 G576 (.A1(W4867), .A2(W3991), .ZN(W11662));
  NOR2X1 G577 (.A1(W36931), .A2(I18), .ZN(W39188));
  NOR2X1 G578 (.A1(W16450), .A2(W17546), .ZN(W39161));
  NOR2X1 G579 (.A1(W8108), .A2(W1763), .ZN(W11697));
  NOR2X1 G580 (.A1(W12452), .A2(W18990), .ZN(O10014));
  NOR2X1 G581 (.A1(W6462), .A2(W2515), .ZN(W21464));
  NOR2X1 G582 (.A1(W11566), .A2(W7185), .ZN(W11694));
  NOR2X1 G583 (.A1(W6278), .A2(W2578), .ZN(W11693));
  NOR2X1 G584 (.A1(W3170), .A2(W8333), .ZN(W11692));
  NOR2X1 G585 (.A1(W24199), .A2(W8906), .ZN(W29315));
  NOR2X1 G586 (.A1(W105), .A2(W8343), .ZN(O531));
  NOR2X1 G587 (.A1(W10362), .A2(W6318), .ZN(W11660));
  NOR2X1 G588 (.A1(W12116), .A2(W6138), .ZN(O4828));
  NOR2X1 G589 (.A1(W5035), .A2(W22543), .ZN(O10025));
  NOR2X1 G590 (.A1(W639), .A2(W15), .ZN(W11683));
  NOR2X1 G591 (.A1(W4820), .A2(W11353), .ZN(O4827));
  NOR2X1 G592 (.A1(W11417), .A2(W3322), .ZN(W11681));
  NOR2X1 G593 (.A1(W6347), .A2(I1707), .ZN(W11680));
  NOR2X1 G594 (.A1(W38444), .A2(W2981), .ZN(O10027));
  NOR2X1 G595 (.A1(W34696), .A2(W18215), .ZN(O10052));
  NOR2X1 G596 (.A1(W1366), .A2(W1026), .ZN(W11641));
  NOR2X1 G597 (.A1(W9383), .A2(W3826), .ZN(W11640));
  NOR2X1 G598 (.A1(W9009), .A2(W29748), .ZN(O10047));
  NOR2X1 G599 (.A1(W4713), .A2(W1762), .ZN(W11638));
  NOR2X1 G600 (.A1(W11752), .A2(W7459), .ZN(O2254));
  NOR2X1 G601 (.A1(W28445), .A2(W22711), .ZN(O10049));
  NOR2X1 G602 (.A1(I619), .A2(W1837), .ZN(W11635));
  NOR2X1 G603 (.A1(W10719), .A2(W21211), .ZN(W29298));
  NOR2X1 G604 (.A1(W3448), .A2(W1595), .ZN(O526));
  NOR2X1 G605 (.A1(W12779), .A2(W23751), .ZN(O10055));
  NOR2X1 G606 (.A1(W16731), .A2(W8825), .ZN(W29297));
  NOR2X1 G607 (.A1(W30115), .A2(W25901), .ZN(W39215));
  NOR2X1 G608 (.A1(W3512), .A2(W5937), .ZN(W11628));
  NOR2X1 G609 (.A1(W10318), .A2(W2808), .ZN(O4821));
  NOR2X1 G610 (.A1(W6302), .A2(W28920), .ZN(O10058));
  NOR2X1 G611 (.A1(W17481), .A2(W14817), .ZN(W39220));
  NOR2X1 G612 (.A1(W31283), .A2(W38037), .ZN(O10060));
  NOR2X1 G613 (.A1(W8406), .A2(W9544), .ZN(W39197));
  NOR2X1 G614 (.A1(W31881), .A2(W16655), .ZN(O10037));
  NOR2X1 G615 (.A1(W9616), .A2(W16705), .ZN(O10040));
  NOR2X1 G616 (.A1(W9202), .A2(W5161), .ZN(W11656));
  NOR2X1 G617 (.A1(W3798), .A2(W6151), .ZN(W29302));
  NOR2X1 G618 (.A1(W7510), .A2(W5932), .ZN(W21477));
  NOR2X1 G619 (.A1(W4133), .A2(W8036), .ZN(W11653));
  NOR2X1 G620 (.A1(W5240), .A2(W2907), .ZN(O4822));
  NOR2X1 G621 (.A1(W2692), .A2(W4481), .ZN(W11651));
  NOR2X1 G622 (.A1(I603), .A2(W35028), .ZN(W39157));
  NOR2X1 G623 (.A1(W3276), .A2(I291), .ZN(W11649));
  NOR2X1 G624 (.A1(W13171), .A2(W38698), .ZN(O10045));
  NOR2X1 G625 (.A1(W9690), .A2(W10469), .ZN(W11647));
  NOR2X1 G626 (.A1(W5197), .A2(W785), .ZN(W11646));
  NOR2X1 G627 (.A1(W9153), .A2(W7778), .ZN(W11645));
  NOR2X1 G628 (.A1(W10822), .A2(W306), .ZN(W11644));
  NOR2X1 G629 (.A1(W10012), .A2(I966), .ZN(W29299));
  NOR2X1 G630 (.A1(W30118), .A2(W21449), .ZN(O9976));
  NOR2X1 G631 (.A1(W4701), .A2(W4410), .ZN(W11758));
  NOR2X1 G632 (.A1(W21877), .A2(I829), .ZN(O4842));
  NOR2X1 G633 (.A1(W21001), .A2(W16386), .ZN(W21444));
  NOR2X1 G634 (.A1(W7643), .A2(W1112), .ZN(W11754));
  NOR2X1 G635 (.A1(W20704), .A2(W16602), .ZN(O9973));
  NOR2X1 G636 (.A1(W11070), .A2(W14569), .ZN(W39103));
  NOR2X1 G637 (.A1(W9028), .A2(W7030), .ZN(O535));
  NOR2X1 G638 (.A1(W4584), .A2(W3180), .ZN(W21445));
  NOR2X1 G639 (.A1(W3098), .A2(W2026), .ZN(W21441));
  NOR2X1 G640 (.A1(W10416), .A2(I1161), .ZN(W39107));
  NOR2X1 G641 (.A1(W38560), .A2(W1056), .ZN(W39108));
  NOR2X1 G642 (.A1(W21955), .A2(W36181), .ZN(O9977));
  NOR2X1 G643 (.A1(W9568), .A2(I1761), .ZN(W11745));
  NOR2X1 G644 (.A1(W8295), .A2(W10720), .ZN(W11744));
  NOR2X1 G645 (.A1(W35111), .A2(W22855), .ZN(O9978));
  NOR2X1 G646 (.A1(W13842), .A2(W28315), .ZN(O9981));
  NOR2X1 G647 (.A1(W33213), .A2(W5684), .ZN(O9982));
  NOR2X1 G648 (.A1(W7358), .A2(W4700), .ZN(W21434));
  NOR2X1 G649 (.A1(W2), .A2(W3097), .ZN(W11776));
  NOR2X1 G650 (.A1(W28928), .A2(W27649), .ZN(O9959));
  NOR2X1 G651 (.A1(W3814), .A2(W13479), .ZN(O4849));
  NOR2X1 G652 (.A1(W24142), .A2(W8584), .ZN(O4848));
  NOR2X1 G653 (.A1(W9903), .A2(W21746), .ZN(O9963));
  NOR2X1 G654 (.A1(W2894), .A2(W1011), .ZN(W11771));
  NOR2X1 G655 (.A1(W5159), .A2(W3008), .ZN(W11770));
  NOR2X1 G656 (.A1(W9842), .A2(W4124), .ZN(W11769));
  NOR2X1 G657 (.A1(W21850), .A2(W26520), .ZN(O4839));
  NOR2X1 G658 (.A1(W26213), .A2(W20142), .ZN(O4845));
  NOR2X1 G659 (.A1(W11639), .A2(W4232), .ZN(O4844));
  NOR2X1 G660 (.A1(I456), .A2(I1427), .ZN(W21438));
  NOR2X1 G661 (.A1(W37910), .A2(W34697), .ZN(O9966));
  NOR2X1 G662 (.A1(W3111), .A2(I1166), .ZN(O9967));
  NOR2X1 G663 (.A1(W10362), .A2(W12996), .ZN(O4843));
  NOR2X1 G664 (.A1(W20653), .A2(W20002), .ZN(W29340));
  NOR2X1 G665 (.A1(I1465), .A2(W1301), .ZN(W11709));
  NOR2X1 G666 (.A1(W17773), .A2(W8531), .ZN(W21456));
  NOR2X1 G667 (.A1(W3992), .A2(W11136), .ZN(O2248));
  NOR2X1 G668 (.A1(W27734), .A2(W25122), .ZN(O4834));
  NOR2X1 G669 (.A1(W1440), .A2(W21808), .ZN(W39142));
  NOR2X1 G670 (.A1(W5399), .A2(W26944), .ZN(W29322));
  NOR2X1 G671 (.A1(W37540), .A2(W3923), .ZN(W39146));
  NOR2X1 G672 (.A1(W5016), .A2(W3530), .ZN(O532));
  NOR2X1 G673 (.A1(W9302), .A2(W5752), .ZN(W11710));
  NOR2X1 G674 (.A1(W23396), .A2(W38012), .ZN(O9999));
  NOR2X1 G675 (.A1(W1057), .A2(W347), .ZN(W11707));
  NOR2X1 G676 (.A1(W7554), .A2(W6797), .ZN(W11706));
  NOR2X1 G677 (.A1(W16073), .A2(I263), .ZN(W21462));
  NOR2X1 G678 (.A1(W19020), .A2(W5437), .ZN(O10009));
  NOR2X1 G679 (.A1(W36770), .A2(W24104), .ZN(O10010));
  NOR2X1 G680 (.A1(W5619), .A2(W1649), .ZN(W11701));
  NOR2X1 G681 (.A1(I337), .A2(W16648), .ZN(O10013));
  NOR2X1 G682 (.A1(W6295), .A2(I1239), .ZN(W11699));
  NOR2X1 G683 (.A1(W11632), .A2(I1530), .ZN(W11730));
  NOR2X1 G684 (.A1(W8872), .A2(W20118), .ZN(W21448));
  NOR2X1 G685 (.A1(W10684), .A2(W5709), .ZN(W39120));
  NOR2X1 G686 (.A1(W0), .A2(I310), .ZN(W11736));
  NOR2X1 G687 (.A1(W17395), .A2(W35876), .ZN(O9988));
  NOR2X1 G688 (.A1(W19572), .A2(W19648), .ZN(W21449));
  NOR2X1 G689 (.A1(W27261), .A2(W17787), .ZN(W29332));
  NOR2X1 G690 (.A1(W28954), .A2(W27906), .ZN(W29331));
  NOR2X1 G691 (.A1(W9013), .A2(W31275), .ZN(O9992));
  NOR2X1 G692 (.A1(W18053), .A2(W20533), .ZN(O10062));
  NOR2X1 G693 (.A1(W9045), .A2(W32858), .ZN(W39127));
  NOR2X1 G694 (.A1(W23231), .A2(W8301), .ZN(O9993));
  NOR2X1 G695 (.A1(W5272), .A2(W22301), .ZN(O4837));
  NOR2X1 G696 (.A1(W1175), .A2(W32577), .ZN(O9995));
  NOR2X1 G697 (.A1(W35206), .A2(W20889), .ZN(W39133));
  NOR2X1 G698 (.A1(W25920), .A2(W6843), .ZN(O9997));
  NOR2X1 G699 (.A1(W7413), .A2(W10509), .ZN(W11722));
  NOR2X1 G700 (.A1(W17), .A2(W6376), .ZN(W11513));
  NOR2X1 G701 (.A1(W8004), .A2(W4680), .ZN(W11521));
  NOR2X1 G702 (.A1(W48), .A2(W2155), .ZN(W11520));
  NOR2X1 G703 (.A1(W6119), .A2(W34782), .ZN(W39323));
  NOR2X1 G704 (.A1(W16197), .A2(W11156), .ZN(O10126));
  NOR2X1 G705 (.A1(W2947), .A2(W50), .ZN(W11517));
  NOR2X1 G706 (.A1(W18096), .A2(W25414), .ZN(O4803));
  NOR2X1 G707 (.A1(W5455), .A2(W15654), .ZN(O2269));
  NOR2X1 G708 (.A1(W20361), .A2(W9135), .ZN(W29250));
  NOR2X1 G709 (.A1(W15970), .A2(W9478), .ZN(W39322));
  NOR2X1 G710 (.A1(W1540), .A2(W7041), .ZN(O10132));
  NOR2X1 G711 (.A1(W34871), .A2(W18601), .ZN(O10134));
  NOR2X1 G712 (.A1(W19022), .A2(W14533), .ZN(W21525));
  NOR2X1 G713 (.A1(W4541), .A2(W5405), .ZN(O4802));
  NOR2X1 G714 (.A1(W11060), .A2(W8540), .ZN(W11508));
  NOR2X1 G715 (.A1(W14631), .A2(W9785), .ZN(O2270));
  NOR2X1 G716 (.A1(W16889), .A2(W15492), .ZN(W21529));
  NOR2X1 G717 (.A1(W21375), .A2(W29822), .ZN(W39346));
  NOR2X1 G718 (.A1(I1480), .A2(W4055), .ZN(W11530));
  NOR2X1 G719 (.A1(W26909), .A2(W27375), .ZN(W39301));
  NOR2X1 G720 (.A1(W19663), .A2(W11528), .ZN(W21517));
  NOR2X1 G721 (.A1(W32911), .A2(W20741), .ZN(O10113));
  NOR2X1 G722 (.A1(W37898), .A2(W1998), .ZN(O10115));
  NOR2X1 G723 (.A1(I474), .A2(W1875), .ZN(W11535));
  NOR2X1 G724 (.A1(W3735), .A2(W11226), .ZN(W29257));
  NOR2X1 G725 (.A1(W5104), .A2(W5114), .ZN(W11533));
  NOR2X1 G726 (.A1(W8350), .A2(W158), .ZN(W11532));
  NOR2X1 G727 (.A1(W893), .A2(W160), .ZN(O10142));
  NOR2X1 G728 (.A1(W8832), .A2(W24928), .ZN(W39310));
  NOR2X1 G729 (.A1(W30953), .A2(W23030), .ZN(W39313));
  NOR2X1 G730 (.A1(W3061), .A2(W12577), .ZN(W39314));
  NOR2X1 G731 (.A1(W10281), .A2(W25746), .ZN(O4804));
  NOR2X1 G732 (.A1(W38921), .A2(I286), .ZN(W39319));
  NOR2X1 G733 (.A1(W7040), .A2(I410), .ZN(W11524));
  NOR2X1 G734 (.A1(W36428), .A2(W1586), .ZN(O10122));
  NOR2X1 G735 (.A1(W2831), .A2(W1896), .ZN(W11474));
  NOR2X1 G736 (.A1(W26410), .A2(W28554), .ZN(O10158));
  NOR2X1 G737 (.A1(W1553), .A2(I1272), .ZN(W11482));
  NOR2X1 G738 (.A1(W23103), .A2(W11894), .ZN(W29241));
  NOR2X1 G739 (.A1(I758), .A2(W11455), .ZN(O513));
  NOR2X1 G740 (.A1(W11375), .A2(W9314), .ZN(W11478));
  NOR2X1 G741 (.A1(I171), .A2(W551), .ZN(W11477));
  NOR2X1 G742 (.A1(W6017), .A2(W9536), .ZN(W11476));
  NOR2X1 G743 (.A1(W33080), .A2(W17527), .ZN(O10163));
  NOR2X1 G744 (.A1(W24377), .A2(W7691), .ZN(W39369));
  NOR2X1 G745 (.A1(W16247), .A2(W29363), .ZN(W39376));
  NOR2X1 G746 (.A1(W17913), .A2(W34632), .ZN(O10164));
  NOR2X1 G747 (.A1(W3129), .A2(W756), .ZN(W11471));
  NOR2X1 G748 (.A1(W11766), .A2(I1764), .ZN(W21539));
  NOR2X1 G749 (.A1(W7563), .A2(I481), .ZN(W11468));
  NOR2X1 G750 (.A1(W6565), .A2(W2271), .ZN(W11467));
  NOR2X1 G751 (.A1(W26826), .A2(W11306), .ZN(O10166));
  NOR2X1 G752 (.A1(W33482), .A2(W32430), .ZN(O10167));
  NOR2X1 G753 (.A1(W14035), .A2(W26880), .ZN(O10149));
  NOR2X1 G754 (.A1(W6273), .A2(W21386), .ZN(W21530));
  NOR2X1 G755 (.A1(W8596), .A2(I1770), .ZN(W21531));
  NOR2X1 G756 (.A1(W2350), .A2(W6894), .ZN(W11500));
  NOR2X1 G757 (.A1(W14570), .A2(W10193), .ZN(O2271));
  NOR2X1 G758 (.A1(W9574), .A2(W511), .ZN(W11498));
  NOR2X1 G759 (.A1(W8919), .A2(W29308), .ZN(O10146));
  NOR2X1 G760 (.A1(W16056), .A2(W26236), .ZN(W29243));
  NOR2X1 G761 (.A1(W10425), .A2(W533), .ZN(W11493));
  NOR2X1 G762 (.A1(W38170), .A2(W29154), .ZN(W39298));
  NOR2X1 G763 (.A1(W2650), .A2(W10071), .ZN(W11491));
  NOR2X1 G764 (.A1(W2879), .A2(W17621), .ZN(O10150));
  NOR2X1 G765 (.A1(W21588), .A2(W11036), .ZN(O10151));
  NOR2X1 G766 (.A1(W1785), .A2(W3444), .ZN(W11488));
  NOR2X1 G767 (.A1(W8765), .A2(W12230), .ZN(W21536));
  NOR2X1 G768 (.A1(W11865), .A2(W10579), .ZN(O10153));
  NOR2X1 G769 (.A1(W3057), .A2(W2985), .ZN(O10154));
  NOR2X1 G770 (.A1(W1627), .A2(W15169), .ZN(W21501));
  NOR2X1 G771 (.A1(I790), .A2(I1694), .ZN(W11601));
  NOR2X1 G772 (.A1(W20685), .A2(W23121), .ZN(O10082));
  NOR2X1 G773 (.A1(W2993), .A2(W551), .ZN(W21498));
  NOR2X1 G774 (.A1(W1819), .A2(W19360), .ZN(O10086));
  NOR2X1 G775 (.A1(I468), .A2(W8820), .ZN(O2261));
  NOR2X1 G776 (.A1(W11008), .A2(W10095), .ZN(W11594));
  NOR2X1 G777 (.A1(W32250), .A2(W8452), .ZN(O10087));
  NOR2X1 G778 (.A1(W400), .A2(W3593), .ZN(O522));
  NOR2X1 G779 (.A1(W25945), .A2(W7694), .ZN(O4814));
  NOR2X1 G780 (.A1(W10089), .A2(W442), .ZN(W11590));
  NOR2X1 G781 (.A1(W27232), .A2(W39024), .ZN(W39261));
  NOR2X1 G782 (.A1(W8755), .A2(W38418), .ZN(W39263));
  NOR2X1 G783 (.A1(W12582), .A2(W12099), .ZN(W29272));
  NOR2X1 G784 (.A1(W27264), .A2(W21920), .ZN(O10089));
  NOR2X1 G785 (.A1(W1600), .A2(W270), .ZN(W11584));
  NOR2X1 G786 (.A1(W22557), .A2(W10246), .ZN(O10090));
  NOR2X1 G787 (.A1(W2164), .A2(W921), .ZN(W11582));
  NOR2X1 G788 (.A1(W15948), .A2(W23002), .ZN(W39234));
  NOR2X1 G789 (.A1(W11439), .A2(W1256), .ZN(O4819));
  NOR2X1 G790 (.A1(W3151), .A2(W5823), .ZN(W11620));
  NOR2X1 G791 (.A1(W18593), .A2(W9527), .ZN(W39225));
  NOR2X1 G792 (.A1(I744), .A2(W397), .ZN(O4818));
  NOR2X1 G793 (.A1(W9389), .A2(W14196), .ZN(W29289));
  NOR2X1 G794 (.A1(W3582), .A2(I1766), .ZN(W11616));
  NOR2X1 G795 (.A1(W12768), .A2(W15399), .ZN(O10067));
  NOR2X1 G796 (.A1(W11451), .A2(W12016), .ZN(O2258));
  NOR2X1 G797 (.A1(W2449), .A2(W13087), .ZN(O4812));
  NOR2X1 G798 (.A1(W12964), .A2(W6439), .ZN(W21491));
  NOR2X1 G799 (.A1(W7537), .A2(W5428), .ZN(W11609));
  NOR2X1 G800 (.A1(W6970), .A2(W27661), .ZN(W29282));
  NOR2X1 G801 (.A1(W4794), .A2(W17366), .ZN(O4815));
  NOR2X1 G802 (.A1(W29072), .A2(W33511), .ZN(O10075));
  NOR2X1 G803 (.A1(I504), .A2(W1452), .ZN(O10076));
  NOR2X1 G804 (.A1(W3526), .A2(W37135), .ZN(O10079));
  NOR2X1 G805 (.A1(W1644), .A2(W10064), .ZN(W11552));
  NOR2X1 G806 (.A1(I994), .A2(W5935), .ZN(O521));
  NOR2X1 G807 (.A1(W8018), .A2(W4979), .ZN(O10101));
  NOR2X1 G808 (.A1(W26039), .A2(W38435), .ZN(W39286));
  NOR2X1 G809 (.A1(W1530), .A2(W1918), .ZN(W11559));
  NOR2X1 G810 (.A1(W6730), .A2(W3008), .ZN(W29264));
  NOR2X1 G811 (.A1(W6505), .A2(W5102), .ZN(W11555));
  NOR2X1 G812 (.A1(W14765), .A2(W33296), .ZN(O10103));
  NOR2X1 G813 (.A1(I1033), .A2(I1330), .ZN(W11553));
  NOR2X1 G814 (.A1(W2492), .A2(W220), .ZN(W11563));
  NOR2X1 G815 (.A1(W20384), .A2(W5917), .ZN(W39292));
  NOR2X1 G816 (.A1(W11331), .A2(W5504), .ZN(W11550));
  NOR2X1 G817 (.A1(I196), .A2(W8934), .ZN(O519));
  NOR2X1 G818 (.A1(W11647), .A2(W25133), .ZN(W39294));
  NOR2X1 G819 (.A1(W26926), .A2(W26721), .ZN(W29263));
  NOR2X1 G820 (.A1(W16905), .A2(W28918), .ZN(W29262));
  NOR2X1 G821 (.A1(W5958), .A2(W10129), .ZN(W11544));
  NOR2X1 G822 (.A1(W3464), .A2(W1129), .ZN(W11543));
  NOR2X1 G823 (.A1(W19242), .A2(W4271), .ZN(O4810));
  NOR2X1 G824 (.A1(W21347), .A2(W879), .ZN(O10092));
  NOR2X1 G825 (.A1(W1850), .A2(I750), .ZN(W11579));
  NOR2X1 G826 (.A1(W17933), .A2(W17389), .ZN(O10093));
  NOR2X1 G827 (.A1(W24000), .A2(W17922), .ZN(W39271));
  NOR2X1 G828 (.A1(W818), .A2(W11292), .ZN(W11576));
  NOR2X1 G829 (.A1(W17410), .A2(W5224), .ZN(O4811));
  NOR2X1 G830 (.A1(W10243), .A2(W1914), .ZN(W11574));
  NOR2X1 G831 (.A1(W29145), .A2(W28264), .ZN(W29269));
  NOR2X1 G832 (.A1(W24398), .A2(W36040), .ZN(W39078));
  NOR2X1 G833 (.A1(W9388), .A2(I1340), .ZN(W11571));
  NOR2X1 G834 (.A1(W5571), .A2(W11066), .ZN(W11570));
  NOR2X1 G835 (.A1(W20219), .A2(W19066), .ZN(W39279));
  NOR2X1 G836 (.A1(I1753), .A2(W731), .ZN(W11568));
  NOR2X1 G837 (.A1(W5342), .A2(W6747), .ZN(W11567));
  NOR2X1 G838 (.A1(W11964), .A2(W7648), .ZN(W39281));
  NOR2X1 G839 (.A1(W7575), .A2(W21436), .ZN(W21508));
  NOR2X1 G840 (.A1(W19574), .A2(W1016), .ZN(W38890));
  NOR2X1 G841 (.A1(W27372), .A2(W38411), .ZN(W38881));
  NOR2X1 G842 (.A1(W10237), .A2(W18522), .ZN(W21369));
  NOR2X1 G843 (.A1(W5387), .A2(W2202), .ZN(W11983));
  NOR2X1 G844 (.A1(W28584), .A2(W27056), .ZN(O9844));
  NOR2X1 G845 (.A1(W14132), .A2(W17401), .ZN(W29405));
  NOR2X1 G846 (.A1(I694), .A2(W10719), .ZN(W11980));
  NOR2X1 G847 (.A1(W3842), .A2(W12065), .ZN(W21373));
  NOR2X1 G848 (.A1(W4883), .A2(W5477), .ZN(W11976));
  NOR2X1 G849 (.A1(W12559), .A2(W12823), .ZN(O4877));
  NOR2X1 G850 (.A1(W30508), .A2(W576), .ZN(W38892));
  NOR2X1 G851 (.A1(W7824), .A2(W25645), .ZN(O4873));
  NOR2X1 G852 (.A1(W19901), .A2(W21392), .ZN(W38897));
  NOR2X1 G853 (.A1(W33559), .A2(W20468), .ZN(O9853));
  NOR2X1 G854 (.A1(W6476), .A2(W6682), .ZN(W11969));
  NOR2X1 G855 (.A1(W9576), .A2(W27859), .ZN(W38899));
  NOR2X1 G856 (.A1(W15408), .A2(W13876), .ZN(W29399));
  NOR2X1 G857 (.A1(W1218), .A2(W3374), .ZN(W11966));
  NOR2X1 G858 (.A1(I1312), .A2(W11233), .ZN(W11996));
  NOR2X1 G859 (.A1(W30343), .A2(W36869), .ZN(W38857));
  NOR2X1 G860 (.A1(W10868), .A2(W10503), .ZN(W21360));
  NOR2X1 G861 (.A1(W1023), .A2(W4084), .ZN(O557));
  NOR2X1 G862 (.A1(W19039), .A2(W9028), .ZN(W21362));
  NOR2X1 G863 (.A1(W32501), .A2(W5067), .ZN(O9835));
  NOR2X1 G864 (.A1(W9225), .A2(W5434), .ZN(W11999));
  NOR2X1 G865 (.A1(W3619), .A2(W9126), .ZN(W11998));
  NOR2X1 G866 (.A1(W9088), .A2(W25164), .ZN(O9838));
  NOR2X1 G867 (.A1(W8722), .A2(W10114), .ZN(O4872));
  NOR2X1 G868 (.A1(W14465), .A2(W20305), .ZN(W29416));
  NOR2X1 G869 (.A1(W7354), .A2(W36674), .ZN(W38870));
  NOR2X1 G870 (.A1(W7077), .A2(W23396), .ZN(O4880));
  NOR2X1 G871 (.A1(W15885), .A2(W23089), .ZN(O4879));
  NOR2X1 G872 (.A1(W10699), .A2(W23353), .ZN(O9841));
  NOR2X1 G873 (.A1(W37890), .A2(W10826), .ZN(W38876));
  NOR2X1 G874 (.A1(W31081), .A2(W33415), .ZN(W38877));
  NOR2X1 G875 (.A1(W26109), .A2(W6379), .ZN(O9873));
  NOR2X1 G876 (.A1(W15336), .A2(W20346), .ZN(O4869));
  NOR2X1 G877 (.A1(W19333), .A2(W19839), .ZN(O2230));
  NOR2X1 G878 (.A1(W2614), .A2(W37572), .ZN(O9866));
  NOR2X1 G879 (.A1(W15720), .A2(W16981), .ZN(O9868));
  NOR2X1 G880 (.A1(W1178), .A2(W33055), .ZN(O9870));
  NOR2X1 G881 (.A1(W12367), .A2(W8545), .ZN(O9871));
  NOR2X1 G882 (.A1(W17518), .A2(W6843), .ZN(O2231));
  NOR2X1 G883 (.A1(W123), .A2(W4070), .ZN(W11939));
  NOR2X1 G884 (.A1(W7423), .A2(W11597), .ZN(W11947));
  NOR2X1 G885 (.A1(W2215), .A2(W3916), .ZN(W11937));
  NOR2X1 G886 (.A1(W666), .A2(W35963), .ZN(O9876));
  NOR2X1 G887 (.A1(W8057), .A2(I448), .ZN(O550));
  NOR2X1 G888 (.A1(W2915), .A2(W800), .ZN(W21389));
  NOR2X1 G889 (.A1(W23898), .A2(W34874), .ZN(O9884));
  NOR2X1 G890 (.A1(W9185), .A2(W3804), .ZN(W11931));
  NOR2X1 G891 (.A1(W1242), .A2(I1216), .ZN(W11930));
  NOR2X1 G892 (.A1(W5364), .A2(W23840), .ZN(W38949));
  NOR2X1 G893 (.A1(W7344), .A2(W3902), .ZN(O9861));
  NOR2X1 G894 (.A1(W6242), .A2(W27992), .ZN(W29396));
  NOR2X1 G895 (.A1(W12356), .A2(W18483), .ZN(W38904));
  NOR2X1 G896 (.A1(W12897), .A2(W34362), .ZN(O9858));
  NOR2X1 G897 (.A1(W10547), .A2(W1110), .ZN(O552));
  NOR2X1 G898 (.A1(W14701), .A2(W6444), .ZN(W38906));
  NOR2X1 G899 (.A1(W4139), .A2(W8062), .ZN(W21379));
  NOR2X1 G900 (.A1(W25505), .A2(W18193), .ZN(W29394));
  NOR2X1 G901 (.A1(W17466), .A2(W10043), .ZN(W21381));
  NOR2X1 G902 (.A1(W8379), .A2(W36118), .ZN(O9830));
  NOR2X1 G903 (.A1(W11555), .A2(W8208), .ZN(W11954));
  NOR2X1 G904 (.A1(W3864), .A2(I868), .ZN(O4870));
  NOR2X1 G905 (.A1(W32507), .A2(W22921), .ZN(W38916));
  NOR2X1 G906 (.A1(W22798), .A2(W27482), .ZN(W38917));
  NOR2X1 G907 (.A1(W11170), .A2(W22616), .ZN(W29391));
  NOR2X1 G908 (.A1(I1069), .A2(W10620), .ZN(W11949));
  NOR2X1 G909 (.A1(W19022), .A2(W8809), .ZN(W21385));
  NOR2X1 G910 (.A1(I579), .A2(W247), .ZN(W12058));
  NOR2X1 G911 (.A1(W19874), .A2(W5490), .ZN(W38787));
  NOR2X1 G912 (.A1(W6088), .A2(W10750), .ZN(W12065));
  NOR2X1 G913 (.A1(W19077), .A2(I1270), .ZN(O4892));
  NOR2X1 G914 (.A1(I1993), .A2(W1190), .ZN(W21334));
  NOR2X1 G915 (.A1(W27986), .A2(W11130), .ZN(O9789));
  NOR2X1 G916 (.A1(W35903), .A2(W34408), .ZN(O9790));
  NOR2X1 G917 (.A1(W10991), .A2(I1138), .ZN(W12060));
  NOR2X1 G918 (.A1(W37515), .A2(W14566), .ZN(O9791));
  NOR2X1 G919 (.A1(W8677), .A2(W2083), .ZN(W12067));
  NOR2X1 G920 (.A1(W6641), .A2(W5979), .ZN(W12057));
  NOR2X1 G921 (.A1(W38251), .A2(W20270), .ZN(W38794));
  NOR2X1 G922 (.A1(W29297), .A2(W19681), .ZN(O9792));
  NOR2X1 G923 (.A1(W745), .A2(W17530), .ZN(O4891));
  NOR2X1 G924 (.A1(W851), .A2(W5899), .ZN(W12053));
  NOR2X1 G925 (.A1(W16470), .A2(W27523), .ZN(W29434));
  NOR2X1 G926 (.A1(I729), .A2(W2420), .ZN(W12051));
  NOR2X1 G927 (.A1(W27321), .A2(W32330), .ZN(O9798));
  NOR2X1 G928 (.A1(W24492), .A2(W17659), .ZN(W38771));
  NOR2X1 G929 (.A1(W858), .A2(W4368), .ZN(O4895));
  NOR2X1 G930 (.A1(W25033), .A2(W18366), .ZN(W38767));
  NOR2X1 G931 (.A1(W3746), .A2(W389), .ZN(W12084));
  NOR2X1 G932 (.A1(W3867), .A2(W11321), .ZN(W12083));
  NOR2X1 G933 (.A1(W3444), .A2(W10912), .ZN(W12081));
  NOR2X1 G934 (.A1(W1252), .A2(W3001), .ZN(W12080));
  NOR2X1 G935 (.A1(W6586), .A2(W2756), .ZN(W12079));
  NOR2X1 G936 (.A1(W1026), .A2(W10666), .ZN(O565));
  NOR2X1 G937 (.A1(I52), .A2(W11379), .ZN(W21337));
  NOR2X1 G938 (.A1(W22511), .A2(W6426), .ZN(O9779));
  NOR2X1 G939 (.A1(W9649), .A2(W16796), .ZN(W21329));
  NOR2X1 G940 (.A1(W6639), .A2(W4068), .ZN(W12073));
  NOR2X1 G941 (.A1(W489), .A2(W3829), .ZN(O4894));
  NOR2X1 G942 (.A1(W11211), .A2(W29601), .ZN(O9782));
  NOR2X1 G943 (.A1(W9049), .A2(W7253), .ZN(W21331));
  NOR2X1 G944 (.A1(W7883), .A2(W10753), .ZN(W12069));
  NOR2X1 G945 (.A1(W5508), .A2(W3903), .ZN(W12018));
  NOR2X1 G946 (.A1(W36772), .A2(W13637), .ZN(O9819));
  NOR2X1 G947 (.A1(W29308), .A2(W17646), .ZN(W38839));
  NOR2X1 G948 (.A1(W12161), .A2(I530), .ZN(O2221));
  NOR2X1 G949 (.A1(W9285), .A2(W28281), .ZN(O9822));
  NOR2X1 G950 (.A1(W6897), .A2(W906), .ZN(W12022));
  NOR2X1 G951 (.A1(W23717), .A2(W1635), .ZN(W29423));
  NOR2X1 G952 (.A1(I104), .A2(W8026), .ZN(O559));
  NOR2X1 G953 (.A1(W11900), .A2(W5162), .ZN(W12019));
  NOR2X1 G954 (.A1(W17164), .A2(W8001), .ZN(O9818));
  NOR2X1 G955 (.A1(W15599), .A2(W5574), .ZN(W21353));
  NOR2X1 G956 (.A1(W20054), .A2(W6937), .ZN(W21354));
  NOR2X1 G957 (.A1(W6507), .A2(W18106), .ZN(W29421));
  NOR2X1 G958 (.A1(W10475), .A2(I239), .ZN(W12013));
  NOR2X1 G959 (.A1(W12110), .A2(W2234), .ZN(W21357));
  NOR2X1 G960 (.A1(W33929), .A2(W16159), .ZN(W38852));
  NOR2X1 G961 (.A1(W8403), .A2(I463), .ZN(W12010));
  NOR2X1 G962 (.A1(W7105), .A2(W9003), .ZN(W12009));
  NOR2X1 G963 (.A1(W1481), .A2(W13005), .ZN(O2220));
  NOR2X1 G964 (.A1(W14577), .A2(W18517), .ZN(W21338));
  NOR2X1 G965 (.A1(W3447), .A2(I1719), .ZN(W12047));
  NOR2X1 G966 (.A1(W20443), .A2(W18020), .ZN(O4889));
  NOR2X1 G967 (.A1(W10706), .A2(W20064), .ZN(W21342));
  NOR2X1 G968 (.A1(W9753), .A2(W11276), .ZN(W21343));
  NOR2X1 G969 (.A1(W7557), .A2(W3888), .ZN(W12040));
  NOR2X1 G970 (.A1(W16390), .A2(W28491), .ZN(W38818));
  NOR2X1 G971 (.A1(W233), .A2(W6486), .ZN(W21345));
  NOR2X1 G972 (.A1(W16479), .A2(I919), .ZN(W21391));
  NOR2X1 G973 (.A1(W2340), .A2(W1865), .ZN(W12036));
  NOR2X1 G974 (.A1(W18047), .A2(W36841), .ZN(O9809));
  NOR2X1 G975 (.A1(W5889), .A2(W8510), .ZN(W21347));
  NOR2X1 G976 (.A1(W13723), .A2(W38067), .ZN(O9811));
  NOR2X1 G977 (.A1(W213), .A2(W10181), .ZN(W38828));
  NOR2X1 G978 (.A1(W26515), .A2(W3602), .ZN(O4886));
  NOR2X1 G979 (.A1(W16341), .A2(W5666), .ZN(O9817));
  NOR2X1 G980 (.A1(W2814), .A2(W8669), .ZN(W11825));
  NOR2X1 G981 (.A1(W4305), .A2(I1344), .ZN(W11833));
  NOR2X1 G982 (.A1(W3043), .A2(W1167), .ZN(W11832));
  NOR2X1 G983 (.A1(W7576), .A2(W2426), .ZN(W11831));
  NOR2X1 G984 (.A1(W7843), .A2(W8547), .ZN(W11830));
  NOR2X1 G985 (.A1(W6419), .A2(W1419), .ZN(W11829));
  NOR2X1 G986 (.A1(W2619), .A2(W3936), .ZN(W11828));
  NOR2X1 G987 (.A1(W1278), .A2(W3896), .ZN(W11827));
  NOR2X1 G988 (.A1(W33275), .A2(W6898), .ZN(W39039));
  NOR2X1 G989 (.A1(W27458), .A2(W22615), .ZN(O9933));
  NOR2X1 G990 (.A1(W28869), .A2(W38442), .ZN(O9935));
  NOR2X1 G991 (.A1(W3263), .A2(W9083), .ZN(O540));
  NOR2X1 G992 (.A1(W21196), .A2(I305), .ZN(O4856));
  NOR2X1 G993 (.A1(W30149), .A2(W24653), .ZN(W39045));
  NOR2X1 G994 (.A1(W2410), .A2(W10547), .ZN(W11819));
  NOR2X1 G995 (.A1(W11542), .A2(W9692), .ZN(W11818));
  NOR2X1 G996 (.A1(W6835), .A2(W7713), .ZN(W11817));
  NOR2X1 G997 (.A1(W15249), .A2(W1878), .ZN(W21419));
  NOR2X1 G998 (.A1(W26945), .A2(W25840), .ZN(W39031));
  NOR2X1 G999 (.A1(W15302), .A2(W33604), .ZN(W39022));
  NOR2X1 G1000 (.A1(W17394), .A2(W20102), .ZN(O4857));
  NOR2X1 G1001 (.A1(W5092), .A2(W10302), .ZN(O543));
  NOR2X1 G1002 (.A1(W2277), .A2(W6550), .ZN(W21413));
  NOR2X1 G1003 (.A1(W4960), .A2(W2568), .ZN(W39026));
  NOR2X1 G1004 (.A1(W7473), .A2(W9981), .ZN(W11846));
  NOR2X1 G1005 (.A1(W6386), .A2(W30824), .ZN(O9927));
  NOR2X1 G1006 (.A1(W9943), .A2(W9245), .ZN(W21414));
  NOR2X1 G1007 (.A1(W6609), .A2(W28784), .ZN(O9938));
  NOR2X1 G1008 (.A1(W38259), .A2(W7857), .ZN(O9931));
  NOR2X1 G1009 (.A1(W2398), .A2(W1642), .ZN(W11840));
  NOR2X1 G1010 (.A1(I447), .A2(W4933), .ZN(W11839));
  NOR2X1 G1011 (.A1(W1946), .A2(W9311), .ZN(W21416));
  NOR2X1 G1012 (.A1(W6905), .A2(W10846), .ZN(W11837));
  NOR2X1 G1013 (.A1(W16482), .A2(W33355), .ZN(W39036));
  NOR2X1 G1014 (.A1(W598), .A2(I1263), .ZN(O542));
  NOR2X1 G1015 (.A1(W37368), .A2(W8995), .ZN(W39070));
  NOR2X1 G1016 (.A1(W4850), .A2(W5699), .ZN(W11795));
  NOR2X1 G1017 (.A1(W12248), .A2(I587), .ZN(O9946));
  NOR2X1 G1018 (.A1(W5123), .A2(W37070), .ZN(O9947));
  NOR2X1 G1019 (.A1(W36347), .A2(W21719), .ZN(O9949));
  NOR2X1 G1020 (.A1(W29416), .A2(W15296), .ZN(O9950));
  NOR2X1 G1021 (.A1(W2867), .A2(W5018), .ZN(W11789));
  NOR2X1 G1022 (.A1(W4108), .A2(W20865), .ZN(O4852));
  NOR2X1 G1023 (.A1(I1209), .A2(W17779), .ZN(W21428));
  NOR2X1 G1024 (.A1(W12367), .A2(W20123), .ZN(W21425));
  NOR2X1 G1025 (.A1(W12056), .A2(W6619), .ZN(O4850));
  NOR2X1 G1026 (.A1(W8243), .A2(I1391), .ZN(W11784));
  NOR2X1 G1027 (.A1(W8383), .A2(W9399), .ZN(W11783));
  NOR2X1 G1028 (.A1(W7370), .A2(W6108), .ZN(W11782));
  NOR2X1 G1029 (.A1(W8317), .A2(W13477), .ZN(W21430));
  NOR2X1 G1030 (.A1(W34416), .A2(W5430), .ZN(O9955));
  NOR2X1 G1031 (.A1(W22856), .A2(W2483), .ZN(W39074));
  NOR2X1 G1032 (.A1(W16672), .A2(W20871), .ZN(W21431));
  NOR2X1 G1033 (.A1(W10275), .A2(W11211), .ZN(W11805));
  NOR2X1 G1034 (.A1(W19181), .A2(W17758), .ZN(W21421));
  NOR2X1 G1035 (.A1(I1572), .A2(I842), .ZN(W11812));
  NOR2X1 G1036 (.A1(W13880), .A2(W5099), .ZN(W21422));
  NOR2X1 G1037 (.A1(W9468), .A2(I36), .ZN(W11810));
  NOR2X1 G1038 (.A1(W11127), .A2(W10441), .ZN(W11809));
  NOR2X1 G1039 (.A1(W597), .A2(W9), .ZN(W11808));
  NOR2X1 G1040 (.A1(W13094), .A2(W18220), .ZN(W39053));
  NOR2X1 G1041 (.A1(W24202), .A2(W28411), .ZN(O9941));
  NOR2X1 G1042 (.A1(W11287), .A2(W23836), .ZN(W29362));
  NOR2X1 G1043 (.A1(W6880), .A2(W7321), .ZN(W11804));
  NOR2X1 G1044 (.A1(W16990), .A2(W18461), .ZN(W29355));
  NOR2X1 G1045 (.A1(W25410), .A2(W34343), .ZN(O9943));
  NOR2X1 G1046 (.A1(W6493), .A2(W858), .ZN(W11801));
  NOR2X1 G1047 (.A1(W6067), .A2(W2320), .ZN(W11800));
  NOR2X1 G1048 (.A1(W8912), .A2(W10248), .ZN(W11799));
  NOR2X1 G1049 (.A1(W2924), .A2(W3459), .ZN(W11797));
  NOR2X1 G1050 (.A1(W1373), .A2(W21770), .ZN(O9906));
  NOR2X1 G1051 (.A1(W2964), .A2(W9439), .ZN(O9898));
  NOR2X1 G1052 (.A1(W1279), .A2(W5370), .ZN(W11908));
  NOR2X1 G1053 (.A1(W17859), .A2(W12079), .ZN(O9899));
  NOR2X1 G1054 (.A1(W20209), .A2(W12234), .ZN(W21399));
  NOR2X1 G1055 (.A1(W11708), .A2(W5695), .ZN(W11905));
  NOR2X1 G1056 (.A1(W31103), .A2(I929), .ZN(O9902));
  NOR2X1 G1057 (.A1(W22884), .A2(I1620), .ZN(W38980));
  NOR2X1 G1058 (.A1(W3884), .A2(W27277), .ZN(W29376));
  NOR2X1 G1059 (.A1(I429), .A2(W21034), .ZN(O4867));
  NOR2X1 G1060 (.A1(W10270), .A2(W3671), .ZN(W11898));
  NOR2X1 G1061 (.A1(W33151), .A2(W753), .ZN(W38987));
  NOR2X1 G1062 (.A1(W36319), .A2(W9175), .ZN(O9907));
  NOR2X1 G1063 (.A1(W5178), .A2(W10045), .ZN(W11895));
  NOR2X1 G1064 (.A1(W9447), .A2(W10285), .ZN(W11894));
  NOR2X1 G1065 (.A1(W30738), .A2(W12284), .ZN(W38989));
  NOR2X1 G1066 (.A1(W35376), .A2(W8598), .ZN(O9908));
  NOR2X1 G1067 (.A1(W833), .A2(W3556), .ZN(W11891));
  NOR2X1 G1068 (.A1(I1098), .A2(W4480), .ZN(O549));
  NOR2X1 G1069 (.A1(W4625), .A2(W2203), .ZN(W11927));
  NOR2X1 G1070 (.A1(W25986), .A2(W22057), .ZN(W29387));
  NOR2X1 G1071 (.A1(W6384), .A2(W27901), .ZN(W29385));
  NOR2X1 G1072 (.A1(W324), .A2(W558), .ZN(W11924));
  NOR2X1 G1073 (.A1(W18426), .A2(W2653), .ZN(O2234));
  NOR2X1 G1074 (.A1(W6520), .A2(W3123), .ZN(W29384));
  NOR2X1 G1075 (.A1(W11570), .A2(W773), .ZN(W11921));
  NOR2X1 G1076 (.A1(W13270), .A2(W30499), .ZN(W38956));
  NOR2X1 G1077 (.A1(W2445), .A2(W9012), .ZN(O9910));
  NOR2X1 G1078 (.A1(I1811), .A2(W36130), .ZN(W38961));
  NOR2X1 G1079 (.A1(W143), .A2(W8027), .ZN(W21396));
  NOR2X1 G1080 (.A1(W20099), .A2(W10939), .ZN(W38965));
  NOR2X1 G1081 (.A1(W22325), .A2(W30076), .ZN(O9893));
  NOR2X1 G1082 (.A1(W28799), .A2(W19860), .ZN(O9895));
  NOR2X1 G1083 (.A1(W9921), .A2(W6890), .ZN(W11913));
  NOR2X1 G1084 (.A1(W8856), .A2(I1220), .ZN(O548));
  NOR2X1 G1085 (.A1(W1538), .A2(W5994), .ZN(W11862));
  NOR2X1 G1086 (.A1(W6070), .A2(W7238), .ZN(W11871));
  NOR2X1 G1087 (.A1(W4470), .A2(I429), .ZN(W11870));
  NOR2X1 G1088 (.A1(W26979), .A2(W28251), .ZN(O9916));
  NOR2X1 G1089 (.A1(W7355), .A2(W12813), .ZN(O9917));
  NOR2X1 G1090 (.A1(I1802), .A2(W4237), .ZN(W11867));
  NOR2X1 G1091 (.A1(W2880), .A2(W13919), .ZN(W21405));
  NOR2X1 G1092 (.A1(W11644), .A2(W2077), .ZN(W11864));
  NOR2X1 G1093 (.A1(W1379), .A2(W2701), .ZN(W11863));
  NOR2X1 G1094 (.A1(W23373), .A2(W38842), .ZN(O9914));
  NOR2X1 G1095 (.A1(W2982), .A2(W20975), .ZN(W29370));
  NOR2X1 G1096 (.A1(W37638), .A2(W35881), .ZN(W39012));
  NOR2X1 G1097 (.A1(W22979), .A2(W22398), .ZN(O4860));
  NOR2X1 G1098 (.A1(W10849), .A2(W9799), .ZN(W11857));
  NOR2X1 G1099 (.A1(W10902), .A2(W23843), .ZN(O9922));
  NOR2X1 G1100 (.A1(W4854), .A2(W31515), .ZN(O9924));
  NOR2X1 G1101 (.A1(W17579), .A2(W804), .ZN(O9925));
  NOR2X1 G1102 (.A1(W3026), .A2(W4899), .ZN(O544));
  NOR2X1 G1103 (.A1(W4706), .A2(W11139), .ZN(W11888));
  NOR2X1 G1104 (.A1(I953), .A2(W11776), .ZN(W11887));
  NOR2X1 G1105 (.A1(W16823), .A2(W6725), .ZN(O4864));
  NOR2X1 G1106 (.A1(I179), .A2(W34597), .ZN(O9912));
  NOR2X1 G1107 (.A1(W10669), .A2(W1992), .ZN(W11884));
  NOR2X1 G1108 (.A1(W10018), .A2(W30854), .ZN(W38999));
  NOR2X1 G1109 (.A1(W7932), .A2(I1993), .ZN(W11882));
  NOR2X1 G1110 (.A1(W15693), .A2(W10598), .ZN(W39000));
  NOR2X1 G1111 (.A1(W28919), .A2(W26923), .ZN(O9378));
  NOR2X1 G1112 (.A1(W11171), .A2(W7944), .ZN(W11879));
  NOR2X1 G1113 (.A1(I49), .A2(W11768), .ZN(W11878));
  NOR2X1 G1114 (.A1(W26551), .A2(W16759), .ZN(O9913));
  NOR2X1 G1115 (.A1(W2011), .A2(W11529), .ZN(W11876));
  NOR2X1 G1116 (.A1(I1956), .A2(W3420), .ZN(W39002));
  NOR2X1 G1117 (.A1(W5509), .A2(W3066), .ZN(W11874));
  NOR2X1 G1118 (.A1(W9120), .A2(W1802), .ZN(W11873));
  NOR2X1 G1119 (.A1(W16620), .A2(I815), .ZN(W20849));
  NOR2X1 G1120 (.A1(W29780), .A2(W34014), .ZN(W37278));
  NOR2X1 G1121 (.A1(W4875), .A2(W11471), .ZN(W13552));
  NOR2X1 G1122 (.A1(I948), .A2(W6238), .ZN(O755));
  NOR2X1 G1123 (.A1(W4355), .A2(W6555), .ZN(W13550));
  NOR2X1 G1124 (.A1(W4316), .A2(W35423), .ZN(W37279));
  NOR2X1 G1125 (.A1(W5188), .A2(I334), .ZN(W20848));
  NOR2X1 G1126 (.A1(W414), .A2(W7230), .ZN(W13547));
  NOR2X1 G1127 (.A1(W3736), .A2(W13360), .ZN(W13546));
  NOR2X1 G1128 (.A1(W5882), .A2(W3104), .ZN(O757));
  NOR2X1 G1129 (.A1(W19499), .A2(W32824), .ZN(O8886));
  NOR2X1 G1130 (.A1(W20358), .A2(W24704), .ZN(O8887));
  NOR2X1 G1131 (.A1(W18118), .A2(W35035), .ZN(W37287));
  NOR2X1 G1132 (.A1(W4607), .A2(W12342), .ZN(W20851));
  NOR2X1 G1133 (.A1(W25016), .A2(W8771), .ZN(W37293));
  NOR2X1 G1134 (.A1(W3959), .A2(W11394), .ZN(O754));
  NOR2X1 G1135 (.A1(W428), .A2(W8181), .ZN(W13537));
  NOR2X1 G1136 (.A1(W4205), .A2(W1866), .ZN(W37294));
  NOR2X1 G1137 (.A1(W7786), .A2(W31324), .ZN(O8878));
  NOR2X1 G1138 (.A1(W9618), .A2(W9908), .ZN(W13572));
  NOR2X1 G1139 (.A1(W2286), .A2(W5199), .ZN(W13570));
  NOR2X1 G1140 (.A1(I1072), .A2(W7893), .ZN(W13569));
  NOR2X1 G1141 (.A1(W7746), .A2(W7737), .ZN(W13568));
  NOR2X1 G1142 (.A1(W2046), .A2(W6552), .ZN(W13567));
  NOR2X1 G1143 (.A1(W10393), .A2(W24440), .ZN(O8876));
  NOR2X1 G1144 (.A1(W10192), .A2(W7947), .ZN(O759));
  NOR2X1 G1145 (.A1(I168), .A2(W4393), .ZN(W13564));
  NOR2X1 G1146 (.A1(W8396), .A2(W25270), .ZN(O5110));
  NOR2X1 G1147 (.A1(W11431), .A2(I314), .ZN(W13562));
  NOR2X1 G1148 (.A1(W31349), .A2(W12070), .ZN(O8879));
  NOR2X1 G1149 (.A1(W25776), .A2(W10955), .ZN(O8881));
  NOR2X1 G1150 (.A1(W2305), .A2(W9386), .ZN(W13559));
  NOR2X1 G1151 (.A1(W5805), .A2(W10842), .ZN(W13558));
  NOR2X1 G1152 (.A1(W9854), .A2(W7438), .ZN(W37274));
  NOR2X1 G1153 (.A1(W3942), .A2(W11283), .ZN(W13556));
  NOR2X1 G1154 (.A1(W8557), .A2(W7555), .ZN(W13507));
  NOR2X1 G1155 (.A1(W27681), .A2(W18923), .ZN(O8913));
  NOR2X1 G1156 (.A1(I989), .A2(W2333), .ZN(W13515));
  NOR2X1 G1157 (.A1(W9978), .A2(W9142), .ZN(W13514));
  NOR2X1 G1158 (.A1(W7005), .A2(W19052), .ZN(W20857));
  NOR2X1 G1159 (.A1(W1687), .A2(W9742), .ZN(W13512));
  NOR2X1 G1160 (.A1(W395), .A2(W10001), .ZN(W13511));
  NOR2X1 G1161 (.A1(W2950), .A2(W12998), .ZN(W13510));
  NOR2X1 G1162 (.A1(W25809), .A2(W20190), .ZN(O8914));
  NOR2X1 G1163 (.A1(W15898), .A2(W1048), .ZN(O8910));
  NOR2X1 G1164 (.A1(W11829), .A2(W11606), .ZN(O5106));
  NOR2X1 G1165 (.A1(W2600), .A2(W15026), .ZN(W20860));
  NOR2X1 G1166 (.A1(W12506), .A2(W20486), .ZN(W29908));
  NOR2X1 G1167 (.A1(W26238), .A2(W10531), .ZN(O8920));
  NOR2X1 G1168 (.A1(W9012), .A2(W2359), .ZN(W13501));
  NOR2X1 G1169 (.A1(W27892), .A2(W16876), .ZN(O8922));
  NOR2X1 G1170 (.A1(W6087), .A2(W8593), .ZN(W37338));
  NOR2X1 G1171 (.A1(W31417), .A2(W1088), .ZN(O8923));
  NOR2X1 G1172 (.A1(W32217), .A2(W11564), .ZN(W37307));
  NOR2X1 G1173 (.A1(W18078), .A2(W28769), .ZN(O8898));
  NOR2X1 G1174 (.A1(W8341), .A2(W10019), .ZN(W13533));
  NOR2X1 G1175 (.A1(W2566), .A2(W19854), .ZN(O8900));
  NOR2X1 G1176 (.A1(W646), .A2(W11513), .ZN(W37301));
  NOR2X1 G1177 (.A1(W1792), .A2(W9417), .ZN(O8902));
  NOR2X1 G1178 (.A1(W30581), .A2(W15866), .ZN(W37304));
  NOR2X1 G1179 (.A1(W3091), .A2(W25022), .ZN(O8903));
  NOR2X1 G1180 (.A1(W3991), .A2(W23001), .ZN(O5108));
  NOR2X1 G1181 (.A1(W4577), .A2(W11477), .ZN(W13573));
  NOR2X1 G1182 (.A1(I136), .A2(W27905), .ZN(W37308));
  NOR2X1 G1183 (.A1(W20478), .A2(W17188), .ZN(W37309));
  NOR2X1 G1184 (.A1(W12660), .A2(W1545), .ZN(O8906));
  NOR2X1 G1185 (.A1(W14926), .A2(W17703), .ZN(W20855));
  NOR2X1 G1186 (.A1(W2841), .A2(I923), .ZN(O8907));
  NOR2X1 G1187 (.A1(W9185), .A2(W8894), .ZN(W13519));
  NOR2X1 G1188 (.A1(W13142), .A2(W6681), .ZN(W29913));
  NOR2X1 G1189 (.A1(W17048), .A2(W1876), .ZN(W37215));
  NOR2X1 G1190 (.A1(W19458), .A2(W15908), .ZN(O8844));
  NOR2X1 G1191 (.A1(I871), .A2(W13884), .ZN(O8846));
  NOR2X1 G1192 (.A1(I14), .A2(W9369), .ZN(W13627));
  NOR2X1 G1193 (.A1(W2260), .A2(W13182), .ZN(W13626));
  NOR2X1 G1194 (.A1(W11658), .A2(W3916), .ZN(W13625));
  NOR2X1 G1195 (.A1(I1000), .A2(W9460), .ZN(W13624));
  NOR2X1 G1196 (.A1(W36880), .A2(W16317), .ZN(W37214));
  NOR2X1 G1197 (.A1(W5413), .A2(W7811), .ZN(W13622));
  NOR2X1 G1198 (.A1(W1917), .A2(W30631), .ZN(W37208));
  NOR2X1 G1199 (.A1(W1457), .A2(W8970), .ZN(W13620));
  NOR2X1 G1200 (.A1(W766), .A2(W2407), .ZN(W20831));
  NOR2X1 G1201 (.A1(W2872), .A2(W2860), .ZN(W29938));
  NOR2X1 G1202 (.A1(W12483), .A2(W20215), .ZN(O5117));
  NOR2X1 G1203 (.A1(W10862), .A2(W6389), .ZN(W13616));
  NOR2X1 G1204 (.A1(W18555), .A2(W25771), .ZN(W29936));
  NOR2X1 G1205 (.A1(W22825), .A2(W4541), .ZN(O8850));
  NOR2X1 G1206 (.A1(W7585), .A2(W20873), .ZN(W37224));
  NOR2X1 G1207 (.A1(W21373), .A2(W2979), .ZN(O8833));
  NOR2X1 G1208 (.A1(W6634), .A2(W4852), .ZN(W13648));
  NOR2X1 G1209 (.A1(W15994), .A2(W1040), .ZN(O2093));
  NOR2X1 G1210 (.A1(W8716), .A2(W12679), .ZN(W13646));
  NOR2X1 G1211 (.A1(W586), .A2(I952), .ZN(W13645));
  NOR2X1 G1212 (.A1(W31568), .A2(W26435), .ZN(W37186));
  NOR2X1 G1213 (.A1(W16537), .A2(W35228), .ZN(O8832));
  NOR2X1 G1214 (.A1(I29), .A2(W27039), .ZN(O5119));
  NOR2X1 G1215 (.A1(W4795), .A2(W18762), .ZN(W37191));
  NOR2X1 G1216 (.A1(W3033), .A2(W36386), .ZN(O8851));
  NOR2X1 G1217 (.A1(W4140), .A2(W1013), .ZN(W13639));
  NOR2X1 G1218 (.A1(W10208), .A2(I238), .ZN(W20825));
  NOR2X1 G1219 (.A1(W11973), .A2(W7178), .ZN(W20826));
  NOR2X1 G1220 (.A1(W5796), .A2(W31686), .ZN(W37198));
  NOR2X1 G1221 (.A1(W14421), .A2(I1442), .ZN(O2094));
  NOR2X1 G1222 (.A1(W23994), .A2(W3361), .ZN(W29941));
  NOR2X1 G1223 (.A1(W15639), .A2(W14202), .ZN(O8843));
  NOR2X1 G1224 (.A1(W26305), .A2(W22640), .ZN(W37255));
  NOR2X1 G1225 (.A1(W3033), .A2(W2169), .ZN(W13593));
  NOR2X1 G1226 (.A1(W8922), .A2(W7999), .ZN(O763));
  NOR2X1 G1227 (.A1(W9743), .A2(W7619), .ZN(W13591));
  NOR2X1 G1228 (.A1(W17576), .A2(W29368), .ZN(O8870));
  NOR2X1 G1229 (.A1(W33405), .A2(W4185), .ZN(W37249));
  NOR2X1 G1230 (.A1(W25025), .A2(W2531), .ZN(O8871));
  NOR2X1 G1231 (.A1(W20656), .A2(W2046), .ZN(W37252));
  NOR2X1 G1232 (.A1(W20497), .A2(W7610), .ZN(O5113));
  NOR2X1 G1233 (.A1(W6791), .A2(W9388), .ZN(W37245));
  NOR2X1 G1234 (.A1(W13921), .A2(W9677), .ZN(W20841));
  NOR2X1 G1235 (.A1(W2656), .A2(I1454), .ZN(W13581));
  NOR2X1 G1236 (.A1(W9100), .A2(W8448), .ZN(O2097));
  NOR2X1 G1237 (.A1(W13526), .A2(W17773), .ZN(W37258));
  NOR2X1 G1238 (.A1(W33835), .A2(I1377), .ZN(W37259));
  NOR2X1 G1239 (.A1(W18864), .A2(W29096), .ZN(W29929));
  NOR2X1 G1240 (.A1(W10911), .A2(W27189), .ZN(W37261));
  NOR2X1 G1241 (.A1(W21123), .A2(W5424), .ZN(W29928));
  NOR2X1 G1242 (.A1(I1182), .A2(W10277), .ZN(O765));
  NOR2X1 G1243 (.A1(W948), .A2(W1284), .ZN(W13611));
  NOR2X1 G1244 (.A1(W760), .A2(W17096), .ZN(O5116));
  NOR2X1 G1245 (.A1(W1359), .A2(W5918), .ZN(W13609));
  NOR2X1 G1246 (.A1(W4987), .A2(W249), .ZN(W13608));
  NOR2X1 G1247 (.A1(W8600), .A2(W10616), .ZN(W13607));
  NOR2X1 G1248 (.A1(W4119), .A2(W32642), .ZN(O8857));
  NOR2X1 G1249 (.A1(W4051), .A2(W11193), .ZN(W13605));
  NOR2X1 G1250 (.A1(W13063), .A2(W34789), .ZN(W37233));
  NOR2X1 G1251 (.A1(W6793), .A2(W2909), .ZN(W13496));
  NOR2X1 G1252 (.A1(W24407), .A2(W25836), .ZN(O8859));
  NOR2X1 G1253 (.A1(W3752), .A2(W12849), .ZN(O8861));
  NOR2X1 G1254 (.A1(W7909), .A2(W2001), .ZN(O8862));
  NOR2X1 G1255 (.A1(W28071), .A2(W19338), .ZN(O8864));
  NOR2X1 G1256 (.A1(W19769), .A2(W61), .ZN(O5115));
  NOR2X1 G1257 (.A1(W21719), .A2(W35968), .ZN(O8866));
  NOR2X1 G1258 (.A1(W10180), .A2(W4267), .ZN(O8868));
  NOR2X1 G1259 (.A1(W11163), .A2(W18384), .ZN(W29870));
  NOR2X1 G1260 (.A1(W7835), .A2(W1356), .ZN(W13396));
  NOR2X1 G1261 (.A1(W26060), .A2(W34678), .ZN(W37445));
  NOR2X1 G1262 (.A1(W29024), .A2(W1638), .ZN(O8985));
  NOR2X1 G1263 (.A1(W6367), .A2(W5945), .ZN(W20890));
  NOR2X1 G1264 (.A1(W3311), .A2(W15595), .ZN(W20891));
  NOR2X1 G1265 (.A1(W4014), .A2(W4998), .ZN(W29871));
  NOR2X1 G1266 (.A1(W4231), .A2(W9328), .ZN(W13389));
  NOR2X1 G1267 (.A1(W26658), .A2(W21292), .ZN(O8990));
  NOR2X1 G1268 (.A1(W5132), .A2(W25611), .ZN(O8982));
  NOR2X1 G1269 (.A1(W14840), .A2(W7555), .ZN(W37456));
  NOR2X1 G1270 (.A1(W222), .A2(I1450), .ZN(W13385));
  NOR2X1 G1271 (.A1(W18098), .A2(W23517), .ZN(W37457));
  NOR2X1 G1272 (.A1(W19840), .A2(W8399), .ZN(O5088));
  NOR2X1 G1273 (.A1(W4197), .A2(W30020), .ZN(O8993));
  NOR2X1 G1274 (.A1(W19533), .A2(W5348), .ZN(W37462));
  NOR2X1 G1275 (.A1(W12851), .A2(W6198), .ZN(W13380));
  NOR2X1 G1276 (.A1(W8638), .A2(W3667), .ZN(O5087));
  NOR2X1 G1277 (.A1(W5397), .A2(W7008), .ZN(W13407));
  NOR2X1 G1278 (.A1(I1532), .A2(W2235), .ZN(W13416));
  NOR2X1 G1279 (.A1(W10670), .A2(W11726), .ZN(W37426));
  NOR2X1 G1280 (.A1(I830), .A2(W12210), .ZN(W13414));
  NOR2X1 G1281 (.A1(W16458), .A2(W11043), .ZN(O8975));
  NOR2X1 G1282 (.A1(W7452), .A2(W1556), .ZN(W13411));
  NOR2X1 G1283 (.A1(W3212), .A2(W18640), .ZN(O2105));
  NOR2X1 G1284 (.A1(W23336), .A2(W32452), .ZN(W37432));
  NOR2X1 G1285 (.A1(W12295), .A2(W15212), .ZN(W37435));
  NOR2X1 G1286 (.A1(W6201), .A2(I1087), .ZN(W13378));
  NOR2X1 G1287 (.A1(W6140), .A2(W6434), .ZN(W13406));
  NOR2X1 G1288 (.A1(W28507), .A2(W21212), .ZN(O8980));
  NOR2X1 G1289 (.A1(I1984), .A2(W2064), .ZN(W13404));
  NOR2X1 G1290 (.A1(W23283), .A2(W18213), .ZN(W29876));
  NOR2X1 G1291 (.A1(W14194), .A2(W34079), .ZN(W37441));
  NOR2X1 G1292 (.A1(W12105), .A2(I1917), .ZN(W13401));
  NOR2X1 G1293 (.A1(W4190), .A2(W7433), .ZN(W13400));
  NOR2X1 G1294 (.A1(W6478), .A2(W1069), .ZN(O9013));
  NOR2X1 G1295 (.A1(W8110), .A2(W9207), .ZN(W13356));
  NOR2X1 G1296 (.A1(W11540), .A2(W25278), .ZN(W29859));
  NOR2X1 G1297 (.A1(W4135), .A2(W9368), .ZN(W29858));
  NOR2X1 G1298 (.A1(W12646), .A2(W9737), .ZN(W13353));
  NOR2X1 G1299 (.A1(W12848), .A2(I704), .ZN(W13352));
  NOR2X1 G1300 (.A1(W2005), .A2(W945), .ZN(W20906));
  NOR2X1 G1301 (.A1(W7344), .A2(W12323), .ZN(O2107));
  NOR2X1 G1302 (.A1(W627), .A2(W12029), .ZN(W20908));
  NOR2X1 G1303 (.A1(I1126), .A2(W4777), .ZN(O5082));
  NOR2X1 G1304 (.A1(W678), .A2(W2869), .ZN(W13347));
  NOR2X1 G1305 (.A1(W13099), .A2(W1778), .ZN(O9016));
  NOR2X1 G1306 (.A1(W840), .A2(W11885), .ZN(W13343));
  NOR2X1 G1307 (.A1(W3419), .A2(I32), .ZN(O732));
  NOR2X1 G1308 (.A1(W1490), .A2(W10224), .ZN(O5080));
  NOR2X1 G1309 (.A1(W3467), .A2(W28225), .ZN(O9018));
  NOR2X1 G1310 (.A1(W22157), .A2(W13428), .ZN(O5078));
  NOR2X1 G1311 (.A1(W17394), .A2(W23217), .ZN(W29847));
  NOR2X1 G1312 (.A1(W8983), .A2(W4297), .ZN(W13366));
  NOR2X1 G1313 (.A1(W22647), .A2(W11393), .ZN(W29867));
  NOR2X1 G1314 (.A1(W104), .A2(W12364), .ZN(O736));
  NOR2X1 G1315 (.A1(W24510), .A2(W26592), .ZN(O8996));
  NOR2X1 G1316 (.A1(W12946), .A2(W3507), .ZN(W13373));
  NOR2X1 G1317 (.A1(W11287), .A2(W5624), .ZN(W13372));
  NOR2X1 G1318 (.A1(W2659), .A2(W7978), .ZN(W13370));
  NOR2X1 G1319 (.A1(W5429), .A2(W9364), .ZN(O8998));
  NOR2X1 G1320 (.A1(W5851), .A2(W28100), .ZN(W37472));
  NOR2X1 G1321 (.A1(W26965), .A2(W17137), .ZN(W29879));
  NOR2X1 G1322 (.A1(W22076), .A2(I1700), .ZN(O5084));
  NOR2X1 G1323 (.A1(W10914), .A2(I1991), .ZN(W13364));
  NOR2X1 G1324 (.A1(W6625), .A2(W5734), .ZN(W13363));
  NOR2X1 G1325 (.A1(W1136), .A2(W22561), .ZN(O9000));
  NOR2X1 G1326 (.A1(W5814), .A2(W4943), .ZN(O9001));
  NOR2X1 G1327 (.A1(I1612), .A2(W5490), .ZN(W13360));
  NOR2X1 G1328 (.A1(W21449), .A2(W1226), .ZN(W37479));
  NOR2X1 G1329 (.A1(W34502), .A2(W3198), .ZN(O8947));
  NOR2X1 G1330 (.A1(W703), .A2(W30305), .ZN(W37368));
  NOR2X1 G1331 (.A1(W4023), .A2(W25202), .ZN(O8943));
  NOR2X1 G1332 (.A1(W7127), .A2(W819), .ZN(W13472));
  NOR2X1 G1333 (.A1(W7846), .A2(W4582), .ZN(W29894));
  NOR2X1 G1334 (.A1(W1371), .A2(W33101), .ZN(W37372));
  NOR2X1 G1335 (.A1(W1360), .A2(I671), .ZN(W13468));
  NOR2X1 G1336 (.A1(W28545), .A2(W28865), .ZN(W29892));
  NOR2X1 G1337 (.A1(W30631), .A2(W12004), .ZN(O8946));
  NOR2X1 G1338 (.A1(W12090), .A2(W16431), .ZN(W37367));
  NOR2X1 G1339 (.A1(W25305), .A2(W13074), .ZN(O8948));
  NOR2X1 G1340 (.A1(W17121), .A2(W28540), .ZN(O8950));
  NOR2X1 G1341 (.A1(W4624), .A2(W4789), .ZN(W13462));
  NOR2X1 G1342 (.A1(I501), .A2(W6790), .ZN(W13461));
  NOR2X1 G1343 (.A1(W24232), .A2(W8295), .ZN(W37383));
  NOR2X1 G1344 (.A1(W32674), .A2(W20969), .ZN(O8952));
  NOR2X1 G1345 (.A1(W13509), .A2(W2947), .ZN(O8953));
  NOR2X1 G1346 (.A1(W12498), .A2(W7606), .ZN(W13456));
  NOR2X1 G1347 (.A1(W14233), .A2(W10341), .ZN(W37351));
  NOR2X1 G1348 (.A1(W10601), .A2(W9095), .ZN(W13495));
  NOR2X1 G1349 (.A1(I1252), .A2(W16825), .ZN(O8926));
  NOR2X1 G1350 (.A1(W10534), .A2(W1293), .ZN(W13493));
  NOR2X1 G1351 (.A1(W63), .A2(W18564), .ZN(O8927));
  NOR2X1 G1352 (.A1(W354), .A2(I1675), .ZN(W13491));
  NOR2X1 G1353 (.A1(I1820), .A2(W12531), .ZN(W13490));
  NOR2X1 G1354 (.A1(W17727), .A2(W3249), .ZN(O8931));
  NOR2X1 G1355 (.A1(W9601), .A2(W8061), .ZN(W13486));
  NOR2X1 G1356 (.A1(W27655), .A2(W15136), .ZN(W37387));
  NOR2X1 G1357 (.A1(W33413), .A2(W33652), .ZN(O8933));
  NOR2X1 G1358 (.A1(W16597), .A2(W4941), .ZN(O2102));
  NOR2X1 G1359 (.A1(W11922), .A2(W29640), .ZN(W37354));
  NOR2X1 G1360 (.A1(W11730), .A2(W3929), .ZN(W13481));
  NOR2X1 G1361 (.A1(W7379), .A2(W21640), .ZN(W29896));
  NOR2X1 G1362 (.A1(W30294), .A2(W4958), .ZN(O8941));
  NOR2X1 G1363 (.A1(W25575), .A2(W22928), .ZN(O8942));
  NOR2X1 G1364 (.A1(W726), .A2(W34811), .ZN(W37418));
  NOR2X1 G1365 (.A1(W7559), .A2(W12501), .ZN(O5093));
  NOR2X1 G1366 (.A1(W10093), .A2(W3782), .ZN(O741));
  NOR2X1 G1367 (.A1(I890), .A2(W10353), .ZN(O8965));
  NOR2X1 G1368 (.A1(W13386), .A2(W1761), .ZN(W13432));
  NOR2X1 G1369 (.A1(I512), .A2(W6698), .ZN(O8967));
  NOR2X1 G1370 (.A1(W33344), .A2(W25795), .ZN(W37414));
  NOR2X1 G1371 (.A1(W3821), .A2(W8050), .ZN(W13429));
  NOR2X1 G1372 (.A1(W16873), .A2(W35503), .ZN(O8970));
  NOR2X1 G1373 (.A1(W16929), .A2(W6005), .ZN(W20880));
  NOR2X1 G1374 (.A1(W2401), .A2(I186), .ZN(W13426));
  NOR2X1 G1375 (.A1(W8916), .A2(W10153), .ZN(W29881));
  NOR2X1 G1376 (.A1(I1150), .A2(W8400), .ZN(O740));
  NOR2X1 G1377 (.A1(W36881), .A2(W32036), .ZN(O8973));
  NOR2X1 G1378 (.A1(W29704), .A2(W4661), .ZN(W37423));
  NOR2X1 G1379 (.A1(W5595), .A2(W9404), .ZN(W13420));
  NOR2X1 G1380 (.A1(W3047), .A2(W13392), .ZN(W13419));
  NOR2X1 G1381 (.A1(W25635), .A2(W30618), .ZN(O8974));
  NOR2X1 G1382 (.A1(W5353), .A2(W10145), .ZN(W37396));
  NOR2X1 G1383 (.A1(W19033), .A2(W14730), .ZN(W20875));
  NOR2X1 G1384 (.A1(W31067), .A2(W15684), .ZN(O8956));
  NOR2X1 G1385 (.A1(W20868), .A2(W2272), .ZN(O8957));
  NOR2X1 G1386 (.A1(W4981), .A2(W3916), .ZN(W13450));
  NOR2X1 G1387 (.A1(W641), .A2(W8458), .ZN(W13449));
  NOR2X1 G1388 (.A1(W802), .A2(I1813), .ZN(W13448));
  NOR2X1 G1389 (.A1(W11860), .A2(W2877), .ZN(O5097));
  NOR2X1 G1390 (.A1(W20393), .A2(W11338), .ZN(O2104));
  NOR2X1 G1391 (.A1(W11155), .A2(W5316), .ZN(W13649));
  NOR2X1 G1392 (.A1(W22107), .A2(I328), .ZN(O8961));
  NOR2X1 G1393 (.A1(W24552), .A2(W24813), .ZN(O5094));
  NOR2X1 G1394 (.A1(W31863), .A2(W30790), .ZN(W37401));
  NOR2X1 G1395 (.A1(W25819), .A2(W21540), .ZN(O8963));
  NOR2X1 G1396 (.A1(W1269), .A2(W147), .ZN(W13439));
  NOR2X1 G1397 (.A1(W8311), .A2(W794), .ZN(W13438));
  NOR2X1 G1398 (.A1(W8694), .A2(I1738), .ZN(W13437));
  NOR2X1 G1399 (.A1(W25092), .A2(W30653), .ZN(W36972));
  NOR2X1 G1400 (.A1(W12320), .A2(W4298), .ZN(W13868));
  NOR2X1 G1401 (.A1(W2556), .A2(W7075), .ZN(W13867));
  NOR2X1 G1402 (.A1(W22823), .A2(W24542), .ZN(W30024));
  NOR2X1 G1403 (.A1(W6317), .A2(W12506), .ZN(O8707));
  NOR2X1 G1404 (.A1(I1594), .A2(W10054), .ZN(W13864));
  NOR2X1 G1405 (.A1(W9262), .A2(I1034), .ZN(O5158));
  NOR2X1 G1406 (.A1(W25830), .A2(W3679), .ZN(O8709));
  NOR2X1 G1407 (.A1(W9972), .A2(W2034), .ZN(W13861));
  NOR2X1 G1408 (.A1(W4156), .A2(W11767), .ZN(W20746));
  NOR2X1 G1409 (.A1(W3452), .A2(W54), .ZN(O793));
  NOR2X1 G1410 (.A1(W17331), .A2(W3607), .ZN(O8710));
  NOR2X1 G1411 (.A1(W33383), .A2(W27139), .ZN(W36974));
  NOR2X1 G1412 (.A1(W5989), .A2(W2398), .ZN(W13856));
  NOR2X1 G1413 (.A1(W12858), .A2(W14987), .ZN(O5157));
  NOR2X1 G1414 (.A1(W27253), .A2(W7928), .ZN(W36977));
  NOR2X1 G1415 (.A1(W33463), .A2(W22603), .ZN(O8713));
  NOR2X1 G1416 (.A1(W32236), .A2(W18462), .ZN(O8714));
  NOR2X1 G1417 (.A1(W33787), .A2(W7699), .ZN(O8697));
  NOR2X1 G1418 (.A1(W8582), .A2(W15427), .ZN(W30025));
  NOR2X1 G1419 (.A1(W9308), .A2(I1674), .ZN(W13884));
  NOR2X1 G1420 (.A1(W28852), .A2(I481), .ZN(W36938));
  NOR2X1 G1421 (.A1(W3462), .A2(W12582), .ZN(W13882));
  NOR2X1 G1422 (.A1(W18187), .A2(W19633), .ZN(W20743));
  NOR2X1 G1423 (.A1(W17234), .A2(W4551), .ZN(O8689));
  NOR2X1 G1424 (.A1(I8), .A2(W207), .ZN(W13879));
  NOR2X1 G1425 (.A1(W1158), .A2(W31216), .ZN(O8692));
  NOR2X1 G1426 (.A1(W497), .A2(W5780), .ZN(W13851));
  NOR2X1 G1427 (.A1(W25175), .A2(W17892), .ZN(W36955));
  NOR2X1 G1428 (.A1(I1982), .A2(W3282), .ZN(W20744));
  NOR2X1 G1429 (.A1(W4687), .A2(W10147), .ZN(W13874));
  NOR2X1 G1430 (.A1(W10297), .A2(W16615), .ZN(O8699));
  NOR2X1 G1431 (.A1(W11286), .A2(W1162), .ZN(W20745));
  NOR2X1 G1432 (.A1(W6342), .A2(W13832), .ZN(O8702));
  NOR2X1 G1433 (.A1(W2896), .A2(W31345), .ZN(O8704));
  NOR2X1 G1434 (.A1(W19143), .A2(W15135), .ZN(W20761));
  NOR2X1 G1435 (.A1(W8853), .A2(I525), .ZN(W13826));
  NOR2X1 G1436 (.A1(W32903), .A2(W2413), .ZN(O8726));
  NOR2X1 G1437 (.A1(W8658), .A2(W8789), .ZN(W13824));
  NOR2X1 G1438 (.A1(W9620), .A2(W5129), .ZN(W13823));
  NOR2X1 G1439 (.A1(W3763), .A2(W3178), .ZN(W20759));
  NOR2X1 G1440 (.A1(W8455), .A2(W5538), .ZN(O788));
  NOR2X1 G1441 (.A1(W4041), .A2(W7850), .ZN(W13819));
  NOR2X1 G1442 (.A1(W19907), .A2(W26406), .ZN(O8728));
  NOR2X1 G1443 (.A1(W25337), .A2(W35069), .ZN(W37006));
  NOR2X1 G1444 (.A1(W7770), .A2(W9618), .ZN(W13816));
  NOR2X1 G1445 (.A1(W8451), .A2(W27446), .ZN(W30005));
  NOR2X1 G1446 (.A1(I866), .A2(W12400), .ZN(W30003));
  NOR2X1 G1447 (.A1(W8599), .A2(W5754), .ZN(O787));
  NOR2X1 G1448 (.A1(W9182), .A2(W11521), .ZN(W13811));
  NOR2X1 G1449 (.A1(W16659), .A2(W7136), .ZN(O2075));
  NOR2X1 G1450 (.A1(I991), .A2(W18410), .ZN(W20766));
  NOR2X1 G1451 (.A1(W17519), .A2(W7646), .ZN(O2076));
  NOR2X1 G1452 (.A1(W20168), .A2(W2183), .ZN(W37001));
  NOR2X1 G1453 (.A1(W1197), .A2(I1657), .ZN(W13850));
  NOR2X1 G1454 (.A1(I1710), .A2(W30351), .ZN(O8715));
  NOR2X1 G1455 (.A1(W3571), .A2(W27398), .ZN(W30019));
  NOR2X1 G1456 (.A1(W727), .A2(I960), .ZN(W13845));
  NOR2X1 G1457 (.A1(W22271), .A2(W24218), .ZN(W36990));
  NOR2X1 G1458 (.A1(W12230), .A2(W2591), .ZN(W13842));
  NOR2X1 G1459 (.A1(W17242), .A2(W2157), .ZN(O8719));
  NOR2X1 G1460 (.A1(W892), .A2(W1188), .ZN(O8720));
  NOR2X1 G1461 (.A1(W28694), .A2(W8660), .ZN(W36936));
  NOR2X1 G1462 (.A1(W5847), .A2(W35640), .ZN(W37002));
  NOR2X1 G1463 (.A1(W16673), .A2(W24418), .ZN(O5152));
  NOR2X1 G1464 (.A1(W35694), .A2(W19244), .ZN(O8725));
  NOR2X1 G1465 (.A1(W11140), .A2(W1897), .ZN(W13831));
  NOR2X1 G1466 (.A1(W12783), .A2(W10283), .ZN(W13830));
  NOR2X1 G1467 (.A1(W2185), .A2(W4568), .ZN(W13829));
  NOR2X1 G1468 (.A1(W5748), .A2(W12468), .ZN(W13828));
  NOR2X1 G1469 (.A1(W10865), .A2(W19662), .ZN(O2069));
  NOR2X1 G1470 (.A1(W10503), .A2(W1267), .ZN(W13940));
  NOR2X1 G1471 (.A1(W13751), .A2(W3485), .ZN(W36880));
  NOR2X1 G1472 (.A1(W1853), .A2(W7657), .ZN(W13938));
  NOR2X1 G1473 (.A1(W8607), .A2(I868), .ZN(O807));
  NOR2X1 G1474 (.A1(W4644), .A2(W2798), .ZN(W13936));
  NOR2X1 G1475 (.A1(W36123), .A2(W7182), .ZN(W36881));
  NOR2X1 G1476 (.A1(W28232), .A2(W29503), .ZN(O8649));
  NOR2X1 G1477 (.A1(W18018), .A2(W33517), .ZN(O8650));
  NOR2X1 G1478 (.A1(W5576), .A2(W7066), .ZN(W13941));
  NOR2X1 G1479 (.A1(W5877), .A2(W4285), .ZN(W13931));
  NOR2X1 G1480 (.A1(W20710), .A2(W12444), .ZN(W30039));
  NOR2X1 G1481 (.A1(W7416), .A2(W21018), .ZN(O5165));
  NOR2X1 G1482 (.A1(W33542), .A2(W7443), .ZN(W36890));
  NOR2X1 G1483 (.A1(W10857), .A2(W4475), .ZN(O8655));
  NOR2X1 G1484 (.A1(W8589), .A2(W2718), .ZN(W13926));
  NOR2X1 G1485 (.A1(W13183), .A2(W13386), .ZN(W13925));
  NOR2X1 G1486 (.A1(W826), .A2(W7297), .ZN(W13924));
  NOR2X1 G1487 (.A1(W22177), .A2(W34712), .ZN(W36863));
  NOR2X1 G1488 (.A1(W15082), .A2(W33128), .ZN(O8635));
  NOR2X1 G1489 (.A1(W6649), .A2(W3408), .ZN(O8636));
  NOR2X1 G1490 (.A1(W7801), .A2(W6140), .ZN(O8637));
  NOR2X1 G1491 (.A1(W1645), .A2(W12264), .ZN(O2067));
  NOR2X1 G1492 (.A1(I1975), .A2(I1959), .ZN(W13954));
  NOR2X1 G1493 (.A1(W10718), .A2(W6075), .ZN(W13953));
  NOR2X1 G1494 (.A1(W5681), .A2(W4034), .ZN(O809));
  NOR2X1 G1495 (.A1(W19070), .A2(W1024), .ZN(W36862));
  NOR2X1 G1496 (.A1(W13367), .A2(W4421), .ZN(W36892));
  NOR2X1 G1497 (.A1(W10125), .A2(W835), .ZN(O8640));
  NOR2X1 G1498 (.A1(W19350), .A2(W19266), .ZN(O8643));
  NOR2X1 G1499 (.A1(W1311), .A2(W14450), .ZN(O8644));
  NOR2X1 G1500 (.A1(I120), .A2(W5899), .ZN(O808));
  NOR2X1 G1501 (.A1(W1322), .A2(W8641), .ZN(O2068));
  NOR2X1 G1502 (.A1(W23616), .A2(W36347), .ZN(O8646));
  NOR2X1 G1503 (.A1(W1816), .A2(W21065), .ZN(W30041));
  NOR2X1 G1504 (.A1(W3127), .A2(W6465), .ZN(W13896));
  NOR2X1 G1505 (.A1(W7393), .A2(W18292), .ZN(O8672));
  NOR2X1 G1506 (.A1(W19556), .A2(W10078), .ZN(W30030));
  NOR2X1 G1507 (.A1(W6954), .A2(W24114), .ZN(O8676));
  NOR2X1 G1508 (.A1(I659), .A2(W12770), .ZN(W13901));
  NOR2X1 G1509 (.A1(W9222), .A2(W8264), .ZN(W13900));
  NOR2X1 G1510 (.A1(W12292), .A2(W5875), .ZN(W13899));
  NOR2X1 G1511 (.A1(W6837), .A2(W1310), .ZN(O799));
  NOR2X1 G1512 (.A1(W20589), .A2(W30509), .ZN(W36926));
  NOR2X1 G1513 (.A1(W26298), .A2(W25167), .ZN(O8671));
  NOR2X1 G1514 (.A1(W12972), .A2(W10761), .ZN(W13895));
  NOR2X1 G1515 (.A1(W12161), .A2(W9127), .ZN(W13894));
  NOR2X1 G1516 (.A1(W1655), .A2(W4016), .ZN(W13893));
  NOR2X1 G1517 (.A1(W18731), .A2(W6952), .ZN(O8682));
  NOR2X1 G1518 (.A1(W7239), .A2(W9478), .ZN(W13891));
  NOR2X1 G1519 (.A1(W13303), .A2(W6899), .ZN(O798));
  NOR2X1 G1520 (.A1(W5169), .A2(W18842), .ZN(O5159));
  NOR2X1 G1521 (.A1(W16863), .A2(W1210), .ZN(O8686));
  NOR2X1 G1522 (.A1(I386), .A2(W32353), .ZN(O8665));
  NOR2X1 G1523 (.A1(W30522), .A2(W1437), .ZN(O8657));
  NOR2X1 G1524 (.A1(W16831), .A2(W27408), .ZN(O8658));
  NOR2X1 G1525 (.A1(W11239), .A2(W729), .ZN(W30035));
  NOR2X1 G1526 (.A1(I1079), .A2(W6380), .ZN(W13919));
  NOR2X1 G1527 (.A1(W26834), .A2(W1644), .ZN(W36897));
  NOR2X1 G1528 (.A1(W5039), .A2(I635), .ZN(W13917));
  NOR2X1 G1529 (.A1(W23055), .A2(W28749), .ZN(O8660));
  NOR2X1 G1530 (.A1(W20107), .A2(W1409), .ZN(O5163));
  NOR2X1 G1531 (.A1(W3385), .A2(W9855), .ZN(W13806));
  NOR2X1 G1532 (.A1(I1250), .A2(W3984), .ZN(W36908));
  NOR2X1 G1533 (.A1(W9645), .A2(W2341), .ZN(W20737));
  NOR2X1 G1534 (.A1(W231), .A2(W15734), .ZN(W36911));
  NOR2X1 G1535 (.A1(W24406), .A2(W25073), .ZN(W36912));
  NOR2X1 G1536 (.A1(I1862), .A2(W108), .ZN(W20738));
  NOR2X1 G1537 (.A1(W31604), .A2(W21300), .ZN(O8670));
  NOR2X1 G1538 (.A1(W10061), .A2(W13222), .ZN(W13906));
  NOR2X1 G1539 (.A1(W35893), .A2(W35098), .ZN(W37135));
  NOR2X1 G1540 (.A1(W3528), .A2(W4654), .ZN(W13708));
  NOR2X1 G1541 (.A1(W20002), .A2(W11493), .ZN(O8797));
  NOR2X1 G1542 (.A1(W14746), .A2(W9290), .ZN(W37130));
  NOR2X1 G1543 (.A1(W16962), .A2(W32775), .ZN(O8798));
  NOR2X1 G1544 (.A1(W6453), .A2(W1726), .ZN(W13704));
  NOR2X1 G1545 (.A1(W16569), .A2(I80), .ZN(W20803));
  NOR2X1 G1546 (.A1(I410), .A2(W8246), .ZN(W13702));
  NOR2X1 G1547 (.A1(W19217), .A2(W9167), .ZN(W37134));
  NOR2X1 G1548 (.A1(W16598), .A2(W30636), .ZN(W37126));
  NOR2X1 G1549 (.A1(W9171), .A2(W611), .ZN(W13699));
  NOR2X1 G1550 (.A1(W277), .A2(W11002), .ZN(W13698));
  NOR2X1 G1551 (.A1(W12537), .A2(W5208), .ZN(W20805));
  NOR2X1 G1552 (.A1(W1647), .A2(W24522), .ZN(W37139));
  NOR2X1 G1553 (.A1(I1079), .A2(W13108), .ZN(W13693));
  NOR2X1 G1554 (.A1(W1766), .A2(W8896), .ZN(W13692));
  NOR2X1 G1555 (.A1(W1877), .A2(W3401), .ZN(W13691));
  NOR2X1 G1556 (.A1(W15610), .A2(W29781), .ZN(W29955));
  NOR2X1 G1557 (.A1(I929), .A2(W7376), .ZN(W13717));
  NOR2X1 G1558 (.A1(W15143), .A2(W6911), .ZN(O5129));
  NOR2X1 G1559 (.A1(W5099), .A2(W10122), .ZN(W13726));
  NOR2X1 G1560 (.A1(W7315), .A2(W8149), .ZN(W13725));
  NOR2X1 G1561 (.A1(W20038), .A2(W27032), .ZN(W37115));
  NOR2X1 G1562 (.A1(W4214), .A2(W8374), .ZN(W13723));
  NOR2X1 G1563 (.A1(W34288), .A2(W3845), .ZN(O8788));
  NOR2X1 G1564 (.A1(W1564), .A2(W26132), .ZN(W29961));
  NOR2X1 G1565 (.A1(W11364), .A2(W11395), .ZN(W13718));
  NOR2X1 G1566 (.A1(W29576), .A2(W5689), .ZN(O8804));
  NOR2X1 G1567 (.A1(W12280), .A2(W6102), .ZN(W20801));
  NOR2X1 G1568 (.A1(W36578), .A2(I1112), .ZN(W37122));
  NOR2X1 G1569 (.A1(W11646), .A2(W9382), .ZN(W13714));
  NOR2X1 G1570 (.A1(W12914), .A2(W14565), .ZN(W20802));
  NOR2X1 G1571 (.A1(W9765), .A2(W36696), .ZN(W37124));
  NOR2X1 G1572 (.A1(W7894), .A2(W10435), .ZN(W13711));
  NOR2X1 G1573 (.A1(I206), .A2(W7407), .ZN(O8795));
  NOR2X1 G1574 (.A1(W23999), .A2(W10364), .ZN(W37175));
  NOR2X1 G1575 (.A1(W182), .A2(W7837), .ZN(W13669));
  NOR2X1 G1576 (.A1(W411), .A2(W13093), .ZN(O772));
  NOR2X1 G1577 (.A1(W10009), .A2(W20485), .ZN(O2089));
  NOR2X1 G1578 (.A1(W3306), .A2(W5436), .ZN(W13665));
  NOR2X1 G1579 (.A1(W6624), .A2(W6233), .ZN(W13664));
  NOR2X1 G1580 (.A1(W3775), .A2(W30947), .ZN(O8817));
  NOR2X1 G1581 (.A1(W31287), .A2(W20001), .ZN(O8819));
  NOR2X1 G1582 (.A1(W32125), .A2(W28275), .ZN(O8820));
  NOR2X1 G1583 (.A1(W3460), .A2(W13315), .ZN(O8815));
  NOR2X1 G1584 (.A1(W7533), .A2(W13978), .ZN(O2091));
  NOR2X1 G1585 (.A1(W7521), .A2(W2262), .ZN(W20818));
  NOR2X1 G1586 (.A1(W28906), .A2(W26197), .ZN(O8825));
  NOR2X1 G1587 (.A1(W11590), .A2(W2961), .ZN(W20820));
  NOR2X1 G1588 (.A1(W276), .A2(W8112), .ZN(W13653));
  NOR2X1 G1589 (.A1(W9201), .A2(W6833), .ZN(O769));
  NOR2X1 G1590 (.A1(W9211), .A2(W9994), .ZN(W20821));
  NOR2X1 G1591 (.A1(W7506), .A2(W5701), .ZN(O2092));
  NOR2X1 G1592 (.A1(I1868), .A2(I1706), .ZN(W37149));
  NOR2X1 G1593 (.A1(W32899), .A2(W27613), .ZN(O8805));
  NOR2X1 G1594 (.A1(W7576), .A2(W2277), .ZN(W13687));
  NOR2X1 G1595 (.A1(W35088), .A2(W8570), .ZN(W37144));
  NOR2X1 G1596 (.A1(W9102), .A2(W32955), .ZN(W37145));
  NOR2X1 G1597 (.A1(W2211), .A2(W29908), .ZN(W37147));
  NOR2X1 G1598 (.A1(W6548), .A2(W6727), .ZN(W13683));
  NOR2X1 G1599 (.A1(W15960), .A2(W15241), .ZN(W37148));
  NOR2X1 G1600 (.A1(W12436), .A2(W3332), .ZN(W13681));
  NOR2X1 G1601 (.A1(W14827), .A2(W24606), .ZN(W37111));
  NOR2X1 G1602 (.A1(W19789), .A2(W504), .ZN(W20808));
  NOR2X1 G1603 (.A1(W12749), .A2(W14604), .ZN(O2087));
  NOR2X1 G1604 (.A1(W2511), .A2(W4469), .ZN(W20812));
  NOR2X1 G1605 (.A1(W25142), .A2(W20821), .ZN(O8813));
  NOR2X1 G1606 (.A1(W12273), .A2(I1161), .ZN(W29952));
  NOR2X1 G1607 (.A1(W8775), .A2(W182), .ZN(W13672));
  NOR2X1 G1608 (.A1(W10608), .A2(W11738), .ZN(O773));
  NOR2X1 G1609 (.A1(W32373), .A2(W18556), .ZN(O8746));
  NOR2X1 G1610 (.A1(W4757), .A2(I252), .ZN(O784));
  NOR2X1 G1611 (.A1(W2008), .A2(W12443), .ZN(W13786));
  NOR2X1 G1612 (.A1(W35534), .A2(W28860), .ZN(W37043));
  NOR2X1 G1613 (.A1(W4766), .A2(W19706), .ZN(W20774));
  NOR2X1 G1614 (.A1(W13000), .A2(W8386), .ZN(W13782));
  NOR2X1 G1615 (.A1(W35135), .A2(W23106), .ZN(W37046));
  NOR2X1 G1616 (.A1(W12136), .A2(W28141), .ZN(W37049));
  NOR2X1 G1617 (.A1(I498), .A2(W1465), .ZN(W13779));
  NOR2X1 G1618 (.A1(W34267), .A2(W12191), .ZN(W37042));
  NOR2X1 G1619 (.A1(W8207), .A2(W6016), .ZN(W13776));
  NOR2X1 G1620 (.A1(W13691), .A2(W16837), .ZN(W29989));
  NOR2X1 G1621 (.A1(W1851), .A2(W8703), .ZN(W13772));
  NOR2X1 G1622 (.A1(W18905), .A2(W3724), .ZN(W20780));
  NOR2X1 G1623 (.A1(W31805), .A2(W2683), .ZN(W37059));
  NOR2X1 G1624 (.A1(W5148), .A2(W11063), .ZN(W13769));
  NOR2X1 G1625 (.A1(W4678), .A2(W26851), .ZN(O8753));
  NOR2X1 G1626 (.A1(W4154), .A2(W6869), .ZN(O783));
  NOR2X1 G1627 (.A1(W2177), .A2(W23357), .ZN(W29998));
  NOR2X1 G1628 (.A1(W6116), .A2(W10691), .ZN(W20769));
  NOR2X1 G1629 (.A1(W20183), .A2(W17511), .ZN(O8735));
  NOR2X1 G1630 (.A1(W503), .A2(I1446), .ZN(W13803));
  NOR2X1 G1631 (.A1(W21068), .A2(W14271), .ZN(O5148));
  NOR2X1 G1632 (.A1(W3576), .A2(W12621), .ZN(W13801));
  NOR2X1 G1633 (.A1(W10212), .A2(W3395), .ZN(W13800));
  NOR2X1 G1634 (.A1(I1881), .A2(W11664), .ZN(W13799));
  NOR2X1 G1635 (.A1(W22294), .A2(W34841), .ZN(W37035));
  NOR2X1 G1636 (.A1(W19778), .A2(W18394), .ZN(O2080));
  NOR2X1 G1637 (.A1(W6952), .A2(W13666), .ZN(W13795));
  NOR2X1 G1638 (.A1(W10410), .A2(W8524), .ZN(O785));
  NOR2X1 G1639 (.A1(W4147), .A2(W11253), .ZN(W13793));
  NOR2X1 G1640 (.A1(W10261), .A2(W5114), .ZN(W13792));
  NOR2X1 G1641 (.A1(W25536), .A2(W16459), .ZN(O5145));
  NOR2X1 G1642 (.A1(W12665), .A2(W30484), .ZN(W37041));
  NOR2X1 G1643 (.A1(W7203), .A2(W2189), .ZN(W13789));
  NOR2X1 G1644 (.A1(W546), .A2(W12992), .ZN(O5131));
  NOR2X1 G1645 (.A1(W3520), .A2(I1258), .ZN(W13746));
  NOR2X1 G1646 (.A1(W27149), .A2(W19956), .ZN(W29976));
  NOR2X1 G1647 (.A1(W8846), .A2(W3419), .ZN(W13742));
  NOR2X1 G1648 (.A1(W34948), .A2(W16923), .ZN(O8775));
  NOR2X1 G1649 (.A1(I660), .A2(W2376), .ZN(W13740));
  NOR2X1 G1650 (.A1(W17678), .A2(W18062), .ZN(O2085));
  NOR2X1 G1651 (.A1(W14631), .A2(W10961), .ZN(O8779));
  NOR2X1 G1652 (.A1(W6684), .A2(W3228), .ZN(O781));
  NOR2X1 G1653 (.A1(W4700), .A2(W11860), .ZN(W13747));
  NOR2X1 G1654 (.A1(W10229), .A2(W7411), .ZN(W13735));
  NOR2X1 G1655 (.A1(W19065), .A2(W2149), .ZN(W20794));
  NOR2X1 G1656 (.A1(W3542), .A2(W6459), .ZN(W13733));
  NOR2X1 G1657 (.A1(I546), .A2(W5743), .ZN(W13732));
  NOR2X1 G1658 (.A1(W18400), .A2(W226), .ZN(W29965));
  NOR2X1 G1659 (.A1(W27798), .A2(W7774), .ZN(W37103));
  NOR2X1 G1660 (.A1(W14912), .A2(W20541), .ZN(W20796));
  NOR2X1 G1661 (.A1(W1175), .A2(W1713), .ZN(W13756));
  NOR2X1 G1662 (.A1(W8627), .A2(W28646), .ZN(W29982));
  NOR2X1 G1663 (.A1(W6533), .A2(W29483), .ZN(W37068));
  NOR2X1 G1664 (.A1(I1667), .A2(W2224), .ZN(W13762));
  NOR2X1 G1665 (.A1(W13290), .A2(W2408), .ZN(O782));
  NOR2X1 G1666 (.A1(W18478), .A2(W15200), .ZN(W20784));
  NOR2X1 G1667 (.A1(W22202), .A2(W33066), .ZN(W37072));
  NOR2X1 G1668 (.A1(W16694), .A2(I1385), .ZN(O2082));
  NOR2X1 G1669 (.A1(W13348), .A2(W12169), .ZN(W13757));
  NOR2X1 G1670 (.A1(W13715), .A2(W7733), .ZN(W37510));
  NOR2X1 G1671 (.A1(W19991), .A2(W7102), .ZN(O8764));
  NOR2X1 G1672 (.A1(W6583), .A2(W1863), .ZN(W13753));
  NOR2X1 G1673 (.A1(W24606), .A2(W7290), .ZN(O5139));
  NOR2X1 G1674 (.A1(W7466), .A2(W7303), .ZN(W13751));
  NOR2X1 G1675 (.A1(W32118), .A2(W34877), .ZN(O8767));
  NOR2X1 G1676 (.A1(W13198), .A2(W13248), .ZN(W29977));
  NOR2X1 G1677 (.A1(W1575), .A2(W7689), .ZN(O8769));
  NOR2X1 G1678 (.A1(W7989), .A2(W5496), .ZN(W12919));
  NOR2X1 G1679 (.A1(W13166), .A2(W4894), .ZN(W29719));
  NOR2X1 G1680 (.A1(W17991), .A2(W3482), .ZN(W21040));
  NOR2X1 G1681 (.A1(W5310), .A2(W4036), .ZN(W12926));
  NOR2X1 G1682 (.A1(W26332), .A2(I1617), .ZN(W37899));
  NOR2X1 G1683 (.A1(W11993), .A2(W8259), .ZN(W12924));
  NOR2X1 G1684 (.A1(W5945), .A2(W2769), .ZN(O665));
  NOR2X1 G1685 (.A1(W2229), .A2(W24858), .ZN(O9265));
  NOR2X1 G1686 (.A1(W8959), .A2(W3384), .ZN(W12920));
  NOR2X1 G1687 (.A1(W15643), .A2(W31788), .ZN(W37895));
  NOR2X1 G1688 (.A1(W5393), .A2(I1038), .ZN(O9266));
  NOR2X1 G1689 (.A1(I1367), .A2(I1273), .ZN(W12917));
  NOR2X1 G1690 (.A1(W26398), .A2(W26433), .ZN(W29715));
  NOR2X1 G1691 (.A1(W24725), .A2(W7159), .ZN(O9267));
  NOR2X1 G1692 (.A1(W4236), .A2(W3461), .ZN(W21043));
  NOR2X1 G1693 (.A1(W12294), .A2(W3466), .ZN(W29714));
  NOR2X1 G1694 (.A1(W18424), .A2(W18051), .ZN(W21045));
  NOR2X1 G1695 (.A1(W1363), .A2(I1892), .ZN(W12911));
  NOR2X1 G1696 (.A1(W12166), .A2(W15405), .ZN(O9253));
  NOR2X1 G1697 (.A1(I1428), .A2(W10311), .ZN(W12947));
  NOR2X1 G1698 (.A1(W6531), .A2(W8702), .ZN(W12946));
  NOR2X1 G1699 (.A1(W10697), .A2(W17922), .ZN(W29723));
  NOR2X1 G1700 (.A1(W10624), .A2(W33514), .ZN(O9250));
  NOR2X1 G1701 (.A1(W8552), .A2(W12005), .ZN(W12943));
  NOR2X1 G1702 (.A1(W9775), .A2(W25111), .ZN(O9251));
  NOR2X1 G1703 (.A1(W152), .A2(W9248), .ZN(W12941));
  NOR2X1 G1704 (.A1(W26627), .A2(W27103), .ZN(O9252));
  NOR2X1 G1705 (.A1(I62), .A2(W10868), .ZN(W29711));
  NOR2X1 G1706 (.A1(W25400), .A2(I1744), .ZN(O9254));
  NOR2X1 G1707 (.A1(W14418), .A2(W34891), .ZN(O9256));
  NOR2X1 G1708 (.A1(W8955), .A2(W4280), .ZN(O666));
  NOR2X1 G1709 (.A1(W2113), .A2(W817), .ZN(W12933));
  NOR2X1 G1710 (.A1(W23062), .A2(W27837), .ZN(O9258));
  NOR2X1 G1711 (.A1(W12024), .A2(W660), .ZN(W12931));
  NOR2X1 G1712 (.A1(W7696), .A2(W20570), .ZN(O5015));
  NOR2X1 G1713 (.A1(W32090), .A2(W9765), .ZN(W37951));
  NOR2X1 G1714 (.A1(W7467), .A2(W17464), .ZN(W29705));
  NOR2X1 G1715 (.A1(W2924), .A2(W5422), .ZN(W12888));
  NOR2X1 G1716 (.A1(W2705), .A2(W969), .ZN(O661));
  NOR2X1 G1717 (.A1(W11777), .A2(W6112), .ZN(O2141));
  NOR2X1 G1718 (.A1(W3502), .A2(W10875), .ZN(O5010));
  NOR2X1 G1719 (.A1(I639), .A2(W25848), .ZN(O9292));
  NOR2X1 G1720 (.A1(W5377), .A2(W11181), .ZN(W12883));
  NOR2X1 G1721 (.A1(W33934), .A2(W29509), .ZN(O9293));
  NOR2X1 G1722 (.A1(I1271), .A2(W4026), .ZN(W12890));
  NOR2X1 G1723 (.A1(W9012), .A2(W14119), .ZN(O5009));
  NOR2X1 G1724 (.A1(W4114), .A2(W10505), .ZN(W21058));
  NOR2X1 G1725 (.A1(W19802), .A2(W8077), .ZN(W21059));
  NOR2X1 G1726 (.A1(W3275), .A2(W11527), .ZN(O5008));
  NOR2X1 G1727 (.A1(W2814), .A2(W9338), .ZN(W12875));
  NOR2X1 G1728 (.A1(W2667), .A2(W19776), .ZN(O9298));
  NOR2X1 G1729 (.A1(W7523), .A2(W10878), .ZN(W12872));
  NOR2X1 G1730 (.A1(W36210), .A2(W26600), .ZN(W37962));
  NOR2X1 G1731 (.A1(W31018), .A2(W14963), .ZN(W37929));
  NOR2X1 G1732 (.A1(W4577), .A2(W5517), .ZN(W37914));
  NOR2X1 G1733 (.A1(W15058), .A2(W10191), .ZN(O9276));
  NOR2X1 G1734 (.A1(W28925), .A2(W1577), .ZN(W29710));
  NOR2X1 G1735 (.A1(W36428), .A2(W8470), .ZN(O9277));
  NOR2X1 G1736 (.A1(W21840), .A2(W15674), .ZN(O9278));
  NOR2X1 G1737 (.A1(W36202), .A2(W23091), .ZN(W37923));
  NOR2X1 G1738 (.A1(W24519), .A2(I1569), .ZN(W37926));
  NOR2X1 G1739 (.A1(W12761), .A2(W8858), .ZN(W12901));
  NOR2X1 G1740 (.A1(W18476), .A2(W3344), .ZN(W21034));
  NOR2X1 G1741 (.A1(W28934), .A2(W2961), .ZN(W37932));
  NOR2X1 G1742 (.A1(W9508), .A2(W1526), .ZN(O9284));
  NOR2X1 G1743 (.A1(W13722), .A2(W9887), .ZN(O2139));
  NOR2X1 G1744 (.A1(W12269), .A2(W12180), .ZN(W12895));
  NOR2X1 G1745 (.A1(W18887), .A2(W13980), .ZN(W21051));
  NOR2X1 G1746 (.A1(W33737), .A2(W6159), .ZN(W37941));
  NOR2X1 G1747 (.A1(W4433), .A2(W4400), .ZN(W37942));
  NOR2X1 G1748 (.A1(W95), .A2(W5569), .ZN(W12994));
  NOR2X1 G1749 (.A1(W3914), .A2(W5581), .ZN(W13002));
  NOR2X1 G1750 (.A1(W19115), .A2(W21567), .ZN(O5021));
  NOR2X1 G1751 (.A1(W10564), .A2(W1252), .ZN(W29740));
  NOR2X1 G1752 (.A1(W4169), .A2(W3700), .ZN(W29739));
  NOR2X1 G1753 (.A1(W15378), .A2(W33500), .ZN(W37837));
  NOR2X1 G1754 (.A1(W29702), .A2(W4366), .ZN(W29738));
  NOR2X1 G1755 (.A1(W24226), .A2(W2163), .ZN(O9224));
  NOR2X1 G1756 (.A1(W18348), .A2(W8660), .ZN(W21022));
  NOR2X1 G1757 (.A1(W431), .A2(W18607), .ZN(O9219));
  NOR2X1 G1758 (.A1(W4049), .A2(W7472), .ZN(W12993));
  NOR2X1 G1759 (.A1(W26393), .A2(W18097), .ZN(O9225));
  NOR2X1 G1760 (.A1(W11529), .A2(W6231), .ZN(W12991));
  NOR2X1 G1761 (.A1(W28946), .A2(W23405), .ZN(O5020));
  NOR2X1 G1762 (.A1(I499), .A2(W1458), .ZN(O677));
  NOR2X1 G1763 (.A1(W9672), .A2(W24615), .ZN(O9227));
  NOR2X1 G1764 (.A1(W17311), .A2(W9651), .ZN(W21024));
  NOR2X1 G1765 (.A1(W5693), .A2(I26), .ZN(W12986));
  NOR2X1 G1766 (.A1(W17364), .A2(W14551), .ZN(W29743));
  NOR2X1 G1767 (.A1(W13641), .A2(W13442), .ZN(W21012));
  NOR2X1 G1768 (.A1(W20063), .A2(W12612), .ZN(O9211));
  NOR2X1 G1769 (.A1(W28930), .A2(W15002), .ZN(O5023));
  NOR2X1 G1770 (.A1(W812), .A2(W1844), .ZN(W13017));
  NOR2X1 G1771 (.A1(W16883), .A2(W20017), .ZN(W37823));
  NOR2X1 G1772 (.A1(I1579), .A2(W5315), .ZN(W13015));
  NOR2X1 G1773 (.A1(W10708), .A2(I54), .ZN(W13014));
  NOR2X1 G1774 (.A1(W15313), .A2(W25792), .ZN(W37825));
  NOR2X1 G1775 (.A1(W16722), .A2(W11469), .ZN(O9228));
  NOR2X1 G1776 (.A1(W5741), .A2(W12201), .ZN(O680));
  NOR2X1 G1777 (.A1(W1151), .A2(W6691), .ZN(W13009));
  NOR2X1 G1778 (.A1(W10950), .A2(W8826), .ZN(W13008));
  NOR2X1 G1779 (.A1(W27714), .A2(I1968), .ZN(O9214));
  NOR2X1 G1780 (.A1(W1906), .A2(W2449), .ZN(W13006));
  NOR2X1 G1781 (.A1(W24270), .A2(W27728), .ZN(O9217));
  NOR2X1 G1782 (.A1(W20685), .A2(W12005), .ZN(W21017));
  NOR2X1 G1783 (.A1(W3442), .A2(W870), .ZN(W12957));
  NOR2X1 G1784 (.A1(W6452), .A2(W1827), .ZN(W12965));
  NOR2X1 G1785 (.A1(W20262), .A2(W12365), .ZN(W21032));
  NOR2X1 G1786 (.A1(W3155), .A2(W5004), .ZN(W12963));
  NOR2X1 G1787 (.A1(W15974), .A2(W42), .ZN(O9245));
  NOR2X1 G1788 (.A1(W4847), .A2(W4986), .ZN(W12961));
  NOR2X1 G1789 (.A1(W1008), .A2(I1603), .ZN(W12960));
  NOR2X1 G1790 (.A1(W8891), .A2(W7959), .ZN(O672));
  NOR2X1 G1791 (.A1(W4729), .A2(W2173), .ZN(W12958));
  NOR2X1 G1792 (.A1(W26404), .A2(W28598), .ZN(W29728));
  NOR2X1 G1793 (.A1(W12505), .A2(W7984), .ZN(W12956));
  NOR2X1 G1794 (.A1(I1073), .A2(W12894), .ZN(W12955));
  NOR2X1 G1795 (.A1(I1737), .A2(W3736), .ZN(W12954));
  NOR2X1 G1796 (.A1(W5083), .A2(W5143), .ZN(W12953));
  NOR2X1 G1797 (.A1(W2615), .A2(W29541), .ZN(O5016));
  NOR2X1 G1798 (.A1(W976), .A2(W9989), .ZN(W12951));
  NOR2X1 G1799 (.A1(I1246), .A2(W11296), .ZN(W12950));
  NOR2X1 G1800 (.A1(W8001), .A2(W4599), .ZN(O9247));
  NOR2X1 G1801 (.A1(W5336), .A2(W8624), .ZN(W12975));
  NOR2X1 G1802 (.A1(W8608), .A2(W6748), .ZN(O5018));
  NOR2X1 G1803 (.A1(W36484), .A2(W1815), .ZN(O9233));
  NOR2X1 G1804 (.A1(W4338), .A2(W8057), .ZN(W12981));
  NOR2X1 G1805 (.A1(W11151), .A2(W12547), .ZN(W12980));
  NOR2X1 G1806 (.A1(W5718), .A2(W12739), .ZN(W12979));
  NOR2X1 G1807 (.A1(W11481), .A2(W5105), .ZN(W29732));
  NOR2X1 G1808 (.A1(W11986), .A2(W5692), .ZN(W12977));
  NOR2X1 G1809 (.A1(W23219), .A2(W26952), .ZN(W29731));
  NOR2X1 G1810 (.A1(I446), .A2(W5100), .ZN(W12870));
  NOR2X1 G1811 (.A1(I1966), .A2(W12521), .ZN(W12974));
  NOR2X1 G1812 (.A1(W4377), .A2(W11555), .ZN(W37859));
  NOR2X1 G1813 (.A1(W11061), .A2(W228), .ZN(W12972));
  NOR2X1 G1814 (.A1(W10978), .A2(W249), .ZN(O673));
  NOR2X1 G1815 (.A1(I1916), .A2(W31210), .ZN(O9239));
  NOR2X1 G1816 (.A1(W9228), .A2(W29552), .ZN(W29729));
  NOR2X1 G1817 (.A1(W671), .A2(I1506), .ZN(W12967));
  NOR2X1 G1818 (.A1(W26498), .A2(W8520), .ZN(W38055));
  NOR2X1 G1819 (.A1(W3040), .A2(W11222), .ZN(W38051));
  NOR2X1 G1820 (.A1(W33275), .A2(W20709), .ZN(O9347));
  NOR2X1 G1821 (.A1(W43), .A2(W14012), .ZN(W29661));
  NOR2X1 G1822 (.A1(W2488), .A2(W6111), .ZN(W12770));
  NOR2X1 G1823 (.A1(W11046), .A2(W4509), .ZN(O647));
  NOR2X1 G1824 (.A1(W30490), .A2(W17954), .ZN(W38054));
  NOR2X1 G1825 (.A1(W397), .A2(W6153), .ZN(W12767));
  NOR2X1 G1826 (.A1(W2022), .A2(W2614), .ZN(O646));
  NOR2X1 G1827 (.A1(W4235), .A2(W6413), .ZN(W12774));
  NOR2X1 G1828 (.A1(W18279), .A2(W13673), .ZN(W38056));
  NOR2X1 G1829 (.A1(W3873), .A2(W7782), .ZN(W12763));
  NOR2X1 G1830 (.A1(W2184), .A2(W27978), .ZN(O9351));
  NOR2X1 G1831 (.A1(W11109), .A2(W4579), .ZN(O2148));
  NOR2X1 G1832 (.A1(W9487), .A2(W36710), .ZN(W38062));
  NOR2X1 G1833 (.A1(W9620), .A2(W3575), .ZN(W12759));
  NOR2X1 G1834 (.A1(W24482), .A2(W21920), .ZN(O9352));
  NOR2X1 G1835 (.A1(W5906), .A2(W10867), .ZN(W12757));
  NOR2X1 G1836 (.A1(W3383), .A2(W11283), .ZN(O9344));
  NOR2X1 G1837 (.A1(W8372), .A2(W11393), .ZN(O9336));
  NOR2X1 G1838 (.A1(W1857), .A2(W24018), .ZN(W38032));
  NOR2X1 G1839 (.A1(W8483), .A2(W26114), .ZN(O4995));
  NOR2X1 G1840 (.A1(I999), .A2(W10697), .ZN(W21089));
  NOR2X1 G1841 (.A1(W494), .A2(W5108), .ZN(O9337));
  NOR2X1 G1842 (.A1(W25683), .A2(W5715), .ZN(W29668));
  NOR2X1 G1843 (.A1(W12010), .A2(W16590), .ZN(W29667));
  NOR2X1 G1844 (.A1(W21236), .A2(W18165), .ZN(O9341));
  NOR2X1 G1845 (.A1(W25586), .A2(W15680), .ZN(W29660));
  NOR2X1 G1846 (.A1(W9721), .A2(W9674), .ZN(O648));
  NOR2X1 G1847 (.A1(W28995), .A2(W6123), .ZN(W29664));
  NOR2X1 G1848 (.A1(W2609), .A2(W19486), .ZN(W21095));
  NOR2X1 G1849 (.A1(W28459), .A2(W22308), .ZN(O9346));
  NOR2X1 G1850 (.A1(W25891), .A2(W11226), .ZN(W38049));
  NOR2X1 G1851 (.A1(I1806), .A2(I647), .ZN(W12776));
  NOR2X1 G1852 (.A1(W13102), .A2(I1014), .ZN(W29662));
  NOR2X1 G1853 (.A1(W17326), .A2(W992), .ZN(O9372));
  NOR2X1 G1854 (.A1(W15184), .A2(W1271), .ZN(O4993));
  NOR2X1 G1855 (.A1(W8903), .A2(W17473), .ZN(W21110));
  NOR2X1 G1856 (.A1(W18433), .A2(W19878), .ZN(W21111));
  NOR2X1 G1857 (.A1(W22838), .A2(W23460), .ZN(W38094));
  NOR2X1 G1858 (.A1(W12946), .A2(W22714), .ZN(O9369));
  NOR2X1 G1859 (.A1(W17326), .A2(W24787), .ZN(O4991));
  NOR2X1 G1860 (.A1(I551), .A2(W11191), .ZN(W12726));
  NOR2X1 G1861 (.A1(W21215), .A2(W29125), .ZN(O9371));
  NOR2X1 G1862 (.A1(W13163), .A2(W17135), .ZN(O9366));
  NOR2X1 G1863 (.A1(W2974), .A2(W11819), .ZN(W12723));
  NOR2X1 G1864 (.A1(W1334), .A2(W18844), .ZN(O9373));
  NOR2X1 G1865 (.A1(W16815), .A2(W18852), .ZN(W21114));
  NOR2X1 G1866 (.A1(W1007), .A2(W8454), .ZN(W12719));
  NOR2X1 G1867 (.A1(W8593), .A2(W7805), .ZN(W12718));
  NOR2X1 G1868 (.A1(W5923), .A2(W1220), .ZN(O9376));
  NOR2X1 G1869 (.A1(W21233), .A2(W37455), .ZN(O9377));
  NOR2X1 G1870 (.A1(I438), .A2(W7295), .ZN(W12714));
  NOR2X1 G1871 (.A1(W26202), .A2(W8622), .ZN(O9363));
  NOR2X1 G1872 (.A1(W6226), .A2(W10414), .ZN(W12754));
  NOR2X1 G1873 (.A1(W7128), .A2(W725), .ZN(O9357));
  NOR2X1 G1874 (.A1(W32419), .A2(W31316), .ZN(O9358));
  NOR2X1 G1875 (.A1(W31830), .A2(W35813), .ZN(W38072));
  NOR2X1 G1876 (.A1(W26003), .A2(W1315), .ZN(W38074));
  NOR2X1 G1877 (.A1(W25837), .A2(W10565), .ZN(W38076));
  NOR2X1 G1878 (.A1(W14921), .A2(W6231), .ZN(O2150));
  NOR2X1 G1879 (.A1(W10693), .A2(W15073), .ZN(W21104));
  NOR2X1 G1880 (.A1(W7803), .A2(W4322), .ZN(W12793));
  NOR2X1 G1881 (.A1(W25931), .A2(W15865), .ZN(O9364));
  NOR2X1 G1882 (.A1(W5644), .A2(W15869), .ZN(W21106));
  NOR2X1 G1883 (.A1(W12420), .A2(W8941), .ZN(O644));
  NOR2X1 G1884 (.A1(W4640), .A2(W2653), .ZN(W12739));
  NOR2X1 G1885 (.A1(W21231), .A2(W20578), .ZN(O9365));
  NOR2X1 G1886 (.A1(W1853), .A2(I1450), .ZN(O643));
  NOR2X1 G1887 (.A1(W12132), .A2(W16961), .ZN(W21107));
  NOR2X1 G1888 (.A1(W502), .A2(W5605), .ZN(W12841));
  NOR2X1 G1889 (.A1(W8668), .A2(W21620), .ZN(W29688));
  NOR2X1 G1890 (.A1(W4988), .A2(W6368), .ZN(W12849));
  NOR2X1 G1891 (.A1(W12469), .A2(W157), .ZN(W12848));
  NOR2X1 G1892 (.A1(W4988), .A2(W6909), .ZN(W12846));
  NOR2X1 G1893 (.A1(W4624), .A2(W5113), .ZN(O9306));
  NOR2X1 G1894 (.A1(I408), .A2(W12246), .ZN(W12844));
  NOR2X1 G1895 (.A1(W24817), .A2(W35508), .ZN(O9309));
  NOR2X1 G1896 (.A1(W619), .A2(W15602), .ZN(O5002));
  NOR2X1 G1897 (.A1(W455), .A2(W8789), .ZN(W21069));
  NOR2X1 G1898 (.A1(W867), .A2(W4171), .ZN(W12840));
  NOR2X1 G1899 (.A1(W32861), .A2(W21082), .ZN(W37987));
  NOR2X1 G1900 (.A1(W4967), .A2(W3344), .ZN(W12838));
  NOR2X1 G1901 (.A1(W37919), .A2(W7498), .ZN(O9311));
  NOR2X1 G1902 (.A1(W17705), .A2(W23509), .ZN(W37990));
  NOR2X1 G1903 (.A1(W6806), .A2(W8768), .ZN(W12835));
  NOR2X1 G1904 (.A1(W8230), .A2(W7942), .ZN(O659));
  NOR2X1 G1905 (.A1(W8185), .A2(W2297), .ZN(W12832));
  NOR2X1 G1906 (.A1(W26353), .A2(W662), .ZN(W29692));
  NOR2X1 G1907 (.A1(W10442), .A2(W12087), .ZN(W12869));
  NOR2X1 G1908 (.A1(W27735), .A2(W28648), .ZN(O9299));
  NOR2X1 G1909 (.A1(W1901), .A2(W8290), .ZN(W21062));
  NOR2X1 G1910 (.A1(W3897), .A2(W8604), .ZN(W12866));
  NOR2X1 G1911 (.A1(W4087), .A2(W4274), .ZN(W12865));
  NOR2X1 G1912 (.A1(W20474), .A2(W18916), .ZN(W29695));
  NOR2X1 G1913 (.A1(W20882), .A2(W9177), .ZN(W29694));
  NOR2X1 G1914 (.A1(W7046), .A2(W10374), .ZN(W12861));
  NOR2X1 G1915 (.A1(W10283), .A2(W8977), .ZN(W12830));
  NOR2X1 G1916 (.A1(I1188), .A2(I1272), .ZN(W12859));
  NOR2X1 G1917 (.A1(I412), .A2(W3701), .ZN(W12858));
  NOR2X1 G1918 (.A1(W30335), .A2(W10830), .ZN(O9301));
  NOR2X1 G1919 (.A1(I1354), .A2(W9509), .ZN(W12856));
  NOR2X1 G1920 (.A1(W6084), .A2(W11047), .ZN(W12855));
  NOR2X1 G1921 (.A1(W11995), .A2(W3354), .ZN(W29691));
  NOR2X1 G1922 (.A1(W7365), .A2(W9264), .ZN(W37975));
  NOR2X1 G1923 (.A1(W5854), .A2(W122), .ZN(W12803));
  NOR2X1 G1924 (.A1(W4646), .A2(W9109), .ZN(O654));
  NOR2X1 G1925 (.A1(W20831), .A2(W1316), .ZN(W21084));
  NOR2X1 G1926 (.A1(W26213), .A2(W23279), .ZN(O9330));
  NOR2X1 G1927 (.A1(I1940), .A2(W1158), .ZN(W12808));
  NOR2X1 G1928 (.A1(W12699), .A2(W10599), .ZN(W12807));
  NOR2X1 G1929 (.A1(W8545), .A2(W11359), .ZN(W12806));
  NOR2X1 G1930 (.A1(W25732), .A2(W13492), .ZN(O9331));
  NOR2X1 G1931 (.A1(I1015), .A2(W10459), .ZN(W12804));
  NOR2X1 G1932 (.A1(W2481), .A2(W11729), .ZN(W21083));
  NOR2X1 G1933 (.A1(W435), .A2(W8240), .ZN(W12802));
  NOR2X1 G1934 (.A1(W16642), .A2(W7708), .ZN(W21086));
  NOR2X1 G1935 (.A1(W9885), .A2(W34392), .ZN(W38024));
  NOR2X1 G1936 (.A1(W7968), .A2(W35442), .ZN(W38025));
  NOR2X1 G1937 (.A1(W3201), .A2(W14586), .ZN(O9333));
  NOR2X1 G1938 (.A1(W2205), .A2(W5702), .ZN(W12796));
  NOR2X1 G1939 (.A1(W2452), .A2(W4909), .ZN(O4998));
  NOR2X1 G1940 (.A1(W32320), .A2(W16831), .ZN(O9335));
  NOR2X1 G1941 (.A1(W9007), .A2(I616), .ZN(W12820));
  NOR2X1 G1942 (.A1(W16073), .A2(W2060), .ZN(O2144));
  NOR2X1 G1943 (.A1(W6903), .A2(W9943), .ZN(W12828));
  NOR2X1 G1944 (.A1(W20500), .A2(W17374), .ZN(W21076));
  NOR2X1 G1945 (.A1(W20192), .A2(W23155), .ZN(O9317));
  NOR2X1 G1946 (.A1(W17515), .A2(W24795), .ZN(W29682));
  NOR2X1 G1947 (.A1(W20126), .A2(W23646), .ZN(O9321));
  NOR2X1 G1948 (.A1(W14791), .A2(W12661), .ZN(W21079));
  NOR2X1 G1949 (.A1(W4018), .A2(W779), .ZN(W21080));
  NOR2X1 G1950 (.A1(W3626), .A2(W7185), .ZN(W13022));
  NOR2X1 G1951 (.A1(W7167), .A2(W23587), .ZN(W29678));
  NOR2X1 G1952 (.A1(W20386), .A2(W13427), .ZN(O9323));
  NOR2X1 G1953 (.A1(W9968), .A2(W3157), .ZN(W38010));
  NOR2X1 G1954 (.A1(W17283), .A2(W5488), .ZN(W38012));
  NOR2X1 G1955 (.A1(W9387), .A2(W14043), .ZN(W29676));
  NOR2X1 G1956 (.A1(W12757), .A2(I158), .ZN(W12814));
  NOR2X1 G1957 (.A1(W12663), .A2(W1715), .ZN(W12813));
  NOR2X1 G1958 (.A1(W7078), .A2(W10561), .ZN(W13229));
  NOR2X1 G1959 (.A1(W5122), .A2(W12790), .ZN(W13237));
  NOR2X1 G1960 (.A1(W11937), .A2(W2142), .ZN(W13236));
  NOR2X1 G1961 (.A1(W33853), .A2(I1895), .ZN(W37597));
  NOR2X1 G1962 (.A1(W15317), .A2(W3161), .ZN(W29812));
  NOR2X1 G1963 (.A1(W4456), .A2(W10270), .ZN(W13233));
  NOR2X1 G1964 (.A1(I1666), .A2(W10538), .ZN(O713));
  NOR2X1 G1965 (.A1(W9247), .A2(W13968), .ZN(W20947));
  NOR2X1 G1966 (.A1(W7670), .A2(W10419), .ZN(W13230));
  NOR2X1 G1967 (.A1(W18423), .A2(W13275), .ZN(W37595));
  NOR2X1 G1968 (.A1(W10792), .A2(W26229), .ZN(O9073));
  NOR2X1 G1969 (.A1(W7149), .A2(W6019), .ZN(O9076));
  NOR2X1 G1970 (.A1(I1682), .A2(W4898), .ZN(W20949));
  NOR2X1 G1971 (.A1(W3369), .A2(W2344), .ZN(W13224));
  NOR2X1 G1972 (.A1(W9744), .A2(W2130), .ZN(W13223));
  NOR2X1 G1973 (.A1(I1675), .A2(W11464), .ZN(W37612));
  NOR2X1 G1974 (.A1(W20254), .A2(W23684), .ZN(O9079));
  NOR2X1 G1975 (.A1(I116), .A2(W4763), .ZN(W37615));
  NOR2X1 G1976 (.A1(W21822), .A2(W939), .ZN(O9067));
  NOR2X1 G1977 (.A1(W8229), .A2(W6351), .ZN(O5062));
  NOR2X1 G1978 (.A1(W6888), .A2(W9109), .ZN(W13255));
  NOR2X1 G1979 (.A1(W13403), .A2(I1809), .ZN(W20941));
  NOR2X1 G1980 (.A1(I933), .A2(W12010), .ZN(O719));
  NOR2X1 G1981 (.A1(W20019), .A2(W331), .ZN(W20942));
  NOR2X1 G1982 (.A1(W583), .A2(W5864), .ZN(W20943));
  NOR2X1 G1983 (.A1(W483), .A2(W14768), .ZN(O5057));
  NOR2X1 G1984 (.A1(W30743), .A2(W11671), .ZN(O9066));
  NOR2X1 G1985 (.A1(W14998), .A2(W26262), .ZN(W29807));
  NOR2X1 G1986 (.A1(W11058), .A2(W4256), .ZN(W13246));
  NOR2X1 G1987 (.A1(W12137), .A2(W34267), .ZN(W37592));
  NOR2X1 G1988 (.A1(I890), .A2(W6812), .ZN(W13244));
  NOR2X1 G1989 (.A1(W5836), .A2(W12498), .ZN(O717));
  NOR2X1 G1990 (.A1(W28221), .A2(W4856), .ZN(O9068));
  NOR2X1 G1991 (.A1(W9182), .A2(W641), .ZN(O716));
  NOR2X1 G1992 (.A1(W19931), .A2(W22347), .ZN(O9069));
  NOR2X1 G1993 (.A1(W11516), .A2(W33888), .ZN(O9092));
  NOR2X1 G1994 (.A1(W31197), .A2(I1512), .ZN(O9086));
  NOR2X1 G1995 (.A1(W9455), .A2(W12168), .ZN(W13199));
  NOR2X1 G1996 (.A1(W19227), .A2(W11171), .ZN(O2120));
  NOR2X1 G1997 (.A1(W11315), .A2(W7991), .ZN(W13197));
  NOR2X1 G1998 (.A1(W241), .A2(I485), .ZN(O9088));
  NOR2X1 G1999 (.A1(W18402), .A2(W28442), .ZN(O9089));
  NOR2X1 G2000 (.A1(W11437), .A2(W20004), .ZN(O9090));
  NOR2X1 G2001 (.A1(I158), .A2(W4086), .ZN(O9091));
  NOR2X1 G2002 (.A1(W36247), .A2(W27221), .ZN(W37626));
  NOR2X1 G2003 (.A1(W7429), .A2(W1233), .ZN(W13190));
  NOR2X1 G2004 (.A1(I309), .A2(W7530), .ZN(W13189));
  NOR2X1 G2005 (.A1(I334), .A2(I1703), .ZN(W13188));
  NOR2X1 G2006 (.A1(W5043), .A2(W12098), .ZN(W13187));
  NOR2X1 G2007 (.A1(W3576), .A2(W12544), .ZN(O2121));
  NOR2X1 G2008 (.A1(W6507), .A2(W7160), .ZN(O9097));
  NOR2X1 G2009 (.A1(W8703), .A2(W941), .ZN(O708));
  NOR2X1 G2010 (.A1(I1014), .A2(W28599), .ZN(W37642));
  NOR2X1 G2011 (.A1(W10152), .A2(W10165), .ZN(W20954));
  NOR2X1 G2012 (.A1(W19448), .A2(W7282), .ZN(W20952));
  NOR2X1 G2013 (.A1(W5286), .A2(W11613), .ZN(W13216));
  NOR2X1 G2014 (.A1(W7565), .A2(W1377), .ZN(O712));
  NOR2X1 G2015 (.A1(W13586), .A2(W24011), .ZN(W37618));
  NOR2X1 G2016 (.A1(W13203), .A2(W9093), .ZN(W13213));
  NOR2X1 G2017 (.A1(W8134), .A2(W35126), .ZN(O9082));
  NOR2X1 G2018 (.A1(W9779), .A2(W2794), .ZN(W13211));
  NOR2X1 G2019 (.A1(W2342), .A2(W7287), .ZN(W20953));
  NOR2X1 G2020 (.A1(W173), .A2(W19177), .ZN(W37579));
  NOR2X1 G2021 (.A1(W7950), .A2(W14766), .ZN(O9084));
  NOR2X1 G2022 (.A1(I884), .A2(W3931), .ZN(W13207));
  NOR2X1 G2023 (.A1(I1784), .A2(W3597), .ZN(W13206));
  NOR2X1 G2024 (.A1(W14465), .A2(W17292), .ZN(W20955));
  NOR2X1 G2025 (.A1(W3514), .A2(W5620), .ZN(W13204));
  NOR2X1 G2026 (.A1(W2769), .A2(W23240), .ZN(W37625));
  NOR2X1 G2027 (.A1(W10637), .A2(W9107), .ZN(W13202));
  NOR2X1 G2028 (.A1(W7764), .A2(I738), .ZN(W13306));
  NOR2X1 G2029 (.A1(W4534), .A2(W12508), .ZN(W13316));
  NOR2X1 G2030 (.A1(W9460), .A2(W6642), .ZN(W13315));
  NOR2X1 G2031 (.A1(W19175), .A2(W26579), .ZN(O9032));
  NOR2X1 G2032 (.A1(W24812), .A2(W14412), .ZN(O5075));
  NOR2X1 G2033 (.A1(W13150), .A2(W22312), .ZN(O5070));
  NOR2X1 G2034 (.A1(W3059), .A2(W3258), .ZN(W20927));
  NOR2X1 G2035 (.A1(W258), .A2(W22212), .ZN(W29833));
  NOR2X1 G2036 (.A1(W12499), .A2(W12090), .ZN(W13307));
  NOR2X1 G2037 (.A1(W15939), .A2(W144), .ZN(O9031));
  NOR2X1 G2038 (.A1(W4392), .A2(W11469), .ZN(W13304));
  NOR2X1 G2039 (.A1(W29146), .A2(W7135), .ZN(O5068));
  NOR2X1 G2040 (.A1(W25178), .A2(W10108), .ZN(O9041));
  NOR2X1 G2041 (.A1(W34997), .A2(W22393), .ZN(W37545));
  NOR2X1 G2042 (.A1(W13158), .A2(W12560), .ZN(W13300));
  NOR2X1 G2043 (.A1(I1208), .A2(W10228), .ZN(W13299));
  NOR2X1 G2044 (.A1(W19841), .A2(W21252), .ZN(O9042));
  NOR2X1 G2045 (.A1(W3208), .A2(I1924), .ZN(O5066));
  NOR2X1 G2046 (.A1(I682), .A2(W18407), .ZN(W20919));
  NOR2X1 G2047 (.A1(W3460), .A2(W11582), .ZN(W13334));
  NOR2X1 G2048 (.A1(W6908), .A2(W8363), .ZN(W13333));
  NOR2X1 G2049 (.A1(W22360), .A2(W14852), .ZN(O9025));
  NOR2X1 G2050 (.A1(W10478), .A2(W3753), .ZN(O729));
  NOR2X1 G2051 (.A1(W17693), .A2(W19576), .ZN(W20917));
  NOR2X1 G2052 (.A1(W11823), .A2(W17663), .ZN(W20918));
  NOR2X1 G2053 (.A1(W24593), .A2(W18171), .ZN(W37517));
  NOR2X1 G2054 (.A1(I320), .A2(W11665), .ZN(W13326));
  NOR2X1 G2055 (.A1(I1526), .A2(I1843), .ZN(W13294));
  NOR2X1 G2056 (.A1(W9526), .A2(W31256), .ZN(O9028));
  NOR2X1 G2057 (.A1(W4519), .A2(I618), .ZN(W20920));
  NOR2X1 G2058 (.A1(W142), .A2(W695), .ZN(W13322));
  NOR2X1 G2059 (.A1(I1136), .A2(W2819), .ZN(O2108));
  NOR2X1 G2060 (.A1(I1166), .A2(W1499), .ZN(O5076));
  NOR2X1 G2061 (.A1(W10869), .A2(W8510), .ZN(O727));
  NOR2X1 G2062 (.A1(I459), .A2(W7555), .ZN(W13318));
  NOR2X1 G2063 (.A1(W22366), .A2(W29526), .ZN(O9058));
  NOR2X1 G2064 (.A1(W29574), .A2(W21013), .ZN(O9055));
  NOR2X1 G2065 (.A1(W11686), .A2(W795), .ZN(O722));
  NOR2X1 G2066 (.A1(W21235), .A2(W24176), .ZN(W37566));
  NOR2X1 G2067 (.A1(W27125), .A2(W24229), .ZN(W29822));
  NOR2X1 G2068 (.A1(W4575), .A2(W287), .ZN(W13270));
  NOR2X1 G2069 (.A1(W3383), .A2(W3615), .ZN(W13269));
  NOR2X1 G2070 (.A1(I815), .A2(W10037), .ZN(W13268));
  NOR2X1 G2071 (.A1(W2520), .A2(W9018), .ZN(W13267));
  NOR2X1 G2072 (.A1(W1292), .A2(W2631), .ZN(W37564));
  NOR2X1 G2073 (.A1(W10773), .A2(W10679), .ZN(W13265));
  NOR2X1 G2074 (.A1(W12425), .A2(W6496), .ZN(W13264));
  NOR2X1 G2075 (.A1(W9066), .A2(W7622), .ZN(W13263));
  NOR2X1 G2076 (.A1(W16127), .A2(W20717), .ZN(W37572));
  NOR2X1 G2077 (.A1(W32846), .A2(W401), .ZN(W37573));
  NOR2X1 G2078 (.A1(W1972), .A2(W31248), .ZN(O9059));
  NOR2X1 G2079 (.A1(W30067), .A2(W20593), .ZN(O9061));
  NOR2X1 G2080 (.A1(W879), .A2(W11171), .ZN(O720));
  NOR2X1 G2081 (.A1(W5816), .A2(W2919), .ZN(W37557));
  NOR2X1 G2082 (.A1(W11950), .A2(W8846), .ZN(O724));
  NOR2X1 G2083 (.A1(W27247), .A2(W19543), .ZN(W37554));
  NOR2X1 G2084 (.A1(W9417), .A2(W5685), .ZN(W13291));
  NOR2X1 G2085 (.A1(W10752), .A2(W5676), .ZN(O2114));
  NOR2X1 G2086 (.A1(W9859), .A2(W9263), .ZN(O723));
  NOR2X1 G2087 (.A1(W10239), .A2(W1878), .ZN(W13287));
  NOR2X1 G2088 (.A1(W5822), .A2(W9959), .ZN(W13286));
  NOR2X1 G2089 (.A1(W7997), .A2(W10058), .ZN(W13285));
  NOR2X1 G2090 (.A1(W11381), .A2(W12963), .ZN(W13182));
  NOR2X1 G2091 (.A1(W7667), .A2(I894), .ZN(W13283));
  NOR2X1 G2092 (.A1(I186), .A2(W35763), .ZN(O9049));
  NOR2X1 G2093 (.A1(W5257), .A2(W26406), .ZN(O9050));
  NOR2X1 G2094 (.A1(W8470), .A2(W381), .ZN(W13280));
  NOR2X1 G2095 (.A1(W14641), .A2(W35585), .ZN(O9051));
  NOR2X1 G2096 (.A1(W2060), .A2(W6756), .ZN(O5063));
  NOR2X1 G2097 (.A1(W1700), .A2(W1980), .ZN(W13277));
  NOR2X1 G2098 (.A1(W5864), .A2(W4017), .ZN(W13072));
  NOR2X1 G2099 (.A1(W33937), .A2(W6194), .ZN(O9168));
  NOR2X1 G2100 (.A1(W16661), .A2(W37208), .ZN(O9169));
  NOR2X1 G2101 (.A1(W8499), .A2(W2796), .ZN(O691));
  NOR2X1 G2102 (.A1(I767), .A2(W23250), .ZN(O9170));
  NOR2X1 G2103 (.A1(W12342), .A2(W16874), .ZN(O5034));
  NOR2X1 G2104 (.A1(W13634), .A2(W18863), .ZN(O9173));
  NOR2X1 G2105 (.A1(W639), .A2(W11952), .ZN(W37767));
  NOR2X1 G2106 (.A1(W18258), .A2(W33651), .ZN(O9177));
  NOR2X1 G2107 (.A1(W2175), .A2(I1108), .ZN(W13082));
  NOR2X1 G2108 (.A1(W4667), .A2(W14664), .ZN(W37771));
  NOR2X1 G2109 (.A1(I1280), .A2(W28308), .ZN(W29763));
  NOR2X1 G2110 (.A1(W11117), .A2(W1964), .ZN(W20998));
  NOR2X1 G2111 (.A1(W9038), .A2(W5457), .ZN(O688));
  NOR2X1 G2112 (.A1(W3497), .A2(W21945), .ZN(O9180));
  NOR2X1 G2113 (.A1(W829), .A2(W313), .ZN(W13065));
  NOR2X1 G2114 (.A1(W8408), .A2(W27669), .ZN(W29761));
  NOR2X1 G2115 (.A1(W4006), .A2(W26962), .ZN(W37778));
  NOR2X1 G2116 (.A1(W20962), .A2(W8439), .ZN(W29771));
  NOR2X1 G2117 (.A1(W15095), .A2(I1618), .ZN(W29777));
  NOR2X1 G2118 (.A1(W636), .A2(W9247), .ZN(W13101));
  NOR2X1 G2119 (.A1(W31872), .A2(W6204), .ZN(W37736));
  NOR2X1 G2120 (.A1(W4369), .A2(W8659), .ZN(W13099));
  NOR2X1 G2121 (.A1(W7657), .A2(W2295), .ZN(W13098));
  NOR2X1 G2122 (.A1(W2936), .A2(W10645), .ZN(W13096));
  NOR2X1 G2123 (.A1(W417), .A2(W3169), .ZN(W29772));
  NOR2X1 G2124 (.A1(W36667), .A2(W7671), .ZN(O9159));
  NOR2X1 G2125 (.A1(W11946), .A2(W963), .ZN(W13062));
  NOR2X1 G2126 (.A1(W11130), .A2(W10208), .ZN(W13091));
  NOR2X1 G2127 (.A1(W4274), .A2(W10895), .ZN(W13088));
  NOR2X1 G2128 (.A1(W25989), .A2(W3095), .ZN(O9164));
  NOR2X1 G2129 (.A1(W9891), .A2(W270), .ZN(O693));
  NOR2X1 G2130 (.A1(W25023), .A2(W33226), .ZN(O9166));
  NOR2X1 G2131 (.A1(W11390), .A2(W29150), .ZN(W37752));
  NOR2X1 G2132 (.A1(W6952), .A2(W3968), .ZN(W13083));
  NOR2X1 G2133 (.A1(W14261), .A2(W8685), .ZN(O2134));
  NOR2X1 G2134 (.A1(W8187), .A2(W632), .ZN(W37796));
  NOR2X1 G2135 (.A1(I1949), .A2(W5051), .ZN(W13043));
  NOR2X1 G2136 (.A1(I1992), .A2(W6857), .ZN(O685));
  NOR2X1 G2137 (.A1(W9602), .A2(W2336), .ZN(W37797));
  NOR2X1 G2138 (.A1(W20063), .A2(W19555), .ZN(O9195));
  NOR2X1 G2139 (.A1(W5178), .A2(W16304), .ZN(W37801));
  NOR2X1 G2140 (.A1(I476), .A2(W17635), .ZN(O9197));
  NOR2X1 G2141 (.A1(W12915), .A2(W5306), .ZN(W13035));
  NOR2X1 G2142 (.A1(W3408), .A2(W7834), .ZN(O2133));
  NOR2X1 G2143 (.A1(W23784), .A2(W9567), .ZN(O5029));
  NOR2X1 G2144 (.A1(W5708), .A2(W7586), .ZN(W13031));
  NOR2X1 G2145 (.A1(W10858), .A2(W3324), .ZN(O681));
  NOR2X1 G2146 (.A1(W5746), .A2(I388), .ZN(W13029));
  NOR2X1 G2147 (.A1(W2750), .A2(W23684), .ZN(O5027));
  NOR2X1 G2148 (.A1(W6889), .A2(I1694), .ZN(W13027));
  NOR2X1 G2149 (.A1(W13958), .A2(W13353), .ZN(W29752));
  NOR2X1 G2150 (.A1(W7726), .A2(W997), .ZN(W13024));
  NOR2X1 G2151 (.A1(W7613), .A2(W35228), .ZN(O9188));
  NOR2X1 G2152 (.A1(W10106), .A2(W11806), .ZN(W13061));
  NOR2X1 G2153 (.A1(W17042), .A2(W6696), .ZN(W21001));
  NOR2X1 G2154 (.A1(W2800), .A2(W35493), .ZN(O9183));
  NOR2X1 G2155 (.A1(W16444), .A2(W34897), .ZN(O9185));
  NOR2X1 G2156 (.A1(W18277), .A2(W7658), .ZN(W37785));
  NOR2X1 G2157 (.A1(W34194), .A2(W5006), .ZN(O9186));
  NOR2X1 G2158 (.A1(W13005), .A2(W33001), .ZN(W37787));
  NOR2X1 G2159 (.A1(W16153), .A2(I1031), .ZN(O9187));
  NOR2X1 G2160 (.A1(W5083), .A2(W934), .ZN(O9155));
  NOR2X1 G2161 (.A1(W31283), .A2(W17417), .ZN(O9189));
  NOR2X1 G2162 (.A1(W8826), .A2(W2265), .ZN(O9190));
  NOR2X1 G2163 (.A1(W22936), .A2(W29278), .ZN(O9192));
  NOR2X1 G2164 (.A1(W6606), .A2(W4546), .ZN(O686));
  NOR2X1 G2165 (.A1(W11278), .A2(W5255), .ZN(O9193));
  NOR2X1 G2166 (.A1(W469), .A2(W900), .ZN(W13047));
  NOR2X1 G2167 (.A1(W806), .A2(I216), .ZN(W13046));
  NOR2X1 G2168 (.A1(W10593), .A2(W12507), .ZN(W13152));
  NOR2X1 G2169 (.A1(W18223), .A2(W37304), .ZN(O9113));
  NOR2X1 G2170 (.A1(W9371), .A2(W6013), .ZN(W20965));
  NOR2X1 G2171 (.A1(W18124), .A2(W5775), .ZN(O9118));
  NOR2X1 G2172 (.A1(W6409), .A2(W4866), .ZN(O9119));
  NOR2X1 G2173 (.A1(I1980), .A2(W16055), .ZN(O9121));
  NOR2X1 G2174 (.A1(W2740), .A2(I144), .ZN(W13157));
  NOR2X1 G2175 (.A1(W8054), .A2(W11292), .ZN(W13155));
  NOR2X1 G2176 (.A1(W2465), .A2(W4246), .ZN(W20968));
  NOR2X1 G2177 (.A1(W11873), .A2(W10264), .ZN(O2122));
  NOR2X1 G2178 (.A1(W22683), .A2(W29537), .ZN(W37681));
  NOR2X1 G2179 (.A1(W6798), .A2(W7508), .ZN(W13150));
  NOR2X1 G2180 (.A1(W4900), .A2(W412), .ZN(O703));
  NOR2X1 G2181 (.A1(W27615), .A2(W19528), .ZN(W37682));
  NOR2X1 G2182 (.A1(W25495), .A2(W22702), .ZN(W37685));
  NOR2X1 G2183 (.A1(W12417), .A2(W8328), .ZN(W13144));
  NOR2X1 G2184 (.A1(I1934), .A2(W12014), .ZN(O2123));
  NOR2X1 G2185 (.A1(W631), .A2(W3684), .ZN(O9130));
  NOR2X1 G2186 (.A1(W33262), .A2(W19758), .ZN(O9103));
  NOR2X1 G2187 (.A1(W17961), .A2(W9760), .ZN(O9099));
  NOR2X1 G2188 (.A1(W1909), .A2(W5948), .ZN(W13179));
  NOR2X1 G2189 (.A1(W17229), .A2(W31440), .ZN(O9100));
  NOR2X1 G2190 (.A1(W17741), .A2(W3877), .ZN(W37649));
  NOR2X1 G2191 (.A1(W1275), .A2(W19645), .ZN(W37650));
  NOR2X1 G2192 (.A1(W27496), .A2(W16151), .ZN(O5051));
  NOR2X1 G2193 (.A1(W6374), .A2(W12593), .ZN(W13174));
  NOR2X1 G2194 (.A1(W2906), .A2(W9128), .ZN(O9101));
  NOR2X1 G2195 (.A1(W5237), .A2(W12260), .ZN(W13141));
  NOR2X1 G2196 (.A1(W5295), .A2(W19719), .ZN(O9104));
  NOR2X1 G2197 (.A1(W12360), .A2(W10113), .ZN(O705));
  NOR2X1 G2198 (.A1(W26363), .A2(W4494), .ZN(W29800));
  NOR2X1 G2199 (.A1(W37518), .A2(W13811), .ZN(W37658));
  NOR2X1 G2200 (.A1(W10811), .A2(W13951), .ZN(O9105));
  NOR2X1 G2201 (.A1(W4286), .A2(W4362), .ZN(W20963));
  NOR2X1 G2202 (.A1(W7870), .A2(W15349), .ZN(O9109));
  NOR2X1 G2203 (.A1(W19116), .A2(I1651), .ZN(W20984));
  NOR2X1 G2204 (.A1(W27480), .A2(W19000), .ZN(W37710));
  NOR2X1 G2205 (.A1(W5201), .A2(W33759), .ZN(O9141));
  NOR2X1 G2206 (.A1(W15482), .A2(W9462), .ZN(O5039));
  NOR2X1 G2207 (.A1(W4192), .A2(W9382), .ZN(O9142));
  NOR2X1 G2208 (.A1(W19708), .A2(I1889), .ZN(O2128));
  NOR2X1 G2209 (.A1(W35133), .A2(W30713), .ZN(W37718));
  NOR2X1 G2210 (.A1(W8408), .A2(W12794), .ZN(W13114));
  NOR2X1 G2211 (.A1(W21010), .A2(W31041), .ZN(O9147));
  NOR2X1 G2212 (.A1(W27652), .A2(W8583), .ZN(W37709));
  NOR2X1 G2213 (.A1(W15217), .A2(W25162), .ZN(W29780));
  NOR2X1 G2214 (.A1(W9906), .A2(W25032), .ZN(W29779));
  NOR2X1 G2215 (.A1(W7167), .A2(W3535), .ZN(W13108));
  NOR2X1 G2216 (.A1(W11571), .A2(W27356), .ZN(O9151));
  NOR2X1 G2217 (.A1(W7091), .A2(W4648), .ZN(O9152));
  NOR2X1 G2218 (.A1(W14053), .A2(W10930), .ZN(O9153));
  NOR2X1 G2219 (.A1(W23129), .A2(W11246), .ZN(W29778));
  NOR2X1 G2220 (.A1(W5941), .A2(W22781), .ZN(W29790));
  NOR2X1 G2221 (.A1(W25803), .A2(W26587), .ZN(O9132));
  NOR2X1 G2222 (.A1(W37059), .A2(W3250), .ZN(W37692));
  NOR2X1 G2223 (.A1(W7829), .A2(W23006), .ZN(O5044));
  NOR2X1 G2224 (.A1(W17245), .A2(W6935), .ZN(W37695));
  NOR2X1 G2225 (.A1(I1851), .A2(W2164), .ZN(W13136));
  NOR2X1 G2226 (.A1(W4129), .A2(W4449), .ZN(W13135));
  NOR2X1 G2227 (.A1(I1865), .A2(W836), .ZN(W13134));
  NOR2X1 G2228 (.A1(W9736), .A2(I554), .ZN(O5043));
  NOR2X1 G2229 (.A1(W27541), .A2(W16041), .ZN(O10168));
  NOR2X1 G2230 (.A1(W2831), .A2(W5060), .ZN(W13131));
  NOR2X1 G2231 (.A1(W19090), .A2(I1815), .ZN(W29789));
  NOR2X1 G2232 (.A1(W13713), .A2(W30700), .ZN(O9137));
  NOR2X1 G2233 (.A1(W6148), .A2(W20098), .ZN(W20976));
  NOR2X1 G2234 (.A1(W1045), .A2(W11599), .ZN(W13127));
  NOR2X1 G2235 (.A1(W6859), .A2(W8942), .ZN(O2125));
  NOR2X1 G2236 (.A1(W9517), .A2(I1445), .ZN(W13123));
  NOR2X1 G2237 (.A1(W8743), .A2(I1284), .ZN(W9802));
  NOR2X1 G2238 (.A1(W3106), .A2(W2872), .ZN(W9810));
  NOR2X1 G2239 (.A1(W6007), .A2(W8720), .ZN(W9809));
  NOR2X1 G2240 (.A1(W8605), .A2(I518), .ZN(W9808));
  NOR2X1 G2241 (.A1(W5188), .A2(W33323), .ZN(O11364));
  NOR2X1 G2242 (.A1(W7672), .A2(W7148), .ZN(W28729));
  NOR2X1 G2243 (.A1(W12413), .A2(W15951), .ZN(O11367));
  NOR2X1 G2244 (.A1(W4522), .A2(I354), .ZN(O329));
  NOR2X1 G2245 (.A1(W5344), .A2(W1469), .ZN(W9803));
  NOR2X1 G2246 (.A1(W9147), .A2(W33080), .ZN(O11362));
  NOR2X1 G2247 (.A1(W34444), .A2(W3146), .ZN(O11369));
  NOR2X1 G2248 (.A1(W20013), .A2(W25498), .ZN(O11370));
  NOR2X1 G2249 (.A1(W11276), .A2(I1122), .ZN(O11372));
  NOR2X1 G2250 (.A1(W17905), .A2(W12009), .ZN(W22051));
  NOR2X1 G2251 (.A1(W7336), .A2(W8930), .ZN(W9797));
  NOR2X1 G2252 (.A1(W4637), .A2(W8457), .ZN(W9796));
  NOR2X1 G2253 (.A1(W25460), .A2(W26827), .ZN(O11377));
  NOR2X1 G2254 (.A1(W194), .A2(W3028), .ZN(O326));
  NOR2X1 G2255 (.A1(W13206), .A2(W7542), .ZN(W41079));
  NOR2X1 G2256 (.A1(W9656), .A2(I1202), .ZN(O331));
  NOR2X1 G2257 (.A1(W159), .A2(I693), .ZN(W28733));
  NOR2X1 G2258 (.A1(W27438), .A2(W27278), .ZN(W41072));
  NOR2X1 G2259 (.A1(W6926), .A2(W1873), .ZN(O330));
  NOR2X1 G2260 (.A1(W37723), .A2(W26451), .ZN(O11345));
  NOR2X1 G2261 (.A1(I185), .A2(W8677), .ZN(W9822));
  NOR2X1 G2262 (.A1(W37618), .A2(W31668), .ZN(O11348));
  NOR2X1 G2263 (.A1(W6652), .A2(W37063), .ZN(O11349));
  NOR2X1 G2264 (.A1(W3135), .A2(W5639), .ZN(W41114));
  NOR2X1 G2265 (.A1(W430), .A2(W4119), .ZN(W9818));
  NOR2X1 G2266 (.A1(W823), .A2(W688), .ZN(W9817));
  NOR2X1 G2267 (.A1(W4982), .A2(W40038), .ZN(O11350));
  NOR2X1 G2268 (.A1(W32660), .A2(W13294), .ZN(O11354));
  NOR2X1 G2269 (.A1(W9533), .A2(W537), .ZN(W9814));
  NOR2X1 G2270 (.A1(I641), .A2(W4785), .ZN(W9813));
  NOR2X1 G2271 (.A1(W23781), .A2(W16187), .ZN(O11360));
  NOR2X1 G2272 (.A1(W24616), .A2(W37969), .ZN(O11401));
  NOR2X1 G2273 (.A1(W36903), .A2(I1979), .ZN(O11393));
  NOR2X1 G2274 (.A1(W17690), .A2(I422), .ZN(W41134));
  NOR2X1 G2275 (.A1(W17742), .A2(W39686), .ZN(O11394));
  NOR2X1 G2276 (.A1(W3476), .A2(W2984), .ZN(W9770));
  NOR2X1 G2277 (.A1(W3078), .A2(W8547), .ZN(W9769));
  NOR2X1 G2278 (.A1(W14423), .A2(W21027), .ZN(O11398));
  NOR2X1 G2279 (.A1(W22300), .A2(W12556), .ZN(O11399));
  NOR2X1 G2280 (.A1(W12232), .A2(W13607), .ZN(W22057));
  NOR2X1 G2281 (.A1(W31235), .A2(W9042), .ZN(O11391));
  NOR2X1 G2282 (.A1(W23831), .A2(W11285), .ZN(O11402));
  NOR2X1 G2283 (.A1(W38504), .A2(W28651), .ZN(O11403));
  NOR2X1 G2284 (.A1(I422), .A2(W3898), .ZN(W9762));
  NOR2X1 G2285 (.A1(W38148), .A2(W5294), .ZN(W41149));
  NOR2X1 G2286 (.A1(W39285), .A2(W16866), .ZN(O11408));
  NOR2X1 G2287 (.A1(W24464), .A2(W30414), .ZN(W41154));
  NOR2X1 G2288 (.A1(W20592), .A2(W17153), .ZN(O2414));
  NOR2X1 G2289 (.A1(W8035), .A2(W660), .ZN(W9757));
  NOR2X1 G2290 (.A1(W2949), .A2(W31344), .ZN(O11388));
  NOR2X1 G2291 (.A1(I630), .A2(W23559), .ZN(W41117));
  NOR2X1 G2292 (.A1(W30050), .A2(W40286), .ZN(O11382));
  NOR2X1 G2293 (.A1(W5724), .A2(W7593), .ZN(W9789));
  NOR2X1 G2294 (.A1(W401), .A2(W2957), .ZN(W9788));
  NOR2X1 G2295 (.A1(W11800), .A2(W28358), .ZN(O4590));
  NOR2X1 G2296 (.A1(W26048), .A2(W36760), .ZN(O11386));
  NOR2X1 G2297 (.A1(W11206), .A2(W2854), .ZN(O11387));
  NOR2X1 G2298 (.A1(W38555), .A2(W22369), .ZN(W41125));
  NOR2X1 G2299 (.A1(W24752), .A2(W16491), .ZN(O11344));
  NOR2X1 G2300 (.A1(W11586), .A2(W11224), .ZN(O2412));
  NOR2X1 G2301 (.A1(W159), .A2(I556), .ZN(W9781));
  NOR2X1 G2302 (.A1(W7061), .A2(W725), .ZN(W9779));
  NOR2X1 G2303 (.A1(W8951), .A2(W8741), .ZN(W9778));
  NOR2X1 G2304 (.A1(W3894), .A2(I1033), .ZN(W9777));
  NOR2X1 G2305 (.A1(W8292), .A2(W309), .ZN(W9776));
  NOR2X1 G2306 (.A1(W21712), .A2(W6998), .ZN(O4589));
  NOR2X1 G2307 (.A1(W4185), .A2(W17664), .ZN(O11317));
  NOR2X1 G2308 (.A1(I1123), .A2(W3700), .ZN(W9885));
  NOR2X1 G2309 (.A1(W21735), .A2(W1910), .ZN(W41026));
  NOR2X1 G2310 (.A1(W27809), .A2(W25006), .ZN(W28750));
  NOR2X1 G2311 (.A1(I431), .A2(W38787), .ZN(O11315));
  NOR2X1 G2312 (.A1(W7889), .A2(W1608), .ZN(W9881));
  NOR2X1 G2313 (.A1(W9132), .A2(W2316), .ZN(W9880));
  NOR2X1 G2314 (.A1(I1391), .A2(W8407), .ZN(W9878));
  NOR2X1 G2315 (.A1(W18973), .A2(W16705), .ZN(W22034));
  NOR2X1 G2316 (.A1(W3614), .A2(W2406), .ZN(W9886));
  NOR2X1 G2317 (.A1(W15671), .A2(W5425), .ZN(W28747));
  NOR2X1 G2318 (.A1(W32420), .A2(W37313), .ZN(W41038));
  NOR2X1 G2319 (.A1(W9411), .A2(W614), .ZN(W9873));
  NOR2X1 G2320 (.A1(W32260), .A2(W31524), .ZN(O11320));
  NOR2X1 G2321 (.A1(W36042), .A2(W31078), .ZN(W41040));
  NOR2X1 G2322 (.A1(W21710), .A2(W9070), .ZN(W22036));
  NOR2X1 G2323 (.A1(W16380), .A2(W14665), .ZN(W22037));
  NOR2X1 G2324 (.A1(W9319), .A2(W5414), .ZN(W9868));
  NOR2X1 G2325 (.A1(W3393), .A2(W18208), .ZN(O2407));
  NOR2X1 G2326 (.A1(W6391), .A2(W9624), .ZN(O4604));
  NOR2X1 G2327 (.A1(W12019), .A2(W33900), .ZN(O11304));
  NOR2X1 G2328 (.A1(W100), .A2(W8526), .ZN(W9901));
  NOR2X1 G2329 (.A1(W21974), .A2(W38033), .ZN(W41012));
  NOR2X1 G2330 (.A1(W8925), .A2(W3921), .ZN(W9899));
  NOR2X1 G2331 (.A1(W5369), .A2(W21801), .ZN(W28753));
  NOR2X1 G2332 (.A1(W28677), .A2(W37001), .ZN(O11306));
  NOR2X1 G2333 (.A1(W5425), .A2(W7005), .ZN(W9896));
  NOR2X1 G2334 (.A1(W19164), .A2(W406), .ZN(W22038));
  NOR2X1 G2335 (.A1(W8816), .A2(W6063), .ZN(W9893));
  NOR2X1 G2336 (.A1(W39893), .A2(W11679), .ZN(O11309));
  NOR2X1 G2337 (.A1(W555), .A2(W5824), .ZN(W9891));
  NOR2X1 G2338 (.A1(W23718), .A2(I455), .ZN(O11310));
  NOR2X1 G2339 (.A1(W8957), .A2(W1930), .ZN(W41022));
  NOR2X1 G2340 (.A1(W19052), .A2(W11992), .ZN(O2408));
  NOR2X1 G2341 (.A1(W3984), .A2(W9485), .ZN(W9887));
  NOR2X1 G2342 (.A1(W9666), .A2(W3464), .ZN(W9838));
  NOR2X1 G2343 (.A1(W22849), .A2(W12152), .ZN(W41054));
  NOR2X1 G2344 (.A1(W1064), .A2(W8653), .ZN(W9846));
  NOR2X1 G2345 (.A1(W18288), .A2(W11165), .ZN(O4601));
  NOR2X1 G2346 (.A1(W31612), .A2(W19807), .ZN(W41056));
  NOR2X1 G2347 (.A1(W6611), .A2(W3907), .ZN(W9843));
  NOR2X1 G2348 (.A1(I247), .A2(W6062), .ZN(W9842));
  NOR2X1 G2349 (.A1(W3362), .A2(W3806), .ZN(W9841));
  NOR2X1 G2350 (.A1(W6394), .A2(I1734), .ZN(W9840));
  NOR2X1 G2351 (.A1(W34779), .A2(W3352), .ZN(W41053));
  NOR2X1 G2352 (.A1(I1938), .A2(W2866), .ZN(W9837));
  NOR2X1 G2353 (.A1(W8597), .A2(W11211), .ZN(W28735));
  NOR2X1 G2354 (.A1(W10253), .A2(W3310), .ZN(O2410));
  NOR2X1 G2355 (.A1(W10325), .A2(W9174), .ZN(W41064));
  NOR2X1 G2356 (.A1(W35230), .A2(W7299), .ZN(O11340));
  NOR2X1 G2357 (.A1(W27969), .A2(W34560), .ZN(O11342));
  NOR2X1 G2358 (.A1(W6431), .A2(W9496), .ZN(W22047));
  NOR2X1 G2359 (.A1(W8866), .A2(W9459), .ZN(W9830));
  NOR2X1 G2360 (.A1(W972), .A2(W7387), .ZN(W9856));
  NOR2X1 G2361 (.A1(W2370), .A2(W3625), .ZN(W9866));
  NOR2X1 G2362 (.A1(I518), .A2(W3336), .ZN(W9865));
  NOR2X1 G2363 (.A1(W6367), .A2(W5055), .ZN(W9863));
  NOR2X1 G2364 (.A1(W4461), .A2(I1719), .ZN(W9862));
  NOR2X1 G2365 (.A1(W5093), .A2(W4865), .ZN(O332));
  NOR2X1 G2366 (.A1(W9217), .A2(W3891), .ZN(W9860));
  NOR2X1 G2367 (.A1(W18235), .A2(W5141), .ZN(W22040));
  NOR2X1 G2368 (.A1(W27032), .A2(W23925), .ZN(O11328));
  NOR2X1 G2369 (.A1(W1967), .A2(W40776), .ZN(O11411));
  NOR2X1 G2370 (.A1(W5771), .A2(W4269), .ZN(W9855));
  NOR2X1 G2371 (.A1(W7010), .A2(W1564), .ZN(W9854));
  NOR2X1 G2372 (.A1(W20736), .A2(W962), .ZN(W22042));
  NOR2X1 G2373 (.A1(W8809), .A2(I1276), .ZN(W9852));
  NOR2X1 G2374 (.A1(W23809), .A2(W2117), .ZN(O11330));
  NOR2X1 G2375 (.A1(W39616), .A2(I821), .ZN(O11331));
  NOR2X1 G2376 (.A1(W33314), .A2(I130), .ZN(O11332));
  NOR2X1 G2377 (.A1(W3588), .A2(W6516), .ZN(W9643));
  NOR2X1 G2378 (.A1(W10270), .A2(W35367), .ZN(O11478));
  NOR2X1 G2379 (.A1(W7889), .A2(W38381), .ZN(O11479));
  NOR2X1 G2380 (.A1(W6540), .A2(W7540), .ZN(O311));
  NOR2X1 G2381 (.A1(W22482), .A2(I233), .ZN(W41266));
  NOR2X1 G2382 (.A1(W30315), .A2(W18921), .ZN(O11480));
  NOR2X1 G2383 (.A1(W19403), .A2(W6885), .ZN(W28677));
  NOR2X1 G2384 (.A1(W5555), .A2(I1069), .ZN(W9645));
  NOR2X1 G2385 (.A1(W21216), .A2(W14731), .ZN(W22095));
  NOR2X1 G2386 (.A1(W2328), .A2(W4935), .ZN(W9653));
  NOR2X1 G2387 (.A1(W4947), .A2(W8365), .ZN(O309));
  NOR2X1 G2388 (.A1(W14488), .A2(W6218), .ZN(O11483));
  NOR2X1 G2389 (.A1(W4458), .A2(W6238), .ZN(W9640));
  NOR2X1 G2390 (.A1(W21014), .A2(W2521), .ZN(O11485));
  NOR2X1 G2391 (.A1(W8145), .A2(I1271), .ZN(W9638));
  NOR2X1 G2392 (.A1(W28644), .A2(W16571), .ZN(O11486));
  NOR2X1 G2393 (.A1(W6), .A2(W9103), .ZN(W9635));
  NOR2X1 G2394 (.A1(W9435), .A2(I996), .ZN(O308));
  NOR2X1 G2395 (.A1(W27927), .A2(W14285), .ZN(O11474));
  NOR2X1 G2396 (.A1(W18027), .A2(W3548), .ZN(W22087));
  NOR2X1 G2397 (.A1(W1124), .A2(W9501), .ZN(W9672));
  NOR2X1 G2398 (.A1(W3543), .A2(W8616), .ZN(W9670));
  NOR2X1 G2399 (.A1(I919), .A2(W29578), .ZN(O11469));
  NOR2X1 G2400 (.A1(I1526), .A2(W4309), .ZN(W9667));
  NOR2X1 G2401 (.A1(W40604), .A2(W3734), .ZN(O11471));
  NOR2X1 G2402 (.A1(W24452), .A2(W9688), .ZN(W28680));
  NOR2X1 G2403 (.A1(W33726), .A2(W3345), .ZN(O11473));
  NOR2X1 G2404 (.A1(W7316), .A2(W1784), .ZN(W9633));
  NOR2X1 G2405 (.A1(I716), .A2(W857), .ZN(W9661));
  NOR2X1 G2406 (.A1(W6962), .A2(W1807), .ZN(W9660));
  NOR2X1 G2407 (.A1(W10435), .A2(W12406), .ZN(W41258));
  NOR2X1 G2408 (.A1(W14497), .A2(W22794), .ZN(W41261));
  NOR2X1 G2409 (.A1(W7120), .A2(W6377), .ZN(W9656));
  NOR2X1 G2410 (.A1(W14522), .A2(W37488), .ZN(O11477));
  NOR2X1 G2411 (.A1(W1819), .A2(W1117), .ZN(W9654));
  NOR2X1 G2412 (.A1(W11173), .A2(W10974), .ZN(W28664));
  NOR2X1 G2413 (.A1(W1698), .A2(W6508), .ZN(W9611));
  NOR2X1 G2414 (.A1(W7800), .A2(W1130), .ZN(W9609));
  NOR2X1 G2415 (.A1(W7528), .A2(W9535), .ZN(W9608));
  NOR2X1 G2416 (.A1(I948), .A2(W30971), .ZN(O11503));
  NOR2X1 G2417 (.A1(W15956), .A2(W36810), .ZN(O11508));
  NOR2X1 G2418 (.A1(W32810), .A2(W27075), .ZN(O11509));
  NOR2X1 G2419 (.A1(W8665), .A2(W1998), .ZN(O305));
  NOR2X1 G2420 (.A1(W9587), .A2(W11187), .ZN(W28665));
  NOR2X1 G2421 (.A1(W18393), .A2(W6885), .ZN(W28669));
  NOR2X1 G2422 (.A1(W39552), .A2(W27738), .ZN(O11517));
  NOR2X1 G2423 (.A1(W12853), .A2(W18199), .ZN(W22112));
  NOR2X1 G2424 (.A1(W27007), .A2(W24396), .ZN(O4571));
  NOR2X1 G2425 (.A1(W6556), .A2(W8179), .ZN(W9592));
  NOR2X1 G2426 (.A1(W28081), .A2(W7011), .ZN(O11525));
  NOR2X1 G2427 (.A1(W26701), .A2(W28180), .ZN(O11528));
  NOR2X1 G2428 (.A1(W28504), .A2(W40211), .ZN(O11529));
  NOR2X1 G2429 (.A1(W6075), .A2(W9077), .ZN(W9586));
  NOR2X1 G2430 (.A1(I1392), .A2(W8601), .ZN(W9624));
  NOR2X1 G2431 (.A1(W31345), .A2(W32396), .ZN(O11487));
  NOR2X1 G2432 (.A1(W38952), .A2(W10284), .ZN(W41280));
  NOR2X1 G2433 (.A1(I1043), .A2(W15959), .ZN(W22097));
  NOR2X1 G2434 (.A1(W6001), .A2(W25851), .ZN(O11488));
  NOR2X1 G2435 (.A1(I1088), .A2(W39983), .ZN(O11489));
  NOR2X1 G2436 (.A1(W23667), .A2(W16827), .ZN(O11490));
  NOR2X1 G2437 (.A1(W19558), .A2(W35220), .ZN(W41287));
  NOR2X1 G2438 (.A1(W41071), .A2(W37709), .ZN(W41288));
  NOR2X1 G2439 (.A1(W38469), .A2(W7203), .ZN(O11466));
  NOR2X1 G2440 (.A1(W1958), .A2(W16270), .ZN(W41290));
  NOR2X1 G2441 (.A1(W9413), .A2(W2417), .ZN(W9621));
  NOR2X1 G2442 (.A1(W7418), .A2(I1568), .ZN(W22100));
  NOR2X1 G2443 (.A1(W23735), .A2(W15524), .ZN(W41293));
  NOR2X1 G2444 (.A1(W22246), .A2(W35631), .ZN(W41294));
  NOR2X1 G2445 (.A1(I1931), .A2(W7244), .ZN(W9615));
  NOR2X1 G2446 (.A1(W26091), .A2(W12864), .ZN(O11497));
  NOR2X1 G2447 (.A1(W2355), .A2(W949), .ZN(W9719));
  NOR2X1 G2448 (.A1(W3779), .A2(W3310), .ZN(W22072));
  NOR2X1 G2449 (.A1(W4442), .A2(W7614), .ZN(O320));
  NOR2X1 G2450 (.A1(W22821), .A2(W11991), .ZN(O4584));
  NOR2X1 G2451 (.A1(W3102), .A2(W23963), .ZN(O11436));
  NOR2X1 G2452 (.A1(W5400), .A2(W8341), .ZN(W9725));
  NOR2X1 G2453 (.A1(W7198), .A2(W2613), .ZN(W9724));
  NOR2X1 G2454 (.A1(W1251), .A2(I212), .ZN(O319));
  NOR2X1 G2455 (.A1(W28043), .A2(W12424), .ZN(W41203));
  NOR2X1 G2456 (.A1(W26766), .A2(W36977), .ZN(W41192));
  NOR2X1 G2457 (.A1(I164), .A2(W9169), .ZN(W9718));
  NOR2X1 G2458 (.A1(W4908), .A2(W11283), .ZN(W22077));
  NOR2X1 G2459 (.A1(I790), .A2(W11706), .ZN(W41207));
  NOR2X1 G2460 (.A1(W2279), .A2(W29938), .ZN(W41209));
  NOR2X1 G2461 (.A1(W5697), .A2(W3228), .ZN(W9714));
  NOR2X1 G2462 (.A1(W26474), .A2(W34269), .ZN(O11444));
  NOR2X1 G2463 (.A1(W6429), .A2(W8525), .ZN(W9712));
  NOR2X1 G2464 (.A1(W4886), .A2(W7852), .ZN(W28692));
  NOR2X1 G2465 (.A1(W18516), .A2(W10391), .ZN(W22064));
  NOR2X1 G2466 (.A1(W6239), .A2(W9423), .ZN(W9755));
  NOR2X1 G2467 (.A1(W4059), .A2(W6570), .ZN(W9754));
  NOR2X1 G2468 (.A1(I55), .A2(W9574), .ZN(W9753));
  NOR2X1 G2469 (.A1(W7408), .A2(W19008), .ZN(O11415));
  NOR2X1 G2470 (.A1(W7303), .A2(W13953), .ZN(O11420));
  NOR2X1 G2471 (.A1(W8783), .A2(W5498), .ZN(W9746));
  NOR2X1 G2472 (.A1(W8323), .A2(W906), .ZN(W9745));
  NOR2X1 G2473 (.A1(W18930), .A2(W20581), .ZN(O4586));
  NOR2X1 G2474 (.A1(W15859), .A2(W16029), .ZN(W41216));
  NOR2X1 G2475 (.A1(W910), .A2(W8691), .ZN(O2418));
  NOR2X1 G2476 (.A1(W11485), .A2(W17777), .ZN(W22069));
  NOR2X1 G2477 (.A1(W20632), .A2(W32673), .ZN(O11429));
  NOR2X1 G2478 (.A1(W27564), .A2(W19374), .ZN(O11431));
  NOR2X1 G2479 (.A1(W6071), .A2(W10042), .ZN(O11432));
  NOR2X1 G2480 (.A1(W19902), .A2(W11494), .ZN(O4585));
  NOR2X1 G2481 (.A1(W5576), .A2(W5108), .ZN(W9732));
  NOR2X1 G2482 (.A1(W12788), .A2(W20733), .ZN(W28687));
  NOR2X1 G2483 (.A1(W2767), .A2(W4129), .ZN(W9691));
  NOR2X1 G2484 (.A1(W17261), .A2(W5925), .ZN(W28689));
  NOR2X1 G2485 (.A1(W4117), .A2(W4664), .ZN(W9689));
  NOR2X1 G2486 (.A1(W5648), .A2(W4042), .ZN(W9688));
  NOR2X1 G2487 (.A1(W4159), .A2(I234), .ZN(W9687));
  NOR2X1 G2488 (.A1(W5031), .A2(W19571), .ZN(W22084));
  NOR2X1 G2489 (.A1(W8145), .A2(W6500), .ZN(W9685));
  NOR2X1 G2490 (.A1(W29955), .A2(W14120), .ZN(W41235));
  NOR2X1 G2491 (.A1(W16472), .A2(W31863), .ZN(O11458));
  NOR2X1 G2492 (.A1(W21039), .A2(W35976), .ZN(O11461));
  NOR2X1 G2493 (.A1(W22457), .A2(W9726), .ZN(W28686));
  NOR2X1 G2494 (.A1(I1697), .A2(W7463), .ZN(W9680));
  NOR2X1 G2495 (.A1(W3647), .A2(W3007), .ZN(W9679));
  NOR2X1 G2496 (.A1(I1974), .A2(W6519), .ZN(W9678));
  NOR2X1 G2497 (.A1(W32388), .A2(W17145), .ZN(O11464));
  NOR2X1 G2498 (.A1(W23519), .A2(W11500), .ZN(O11465));
  NOR2X1 G2499 (.A1(W4641), .A2(W235), .ZN(W9675));
  NOR2X1 G2500 (.A1(W21340), .A2(W1598), .ZN(W22081));
  NOR2X1 G2501 (.A1(W9627), .A2(W4505), .ZN(W9708));
  NOR2X1 G2502 (.A1(W5335), .A2(W22390), .ZN(O11448));
  NOR2X1 G2503 (.A1(W689), .A2(I1872), .ZN(W9706));
  NOR2X1 G2504 (.A1(I647), .A2(W7079), .ZN(W9705));
  NOR2X1 G2505 (.A1(I1542), .A2(W17993), .ZN(O11449));
  NOR2X1 G2506 (.A1(W14512), .A2(W24252), .ZN(W41219));
  NOR2X1 G2507 (.A1(W5386), .A2(W27287), .ZN(W28691));
  NOR2X1 G2508 (.A1(W3202), .A2(W5943), .ZN(W9701));
  NOR2X1 G2509 (.A1(I967), .A2(W5352), .ZN(W9904));
  NOR2X1 G2510 (.A1(W17289), .A2(W9203), .ZN(O11452));
  NOR2X1 G2511 (.A1(W7447), .A2(W1788), .ZN(W9698));
  NOR2X1 G2512 (.A1(W28828), .A2(W3262), .ZN(O11453));
  NOR2X1 G2513 (.A1(W1814), .A2(W4993), .ZN(W9696));
  NOR2X1 G2514 (.A1(W8499), .A2(W6731), .ZN(W9695));
  NOR2X1 G2515 (.A1(W27630), .A2(W3911), .ZN(O11454));
  NOR2X1 G2516 (.A1(W3131), .A2(W5889), .ZN(W22082));
  NOR2X1 G2517 (.A1(W25251), .A2(W2044), .ZN(O11141));
  NOR2X1 G2518 (.A1(W35468), .A2(W18578), .ZN(W40771));
  NOR2X1 G2519 (.A1(W28092), .A2(W26263), .ZN(O11138));
  NOR2X1 G2520 (.A1(I1079), .A2(I1640), .ZN(W10112));
  NOR2X1 G2521 (.A1(W11841), .A2(W5149), .ZN(W28823));
  NOR2X1 G2522 (.A1(W1167), .A2(W8263), .ZN(W10110));
  NOR2X1 G2523 (.A1(W3095), .A2(W18268), .ZN(W21959));
  NOR2X1 G2524 (.A1(W899), .A2(W6158), .ZN(W10107));
  NOR2X1 G2525 (.A1(W9341), .A2(W7321), .ZN(W10106));
  NOR2X1 G2526 (.A1(W3761), .A2(W9460), .ZN(W10115));
  NOR2X1 G2527 (.A1(W20174), .A2(W9892), .ZN(W28821));
  NOR2X1 G2528 (.A1(W1267), .A2(W3875), .ZN(W10103));
  NOR2X1 G2529 (.A1(W9721), .A2(W2217), .ZN(W10102));
  NOR2X1 G2530 (.A1(W37785), .A2(W8468), .ZN(O11143));
  NOR2X1 G2531 (.A1(W30227), .A2(W37863), .ZN(W40781));
  NOR2X1 G2532 (.A1(W14702), .A2(W37712), .ZN(O11144));
  NOR2X1 G2533 (.A1(W18491), .A2(I1654), .ZN(W21961));
  NOR2X1 G2534 (.A1(W9065), .A2(W6311), .ZN(O11145));
  NOR2X1 G2535 (.A1(W19957), .A2(W10543), .ZN(O2384));
  NOR2X1 G2536 (.A1(W22183), .A2(W33175), .ZN(W40757));
  NOR2X1 G2537 (.A1(W6284), .A2(W750), .ZN(W21952));
  NOR2X1 G2538 (.A1(W3907), .A2(W855), .ZN(W10130));
  NOR2X1 G2539 (.A1(W6750), .A2(W5252), .ZN(W10129));
  NOR2X1 G2540 (.A1(W10580), .A2(W35131), .ZN(O11128));
  NOR2X1 G2541 (.A1(W24209), .A2(W879), .ZN(O4630));
  NOR2X1 G2542 (.A1(W7337), .A2(W24058), .ZN(W28825));
  NOR2X1 G2543 (.A1(W5038), .A2(W7868), .ZN(W10125));
  NOR2X1 G2544 (.A1(W9908), .A2(W39978), .ZN(O11146));
  NOR2X1 G2545 (.A1(I1557), .A2(W5572), .ZN(W10122));
  NOR2X1 G2546 (.A1(W8811), .A2(W4489), .ZN(W10121));
  NOR2X1 G2547 (.A1(W140), .A2(W8547), .ZN(O363));
  NOR2X1 G2548 (.A1(W8190), .A2(W2446), .ZN(W10119));
  NOR2X1 G2549 (.A1(W14138), .A2(W4854), .ZN(O11132));
  NOR2X1 G2550 (.A1(W5212), .A2(W7992), .ZN(O11134));
  NOR2X1 G2551 (.A1(W2649), .A2(W20200), .ZN(O11135));
  NOR2X1 G2552 (.A1(W4608), .A2(W7291), .ZN(W10068));
  NOR2X1 G2553 (.A1(W20297), .A2(W33538), .ZN(O11160));
  NOR2X1 G2554 (.A1(W35871), .A2(W24446), .ZN(O11161));
  NOR2X1 G2555 (.A1(W91), .A2(W8587), .ZN(W10075));
  NOR2X1 G2556 (.A1(W4888), .A2(W4230), .ZN(W28816));
  NOR2X1 G2557 (.A1(W976), .A2(W1509), .ZN(W10073));
  NOR2X1 G2558 (.A1(W3567), .A2(W9775), .ZN(O360));
  NOR2X1 G2559 (.A1(W25185), .A2(W2019), .ZN(W40813));
  NOR2X1 G2560 (.A1(W2929), .A2(W10018), .ZN(W10070));
  NOR2X1 G2561 (.A1(W34496), .A2(W36411), .ZN(O11159));
  NOR2X1 G2562 (.A1(W15218), .A2(W9623), .ZN(W40815));
  NOR2X1 G2563 (.A1(W4024), .A2(W3316), .ZN(O358));
  NOR2X1 G2564 (.A1(W5807), .A2(W14593), .ZN(W40816));
  NOR2X1 G2565 (.A1(W7194), .A2(I45), .ZN(W10064));
  NOR2X1 G2566 (.A1(W6087), .A2(W16294), .ZN(O2389));
  NOR2X1 G2567 (.A1(W733), .A2(W4532), .ZN(O4626));
  NOR2X1 G2568 (.A1(W7877), .A2(W10020), .ZN(W10061));
  NOR2X1 G2569 (.A1(W371), .A2(W7545), .ZN(W10059));
  NOR2X1 G2570 (.A1(W13403), .A2(W17244), .ZN(W21964));
  NOR2X1 G2571 (.A1(W11325), .A2(W4822), .ZN(W28820));
  NOR2X1 G2572 (.A1(W4600), .A2(W3711), .ZN(W10094));
  NOR2X1 G2573 (.A1(W16878), .A2(W24913), .ZN(O11148));
  NOR2X1 G2574 (.A1(W2533), .A2(W23276), .ZN(W40792));
  NOR2X1 G2575 (.A1(W987), .A2(W26947), .ZN(O4628));
  NOR2X1 G2576 (.A1(W30566), .A2(W31592), .ZN(O11150));
  NOR2X1 G2577 (.A1(W5293), .A2(W7983), .ZN(W10089));
  NOR2X1 G2578 (.A1(W6992), .A2(W6592), .ZN(W10088));
  NOR2X1 G2579 (.A1(W28933), .A2(W14809), .ZN(O11126));
  NOR2X1 G2580 (.A1(W3450), .A2(W1807), .ZN(W10085));
  NOR2X1 G2581 (.A1(W35469), .A2(W19697), .ZN(W40798));
  NOR2X1 G2582 (.A1(W9855), .A2(I1148), .ZN(W10083));
  NOR2X1 G2583 (.A1(W3792), .A2(W17800), .ZN(O2388));
  NOR2X1 G2584 (.A1(W7102), .A2(W8579), .ZN(W10081));
  NOR2X1 G2585 (.A1(W40249), .A2(W18158), .ZN(O11154));
  NOR2X1 G2586 (.A1(W23834), .A2(W3659), .ZN(O11157));
  NOR2X1 G2587 (.A1(W8805), .A2(W22390), .ZN(O4633));
  NOR2X1 G2588 (.A1(W6865), .A2(W2824), .ZN(W10192));
  NOR2X1 G2589 (.A1(W6232), .A2(I1439), .ZN(W10190));
  NOR2X1 G2590 (.A1(W4524), .A2(W10403), .ZN(W21932));
  NOR2X1 G2591 (.A1(W37767), .A2(W7482), .ZN(W40688));
  NOR2X1 G2592 (.A1(W7456), .A2(W4825), .ZN(O2377));
  NOR2X1 G2593 (.A1(W510), .A2(W10106), .ZN(W10186));
  NOR2X1 G2594 (.A1(W32055), .A2(W13722), .ZN(W40693));
  NOR2X1 G2595 (.A1(W35875), .A2(W23339), .ZN(W40695));
  NOR2X1 G2596 (.A1(W27570), .A2(W7787), .ZN(W40684));
  NOR2X1 G2597 (.A1(W6146), .A2(W26267), .ZN(O11081));
  NOR2X1 G2598 (.A1(W8557), .A2(W11184), .ZN(O4632));
  NOR2X1 G2599 (.A1(W9666), .A2(W20500), .ZN(O11085));
  NOR2X1 G2600 (.A1(I595), .A2(W632), .ZN(O11086));
  NOR2X1 G2601 (.A1(W36737), .A2(W21598), .ZN(O11088));
  NOR2X1 G2602 (.A1(W40124), .A2(W33309), .ZN(O11089));
  NOR2X1 G2603 (.A1(W24118), .A2(W2692), .ZN(O11090));
  NOR2X1 G2604 (.A1(W6703), .A2(W2323), .ZN(W10174));
  NOR2X1 G2605 (.A1(W9879), .A2(W28243), .ZN(W28852));
  NOR2X1 G2606 (.A1(W6928), .A2(W9846), .ZN(W10215));
  NOR2X1 G2607 (.A1(W368), .A2(W7757), .ZN(W21922));
  NOR2X1 G2608 (.A1(W1814), .A2(I692), .ZN(W10213));
  NOR2X1 G2609 (.A1(W14227), .A2(W21297), .ZN(O4639));
  NOR2X1 G2610 (.A1(W37413), .A2(I999), .ZN(O11065));
  NOR2X1 G2611 (.A1(W6329), .A2(W1874), .ZN(W40669));
  NOR2X1 G2612 (.A1(W953), .A2(W5519), .ZN(W10208));
  NOR2X1 G2613 (.A1(W37938), .A2(W38944), .ZN(O11067));
  NOR2X1 G2614 (.A1(W23649), .A2(W11643), .ZN(O11091));
  NOR2X1 G2615 (.A1(W27577), .A2(W38839), .ZN(O11069));
  NOR2X1 G2616 (.A1(W9617), .A2(W1126), .ZN(W10202));
  NOR2X1 G2617 (.A1(W4512), .A2(W252), .ZN(W10200));
  NOR2X1 G2618 (.A1(W6638), .A2(W824), .ZN(W40681));
  NOR2X1 G2619 (.A1(W9097), .A2(W15686), .ZN(O11072));
  NOR2X1 G2620 (.A1(W32265), .A2(W2699), .ZN(W40683));
  NOR2X1 G2621 (.A1(W4259), .A2(W10080), .ZN(W10194));
  NOR2X1 G2622 (.A1(W7381), .A2(I2), .ZN(O365));
  NOR2X1 G2623 (.A1(W29027), .A2(W12316), .ZN(O11108));
  NOR2X1 G2624 (.A1(W17470), .A2(W12946), .ZN(W21942));
  NOR2X1 G2625 (.A1(W3767), .A2(W16298), .ZN(W28834));
  NOR2X1 G2626 (.A1(W17846), .A2(I992), .ZN(W21946));
  NOR2X1 G2627 (.A1(W38412), .A2(W39055), .ZN(O11115));
  NOR2X1 G2628 (.A1(I1780), .A2(I1180), .ZN(W10147));
  NOR2X1 G2629 (.A1(W9827), .A2(W6062), .ZN(W10145));
  NOR2X1 G2630 (.A1(W18725), .A2(W12595), .ZN(O11117));
  NOR2X1 G2631 (.A1(W28555), .A2(W22829), .ZN(O11107));
  NOR2X1 G2632 (.A1(W120), .A2(W8370), .ZN(W10142));
  NOR2X1 G2633 (.A1(W30199), .A2(W23675), .ZN(W40747));
  NOR2X1 G2634 (.A1(W18953), .A2(W20480), .ZN(W28832));
  NOR2X1 G2635 (.A1(W6502), .A2(W3050), .ZN(W10139));
  NOR2X1 G2636 (.A1(W18807), .A2(W13857), .ZN(W28831));
  NOR2X1 G2637 (.A1(W24898), .A2(W27824), .ZN(W40752));
  NOR2X1 G2638 (.A1(I850), .A2(W4085), .ZN(W10135));
  NOR2X1 G2639 (.A1(W18199), .A2(W12553), .ZN(W28829));
  NOR2X1 G2640 (.A1(W13581), .A2(W4191), .ZN(W21941));
  NOR2X1 G2641 (.A1(W24572), .A2(W8077), .ZN(O11092));
  NOR2X1 G2642 (.A1(W12881), .A2(W28158), .ZN(W40714));
  NOR2X1 G2643 (.A1(W18099), .A2(W1677), .ZN(W28840));
  NOR2X1 G2644 (.A1(W7425), .A2(W13490), .ZN(W40716));
  NOR2X1 G2645 (.A1(W9938), .A2(W19496), .ZN(W40721));
  NOR2X1 G2646 (.A1(W15992), .A2(W20869), .ZN(O2380));
  NOR2X1 G2647 (.A1(I1440), .A2(W6399), .ZN(W10165));
  NOR2X1 G2648 (.A1(W4412), .A2(W7176), .ZN(W28838));
  NOR2X1 G2649 (.A1(W887), .A2(W1655), .ZN(O11168));
  NOR2X1 G2650 (.A1(I1368), .A2(I1089), .ZN(W10162));
  NOR2X1 G2651 (.A1(W1793), .A2(W3874), .ZN(W10161));
  NOR2X1 G2652 (.A1(W1432), .A2(W10155), .ZN(W10160));
  NOR2X1 G2653 (.A1(W29282), .A2(W34336), .ZN(O11102));
  NOR2X1 G2654 (.A1(W3299), .A2(W29561), .ZN(O11104));
  NOR2X1 G2655 (.A1(I128), .A2(W8580), .ZN(O11105));
  NOR2X1 G2656 (.A1(W327), .A2(W5348), .ZN(W10156));
  NOR2X1 G2657 (.A1(W8478), .A2(W7524), .ZN(W9955));
  NOR2X1 G2658 (.A1(W36718), .A2(W11087), .ZN(O11258));
  NOR2X1 G2659 (.A1(W16841), .A2(W10285), .ZN(W28774));
  NOR2X1 G2660 (.A1(W34821), .A2(I595), .ZN(O11262));
  NOR2X1 G2661 (.A1(W29337), .A2(W6264), .ZN(W40950));
  NOR2X1 G2662 (.A1(W10446), .A2(W656), .ZN(O4612));
  NOR2X1 G2663 (.A1(W6302), .A2(I1793), .ZN(W9959));
  NOR2X1 G2664 (.A1(I1475), .A2(W3766), .ZN(W9957));
  NOR2X1 G2665 (.A1(W39025), .A2(W16764), .ZN(O11265));
  NOR2X1 G2666 (.A1(W16343), .A2(W36718), .ZN(O11256));
  NOR2X1 G2667 (.A1(W33944), .A2(W13820), .ZN(O11266));
  NOR2X1 G2668 (.A1(W1389), .A2(W8986), .ZN(W9953));
  NOR2X1 G2669 (.A1(W9706), .A2(W24376), .ZN(W40957));
  NOR2X1 G2670 (.A1(W8412), .A2(W21558), .ZN(W22013));
  NOR2X1 G2671 (.A1(I977), .A2(W33366), .ZN(O11270));
  NOR2X1 G2672 (.A1(W12114), .A2(W25617), .ZN(O4611));
  NOR2X1 G2673 (.A1(W424), .A2(W2394), .ZN(W9948));
  NOR2X1 G2674 (.A1(W1153), .A2(W6056), .ZN(W9947));
  NOR2X1 G2675 (.A1(I1038), .A2(W18984), .ZN(W28780));
  NOR2X1 G2676 (.A1(W3350), .A2(W16230), .ZN(O2395));
  NOR2X1 G2677 (.A1(W19503), .A2(W20836), .ZN(W28785));
  NOR2X1 G2678 (.A1(W24866), .A2(W14471), .ZN(W28783));
  NOR2X1 G2679 (.A1(I424), .A2(W19375), .ZN(O11242));
  NOR2X1 G2680 (.A1(W24066), .A2(W16610), .ZN(O11243));
  NOR2X1 G2681 (.A1(W1989), .A2(W2988), .ZN(O347));
  NOR2X1 G2682 (.A1(W31578), .A2(W33268), .ZN(W40923));
  NOR2X1 G2683 (.A1(W1934), .A2(W3634), .ZN(W9977));
  NOR2X1 G2684 (.A1(W4464), .A2(W5892), .ZN(W9946));
  NOR2X1 G2685 (.A1(I1647), .A2(W282), .ZN(W22005));
  NOR2X1 G2686 (.A1(W6165), .A2(W7650), .ZN(W9974));
  NOR2X1 G2687 (.A1(W8580), .A2(W1159), .ZN(W9972));
  NOR2X1 G2688 (.A1(W2592), .A2(W7850), .ZN(W9971));
  NOR2X1 G2689 (.A1(W2301), .A2(W5253), .ZN(W22007));
  NOR2X1 G2690 (.A1(W3591), .A2(W3169), .ZN(W9969));
  NOR2X1 G2691 (.A1(W7884), .A2(W2550), .ZN(W9967));
  NOR2X1 G2692 (.A1(W5015), .A2(W3524), .ZN(W22022));
  NOR2X1 G2693 (.A1(W6359), .A2(W6149), .ZN(W9923));
  NOR2X1 G2694 (.A1(W10568), .A2(W16715), .ZN(W40996));
  NOR2X1 G2695 (.A1(W6640), .A2(I271), .ZN(W9921));
  NOR2X1 G2696 (.A1(W3118), .A2(W4310), .ZN(W9920));
  NOR2X1 G2697 (.A1(W2193), .A2(W16053), .ZN(O2404));
  NOR2X1 G2698 (.A1(W38179), .A2(I1557), .ZN(W40999));
  NOR2X1 G2699 (.A1(W15039), .A2(W32306), .ZN(O11298));
  NOR2X1 G2700 (.A1(W6655), .A2(W6223), .ZN(O338));
  NOR2X1 G2701 (.A1(W30380), .A2(W32353), .ZN(W40990));
  NOR2X1 G2702 (.A1(W2763), .A2(I609), .ZN(W9913));
  NOR2X1 G2703 (.A1(W4873), .A2(I372), .ZN(W9912));
  NOR2X1 G2704 (.A1(W26444), .A2(W1717), .ZN(W41003));
  NOR2X1 G2705 (.A1(W985), .A2(W8089), .ZN(W28757));
  NOR2X1 G2706 (.A1(W12673), .A2(W127), .ZN(W41005));
  NOR2X1 G2707 (.A1(W29147), .A2(W39693), .ZN(W41006));
  NOR2X1 G2708 (.A1(W16290), .A2(W2022), .ZN(O4605));
  NOR2X1 G2709 (.A1(W1316), .A2(W4927), .ZN(W9906));
  NOR2X1 G2710 (.A1(W19424), .A2(W18397), .ZN(O11285));
  NOR2X1 G2711 (.A1(W20140), .A2(W35671), .ZN(O11274));
  NOR2X1 G2712 (.A1(W8143), .A2(W2043), .ZN(W9944));
  NOR2X1 G2713 (.A1(W3337), .A2(W19824), .ZN(O11275));
  NOR2X1 G2714 (.A1(W4681), .A2(W7917), .ZN(O11278));
  NOR2X1 G2715 (.A1(W635), .A2(W3453), .ZN(W9941));
  NOR2X1 G2716 (.A1(W15784), .A2(W16706), .ZN(W28765));
  NOR2X1 G2717 (.A1(I1065), .A2(W1904), .ZN(W9938));
  NOR2X1 G2718 (.A1(W14461), .A2(W11036), .ZN(O11283));
  NOR2X1 G2719 (.A1(W36188), .A2(W18888), .ZN(O11235));
  NOR2X1 G2720 (.A1(I456), .A2(W14307), .ZN(O11286));
  NOR2X1 G2721 (.A1(W7952), .A2(W27257), .ZN(O11287));
  NOR2X1 G2722 (.A1(W23361), .A2(W32371), .ZN(W40982));
  NOR2X1 G2723 (.A1(I635), .A2(W7124), .ZN(W9930));
  NOR2X1 G2724 (.A1(W26340), .A2(W39511), .ZN(O11292));
  NOR2X1 G2725 (.A1(W24431), .A2(W2913), .ZN(O11293));
  NOR2X1 G2726 (.A1(W6052), .A2(W5009), .ZN(O340));
  NOR2X1 G2727 (.A1(I52), .A2(W5026), .ZN(W10032));
  NOR2X1 G2728 (.A1(W4772), .A2(W7880), .ZN(W10040));
  NOR2X1 G2729 (.A1(W24008), .A2(W23157), .ZN(W28802));
  NOR2X1 G2730 (.A1(I658), .A2(W1228), .ZN(O11188));
  NOR2X1 G2731 (.A1(W4170), .A2(W16296), .ZN(O11189));
  NOR2X1 G2732 (.A1(W12166), .A2(W2574), .ZN(W40854));
  NOR2X1 G2733 (.A1(W11511), .A2(W879), .ZN(O11194));
  NOR2X1 G2734 (.A1(W26602), .A2(W35523), .ZN(O11195));
  NOR2X1 G2735 (.A1(W149), .A2(W17308), .ZN(O11196));
  NOR2X1 G2736 (.A1(W19517), .A2(W6018), .ZN(O2392));
  NOR2X1 G2737 (.A1(W7759), .A2(W3413), .ZN(O11197));
  NOR2X1 G2738 (.A1(W17817), .A2(W6966), .ZN(W21984));
  NOR2X1 G2739 (.A1(W4465), .A2(W28305), .ZN(O11200));
  NOR2X1 G2740 (.A1(W33139), .A2(W1956), .ZN(O11201));
  NOR2X1 G2741 (.A1(W7471), .A2(W18168), .ZN(W21986));
  NOR2X1 G2742 (.A1(W29541), .A2(W9249), .ZN(W40867));
  NOR2X1 G2743 (.A1(I1896), .A2(W6402), .ZN(W10024));
  NOR2X1 G2744 (.A1(W35741), .A2(W29424), .ZN(O11203));
  NOR2X1 G2745 (.A1(W37721), .A2(W40284), .ZN(W40833));
  NOR2X1 G2746 (.A1(W24546), .A2(W17230), .ZN(O4625));
  NOR2X1 G2747 (.A1(W10861), .A2(W26855), .ZN(W28808));
  NOR2X1 G2748 (.A1(W19742), .A2(W4018), .ZN(W21974));
  NOR2X1 G2749 (.A1(W15377), .A2(W8751), .ZN(W21975));
  NOR2X1 G2750 (.A1(W31792), .A2(W13290), .ZN(O11174));
  NOR2X1 G2751 (.A1(I1880), .A2(W5091), .ZN(W10052));
  NOR2X1 G2752 (.A1(W10434), .A2(W2424), .ZN(W21976));
  NOR2X1 G2753 (.A1(W17704), .A2(W28096), .ZN(O4624));
  NOR2X1 G2754 (.A1(W4454), .A2(W23756), .ZN(W28799));
  NOR2X1 G2755 (.A1(W16256), .A2(W6765), .ZN(W21978));
  NOR2X1 G2756 (.A1(W11042), .A2(W34435), .ZN(O11180));
  NOR2X1 G2757 (.A1(W15651), .A2(W6142), .ZN(W21979));
  NOR2X1 G2758 (.A1(W20007), .A2(W3049), .ZN(W28804));
  NOR2X1 G2759 (.A1(W1057), .A2(W2610), .ZN(W10044));
  NOR2X1 G2760 (.A1(W22573), .A2(W2928), .ZN(O11183));
  NOR2X1 G2761 (.A1(W10053), .A2(W14405), .ZN(W21981));
  NOR2X1 G2762 (.A1(W34768), .A2(W10712), .ZN(O11232));
  NOR2X1 G2763 (.A1(W5840), .A2(W1693), .ZN(W10003));
  NOR2X1 G2764 (.A1(W10177), .A2(W15610), .ZN(W21994));
  NOR2X1 G2765 (.A1(W23738), .A2(W24183), .ZN(W28793));
  NOR2X1 G2766 (.A1(W9143), .A2(I1098), .ZN(W9999));
  NOR2X1 G2767 (.A1(W1477), .A2(W26200), .ZN(W28791));
  NOR2X1 G2768 (.A1(W8229), .A2(W6880), .ZN(W9997));
  NOR2X1 G2769 (.A1(W8193), .A2(W17332), .ZN(W21997));
  NOR2X1 G2770 (.A1(W9094), .A2(W2696), .ZN(O4619));
  NOR2X1 G2771 (.A1(W14209), .A2(W12373), .ZN(O11221));
  NOR2X1 G2772 (.A1(W1579), .A2(I348), .ZN(W9993));
  NOR2X1 G2773 (.A1(W24802), .A2(W14649), .ZN(O4617));
  NOR2X1 G2774 (.A1(W1086), .A2(W24570), .ZN(W28786));
  NOR2X1 G2775 (.A1(W4435), .A2(W7628), .ZN(W9990));
  NOR2X1 G2776 (.A1(W32461), .A2(W37076), .ZN(O11234));
  NOR2X1 G2777 (.A1(W6887), .A2(W843), .ZN(W9988));
  NOR2X1 G2778 (.A1(W9042), .A2(W2874), .ZN(W9987));
  NOR2X1 G2779 (.A1(W23116), .A2(W459), .ZN(W40913));
  NOR2X1 G2780 (.A1(W32262), .A2(W17581), .ZN(W40886));
  NOR2X1 G2781 (.A1(W3824), .A2(W559), .ZN(W10021));
  NOR2X1 G2782 (.A1(W855), .A2(W21129), .ZN(W40876));
  NOR2X1 G2783 (.A1(W8079), .A2(W2687), .ZN(W10019));
  NOR2X1 G2784 (.A1(W3018), .A2(W3497), .ZN(W28798));
  NOR2X1 G2785 (.A1(W14735), .A2(W13790), .ZN(O11210));
  NOR2X1 G2786 (.A1(W25245), .A2(W40524), .ZN(O11212));
  NOR2X1 G2787 (.A1(W4337), .A2(W5616), .ZN(W10015));
  NOR2X1 G2788 (.A1(W17851), .A2(I1362), .ZN(O4621));
  NOR2X1 G2789 (.A1(W4258), .A2(W3645), .ZN(W9585));
  NOR2X1 G2790 (.A1(W38191), .A2(W40264), .ZN(W40888));
  NOR2X1 G2791 (.A1(W3545), .A2(W12084), .ZN(W21991));
  NOR2X1 G2792 (.A1(W3929), .A2(I1876), .ZN(O2393));
  NOR2X1 G2793 (.A1(W168), .A2(W3561), .ZN(W10008));
  NOR2X1 G2794 (.A1(W5247), .A2(W20855), .ZN(O11219));
  NOR2X1 G2795 (.A1(I1852), .A2(W4148), .ZN(W10006));
  NOR2X1 G2796 (.A1(W13454), .A2(W25185), .ZN(O11220));
  NOR2X1 G2797 (.A1(W22707), .A2(W747), .ZN(W41749));
  NOR2X1 G2798 (.A1(W8660), .A2(W6058), .ZN(W9167));
  NOR2X1 G2799 (.A1(W6344), .A2(W9846), .ZN(O11825));
  NOR2X1 G2800 (.A1(W7087), .A2(W8909), .ZN(W9164));
  NOR2X1 G2801 (.A1(W36103), .A2(W8893), .ZN(W41747));
  NOR2X1 G2802 (.A1(W6238), .A2(W1921), .ZN(W9162));
  NOR2X1 G2803 (.A1(W4202), .A2(I228), .ZN(W9161));
  NOR2X1 G2804 (.A1(I1698), .A2(W6473), .ZN(O271));
  NOR2X1 G2805 (.A1(W7782), .A2(W3354), .ZN(W9158));
  NOR2X1 G2806 (.A1(W5320), .A2(W15498), .ZN(W28499));
  NOR2X1 G2807 (.A1(W22), .A2(W5900), .ZN(W9156));
  NOR2X1 G2808 (.A1(W13455), .A2(W1243), .ZN(W22266));
  NOR2X1 G2809 (.A1(W6178), .A2(W2047), .ZN(W9154));
  NOR2X1 G2810 (.A1(W40952), .A2(W21364), .ZN(W41751));
  NOR2X1 G2811 (.A1(W9508), .A2(W20963), .ZN(O11829));
  NOR2X1 G2812 (.A1(W1327), .A2(W7149), .ZN(W9151));
  NOR2X1 G2813 (.A1(W693), .A2(W8545), .ZN(W9150));
  NOR2X1 G2814 (.A1(W3933), .A2(W21310), .ZN(W22267));
  NOR2X1 G2815 (.A1(W16514), .A2(W27527), .ZN(W28500));
  NOR2X1 G2816 (.A1(W20194), .A2(W11382), .ZN(W41735));
  NOR2X1 G2817 (.A1(I636), .A2(W774), .ZN(O11819));
  NOR2X1 G2818 (.A1(I1611), .A2(W1472), .ZN(O11820));
  NOR2X1 G2819 (.A1(W224), .A2(W1839), .ZN(W9181));
  NOR2X1 G2820 (.A1(W9608), .A2(W24663), .ZN(W28503));
  NOR2X1 G2821 (.A1(W2743), .A2(I1571), .ZN(O4522));
  NOR2X1 G2822 (.A1(I1247), .A2(W2045), .ZN(W9178));
  NOR2X1 G2823 (.A1(W8412), .A2(W6823), .ZN(W9177));
  NOR2X1 G2824 (.A1(W8582), .A2(W5754), .ZN(O2461));
  NOR2X1 G2825 (.A1(W4801), .A2(W8082), .ZN(W9175));
  NOR2X1 G2826 (.A1(W6349), .A2(I276), .ZN(W9174));
  NOR2X1 G2827 (.A1(W5432), .A2(W4249), .ZN(W9173));
  NOR2X1 G2828 (.A1(W2712), .A2(W6444), .ZN(W9172));
  NOR2X1 G2829 (.A1(W6844), .A2(W22151), .ZN(W22262));
  NOR2X1 G2830 (.A1(W3421), .A2(W1452), .ZN(W9170));
  NOR2X1 G2831 (.A1(I389), .A2(I1386), .ZN(W9169));
  NOR2X1 G2832 (.A1(W31923), .A2(W2428), .ZN(O11862));
  NOR2X1 G2833 (.A1(I1299), .A2(W5043), .ZN(W9126));
  NOR2X1 G2834 (.A1(W26757), .A2(W25093), .ZN(O11848));
  NOR2X1 G2835 (.A1(W5990), .A2(W7), .ZN(W9124));
  NOR2X1 G2836 (.A1(W17906), .A2(W1535), .ZN(O11849));
  NOR2X1 G2837 (.A1(W6032), .A2(W9089), .ZN(W9121));
  NOR2X1 G2838 (.A1(W39439), .A2(W29027), .ZN(W41791));
  NOR2X1 G2839 (.A1(W4322), .A2(W4873), .ZN(W9118));
  NOR2X1 G2840 (.A1(I708), .A2(W28886), .ZN(O11861));
  NOR2X1 G2841 (.A1(W322), .A2(W5848), .ZN(W9128));
  NOR2X1 G2842 (.A1(W24533), .A2(W36093), .ZN(W41800));
  NOR2X1 G2843 (.A1(W23343), .A2(W9132), .ZN(W28483));
  NOR2X1 G2844 (.A1(W18729), .A2(W33764), .ZN(W41804));
  NOR2X1 G2845 (.A1(W929), .A2(W4646), .ZN(W9112));
  NOR2X1 G2846 (.A1(W4427), .A2(W7677), .ZN(W22280));
  NOR2X1 G2847 (.A1(W8619), .A2(W2575), .ZN(O264));
  NOR2X1 G2848 (.A1(I486), .A2(W4298), .ZN(O2465));
  NOR2X1 G2849 (.A1(W8702), .A2(W3108), .ZN(W9108));
  NOR2X1 G2850 (.A1(W3907), .A2(W5486), .ZN(W9138));
  NOR2X1 G2851 (.A1(W1177), .A2(I390), .ZN(W9147));
  NOR2X1 G2852 (.A1(W19032), .A2(W13614), .ZN(O11833));
  NOR2X1 G2853 (.A1(W17297), .A2(W33853), .ZN(O11834));
  NOR2X1 G2854 (.A1(W6731), .A2(W19476), .ZN(O11836));
  NOR2X1 G2855 (.A1(W27541), .A2(W26032), .ZN(O4520));
  NOR2X1 G2856 (.A1(W15091), .A2(I1580), .ZN(W28492));
  NOR2X1 G2857 (.A1(I994), .A2(W39545), .ZN(O11838));
  NOR2X1 G2858 (.A1(W17577), .A2(W21275), .ZN(W22272));
  NOR2X1 G2859 (.A1(W4737), .A2(W5966), .ZN(W9186));
  NOR2X1 G2860 (.A1(W2407), .A2(W3481), .ZN(W9137));
  NOR2X1 G2861 (.A1(W10844), .A2(W28147), .ZN(O11843));
  NOR2X1 G2862 (.A1(W25811), .A2(W6420), .ZN(W41772));
  NOR2X1 G2863 (.A1(W4876), .A2(I489), .ZN(O267));
  NOR2X1 G2864 (.A1(W9144), .A2(W34572), .ZN(O11845));
  NOR2X1 G2865 (.A1(W11432), .A2(W927), .ZN(W28490));
  NOR2X1 G2866 (.A1(W41038), .A2(W8867), .ZN(O11846));
  NOR2X1 G2867 (.A1(W8526), .A2(W8901), .ZN(W9237));
  NOR2X1 G2868 (.A1(W20616), .A2(W12753), .ZN(O2458));
  NOR2X1 G2869 (.A1(W34867), .A2(W35160), .ZN(O11777));
  NOR2X1 G2870 (.A1(W21378), .A2(W8503), .ZN(W28520));
  NOR2X1 G2871 (.A1(W8349), .A2(W7264), .ZN(W22240));
  NOR2X1 G2872 (.A1(W5997), .A2(W5825), .ZN(W41681));
  NOR2X1 G2873 (.A1(W8445), .A2(W1448), .ZN(W9240));
  NOR2X1 G2874 (.A1(I52), .A2(W28613), .ZN(O11779));
  NOR2X1 G2875 (.A1(W14584), .A2(W6460), .ZN(W41683));
  NOR2X1 G2876 (.A1(W3906), .A2(W3354), .ZN(W9247));
  NOR2X1 G2877 (.A1(W8322), .A2(W321), .ZN(W9236));
  NOR2X1 G2878 (.A1(W40845), .A2(W36215), .ZN(O11780));
  NOR2X1 G2879 (.A1(W23528), .A2(W33669), .ZN(W41686));
  NOR2X1 G2880 (.A1(W2944), .A2(W7610), .ZN(W22241));
  NOR2X1 G2881 (.A1(W1171), .A2(W6515), .ZN(W9232));
  NOR2X1 G2882 (.A1(W5480), .A2(W6416), .ZN(O4527));
  NOR2X1 G2883 (.A1(W4010), .A2(W6901), .ZN(W9230));
  NOR2X1 G2884 (.A1(W38350), .A2(W10694), .ZN(O11785));
  NOR2X1 G2885 (.A1(W4798), .A2(W7375), .ZN(W9255));
  NOR2X1 G2886 (.A1(W14685), .A2(W1978), .ZN(O4529));
  NOR2X1 G2887 (.A1(W10722), .A2(W38781), .ZN(W41665));
  NOR2X1 G2888 (.A1(W148), .A2(W6188), .ZN(O277));
  NOR2X1 G2889 (.A1(I829), .A2(W8356), .ZN(W28527));
  NOR2X1 G2890 (.A1(W3217), .A2(W29762), .ZN(O11773));
  NOR2X1 G2891 (.A1(W27462), .A2(W650), .ZN(O4528));
  NOR2X1 G2892 (.A1(W1403), .A2(W651), .ZN(W9257));
  NOR2X1 G2893 (.A1(W15914), .A2(W18772), .ZN(W22234));
  NOR2X1 G2894 (.A1(W2891), .A2(W2799), .ZN(W9228));
  NOR2X1 G2895 (.A1(W1916), .A2(I943), .ZN(W9254));
  NOR2X1 G2896 (.A1(W7919), .A2(W2591), .ZN(W28523));
  NOR2X1 G2897 (.A1(W35950), .A2(W30611), .ZN(W41673));
  NOR2X1 G2898 (.A1(W5814), .A2(W31059), .ZN(O11775));
  NOR2X1 G2899 (.A1(I965), .A2(W2698), .ZN(W9250));
  NOR2X1 G2900 (.A1(W10764), .A2(W13830), .ZN(O2457));
  NOR2X1 G2901 (.A1(W5790), .A2(W8950), .ZN(W9248));
  NOR2X1 G2902 (.A1(W24636), .A2(W16066), .ZN(O11804));
  NOR2X1 G2903 (.A1(W12215), .A2(W12229), .ZN(O11798));
  NOR2X1 G2904 (.A1(W2354), .A2(I472), .ZN(W9208));
  NOR2X1 G2905 (.A1(W12401), .A2(W22883), .ZN(W28515));
  NOR2X1 G2906 (.A1(W7473), .A2(W6284), .ZN(O4525));
  NOR2X1 G2907 (.A1(W3130), .A2(W8056), .ZN(W9205));
  NOR2X1 G2908 (.A1(W29294), .A2(W3483), .ZN(W41714));
  NOR2X1 G2909 (.A1(W12540), .A2(W32280), .ZN(O11802));
  NOR2X1 G2910 (.A1(W23631), .A2(W8705), .ZN(O11803));
  NOR2X1 G2911 (.A1(W3276), .A2(W8574), .ZN(W9210));
  NOR2X1 G2912 (.A1(W1628), .A2(I1540), .ZN(W9198));
  NOR2X1 G2913 (.A1(W1286), .A2(W3283), .ZN(O274));
  NOR2X1 G2914 (.A1(W13197), .A2(W32751), .ZN(W41722));
  NOR2X1 G2915 (.A1(W16522), .A2(W4249), .ZN(O11811));
  NOR2X1 G2916 (.A1(W4992), .A2(W6252), .ZN(O273));
  NOR2X1 G2917 (.A1(W20920), .A2(W12747), .ZN(W22254));
  NOR2X1 G2918 (.A1(I714), .A2(W20674), .ZN(W22255));
  NOR2X1 G2919 (.A1(W5424), .A2(W9742), .ZN(W22257));
  NOR2X1 G2920 (.A1(W14106), .A2(W1829), .ZN(W28517));
  NOR2X1 G2921 (.A1(W16926), .A2(W4418), .ZN(W41694));
  NOR2X1 G2922 (.A1(W3629), .A2(W1200), .ZN(W9226));
  NOR2X1 G2923 (.A1(W26954), .A2(W4625), .ZN(O11788));
  NOR2X1 G2924 (.A1(W55), .A2(W7779), .ZN(W9224));
  NOR2X1 G2925 (.A1(W909), .A2(W1011), .ZN(W9223));
  NOR2X1 G2926 (.A1(W28952), .A2(W7501), .ZN(O11789));
  NOR2X1 G2927 (.A1(W15013), .A2(W33557), .ZN(W41700));
  NOR2X1 G2928 (.A1(W29255), .A2(W28896), .ZN(O11791));
  NOR2X1 G2929 (.A1(W36599), .A2(W8881), .ZN(W41807));
  NOR2X1 G2930 (.A1(W21996), .A2(W6729), .ZN(W22245));
  NOR2X1 G2931 (.A1(W5179), .A2(W6359), .ZN(W22246));
  NOR2X1 G2932 (.A1(W516), .A2(W5006), .ZN(W9215));
  NOR2X1 G2933 (.A1(W3738), .A2(W5267), .ZN(W9214));
  NOR2X1 G2934 (.A1(W26891), .A2(I820), .ZN(O11795));
  NOR2X1 G2935 (.A1(W29611), .A2(W32669), .ZN(O11796));
  NOR2X1 G2936 (.A1(W25464), .A2(W21006), .ZN(O11797));
  NOR2X1 G2937 (.A1(W18639), .A2(I1428), .ZN(W22312));
  NOR2X1 G2938 (.A1(W24285), .A2(W21666), .ZN(O11934));
  NOR2X1 G2939 (.A1(I1935), .A2(W816), .ZN(O4505));
  NOR2X1 G2940 (.A1(W24982), .A2(W6224), .ZN(O11935));
  NOR2X1 G2941 (.A1(W29258), .A2(W14598), .ZN(O11937));
  NOR2X1 G2942 (.A1(W41543), .A2(W25272), .ZN(O11938));
  NOR2X1 G2943 (.A1(W74), .A2(W14508), .ZN(O2477));
  NOR2X1 G2944 (.A1(W32426), .A2(W41350), .ZN(W41906));
  NOR2X1 G2945 (.A1(W115), .A2(W5048), .ZN(O4504));
  NOR2X1 G2946 (.A1(W7922), .A2(W1006), .ZN(W9012));
  NOR2X1 G2947 (.A1(W39726), .A2(W3595), .ZN(W41911));
  NOR2X1 G2948 (.A1(W2574), .A2(W8029), .ZN(W9001));
  NOR2X1 G2949 (.A1(W8276), .A2(W2850), .ZN(W9000));
  NOR2X1 G2950 (.A1(W35697), .A2(W7416), .ZN(O11943));
  NOR2X1 G2951 (.A1(W14356), .A2(I1528), .ZN(W28444));
  NOR2X1 G2952 (.A1(W33517), .A2(W34678), .ZN(O11947));
  NOR2X1 G2953 (.A1(W25349), .A2(W4724), .ZN(W28442));
  NOR2X1 G2954 (.A1(W29902), .A2(W22124), .ZN(O11950));
  NOR2X1 G2955 (.A1(W356), .A2(I640), .ZN(W9021));
  NOR2X1 G2956 (.A1(W37650), .A2(W33521), .ZN(O11919));
  NOR2X1 G2957 (.A1(W31237), .A2(W21428), .ZN(W41883));
  NOR2X1 G2958 (.A1(W6840), .A2(W2121), .ZN(O2474));
  NOR2X1 G2959 (.A1(W15974), .A2(W2304), .ZN(O11922));
  NOR2X1 G2960 (.A1(W27303), .A2(W22098), .ZN(O11924));
  NOR2X1 G2961 (.A1(W24080), .A2(W14242), .ZN(O11925));
  NOR2X1 G2962 (.A1(W5937), .A2(W773), .ZN(W9023));
  NOR2X1 G2963 (.A1(W1711), .A2(W3702), .ZN(W9022));
  NOR2X1 G2964 (.A1(W2127), .A2(I1217), .ZN(W41920));
  NOR2X1 G2965 (.A1(I324), .A2(W4828), .ZN(W9020));
  NOR2X1 G2966 (.A1(W8498), .A2(W4571), .ZN(W9019));
  NOR2X1 G2967 (.A1(W28063), .A2(W10497), .ZN(O4506));
  NOR2X1 G2968 (.A1(W19764), .A2(W9280), .ZN(O11930));
  NOR2X1 G2969 (.A1(W748), .A2(W1770), .ZN(W9015));
  NOR2X1 G2970 (.A1(W17325), .A2(W31243), .ZN(O11932));
  NOR2X1 G2971 (.A1(W4578), .A2(W1477), .ZN(W9013));
  NOR2X1 G2972 (.A1(W30538), .A2(W13122), .ZN(O11976));
  NOR2X1 G2973 (.A1(W18061), .A2(W3492), .ZN(W22325));
  NOR2X1 G2974 (.A1(W7193), .A2(W22472), .ZN(O4496));
  NOR2X1 G2975 (.A1(W38258), .A2(W30091), .ZN(O11971));
  NOR2X1 G2976 (.A1(W1440), .A2(W1903), .ZN(W8966));
  NOR2X1 G2977 (.A1(W5875), .A2(W18402), .ZN(O4495));
  NOR2X1 G2978 (.A1(W41656), .A2(W2733), .ZN(O11975));
  NOR2X1 G2979 (.A1(W3222), .A2(W2647), .ZN(W8962));
  NOR2X1 G2980 (.A1(W171), .A2(W8559), .ZN(W8961));
  NOR2X1 G2981 (.A1(W23568), .A2(W25621), .ZN(O11968));
  NOR2X1 G2982 (.A1(W6997), .A2(W3716), .ZN(W28425));
  NOR2X1 G2983 (.A1(W1681), .A2(I1954), .ZN(W8957));
  NOR2X1 G2984 (.A1(W4261), .A2(W4489), .ZN(W8956));
  NOR2X1 G2985 (.A1(W6223), .A2(W2943), .ZN(W8955));
  NOR2X1 G2986 (.A1(W957), .A2(W8064), .ZN(W22331));
  NOR2X1 G2987 (.A1(W6114), .A2(W8123), .ZN(O259));
  NOR2X1 G2988 (.A1(W4185), .A2(W7473), .ZN(W8950));
  NOR2X1 G2989 (.A1(I1865), .A2(W3495), .ZN(W8949));
  NOR2X1 G2990 (.A1(W21983), .A2(W1286), .ZN(O11962));
  NOR2X1 G2991 (.A1(W21753), .A2(W36755), .ZN(O11952));
  NOR2X1 G2992 (.A1(W19535), .A2(W3723), .ZN(O11954));
  NOR2X1 G2993 (.A1(W34770), .A2(W40640), .ZN(O11955));
  NOR2X1 G2994 (.A1(W3597), .A2(W38876), .ZN(W41926));
  NOR2X1 G2995 (.A1(W12223), .A2(W15117), .ZN(O2479));
  NOR2X1 G2996 (.A1(W10020), .A2(W24828), .ZN(O11958));
  NOR2X1 G2997 (.A1(W2980), .A2(I1110), .ZN(O4501));
  NOR2X1 G2998 (.A1(W9249), .A2(W29729), .ZN(O11959));
  NOR2X1 G2999 (.A1(W6666), .A2(W1442), .ZN(W9032));
  NOR2X1 G3000 (.A1(W8546), .A2(I372), .ZN(O11964));
  NOR2X1 G3001 (.A1(W6874), .A2(I753), .ZN(W8978));
  NOR2X1 G3002 (.A1(W4505), .A2(I4), .ZN(W8977));
  NOR2X1 G3003 (.A1(W40304), .A2(W28441), .ZN(W41938));
  NOR2X1 G3004 (.A1(W16587), .A2(W10399), .ZN(O2481));
  NOR2X1 G3005 (.A1(W26152), .A2(W37140), .ZN(O11966));
  NOR2X1 G3006 (.A1(W18121), .A2(W20515), .ZN(W41942));
  NOR2X1 G3007 (.A1(W19977), .A2(W23270), .ZN(W41835));
  NOR2X1 G3008 (.A1(W4727), .A2(I256), .ZN(W9087));
  NOR2X1 G3009 (.A1(W21211), .A2(W4876), .ZN(W28477));
  NOR2X1 G3010 (.A1(W15485), .A2(W1779), .ZN(W28476));
  NOR2X1 G3011 (.A1(W6758), .A2(W21978), .ZN(W28474));
  NOR2X1 G3012 (.A1(W6912), .A2(I460), .ZN(W9083));
  NOR2X1 G3013 (.A1(W7874), .A2(W5643), .ZN(W9082));
  NOR2X1 G3014 (.A1(W486), .A2(I502), .ZN(W28473));
  NOR2X1 G3015 (.A1(W8992), .A2(W23051), .ZN(O11884));
  NOR2X1 G3016 (.A1(W6923), .A2(W725), .ZN(W9088));
  NOR2X1 G3017 (.A1(W23911), .A2(W14872), .ZN(W28471));
  NOR2X1 G3018 (.A1(W15311), .A2(W19106), .ZN(O11891));
  NOR2X1 G3019 (.A1(W41573), .A2(W23334), .ZN(O11892));
  NOR2X1 G3020 (.A1(W5801), .A2(I1078), .ZN(W9074));
  NOR2X1 G3021 (.A1(W2601), .A2(W22880), .ZN(O11893));
  NOR2X1 G3022 (.A1(W2624), .A2(W2142), .ZN(W9072));
  NOR2X1 G3023 (.A1(I1100), .A2(W16686), .ZN(W28470));
  NOR2X1 G3024 (.A1(W38821), .A2(W12582), .ZN(O11895));
  NOR2X1 G3025 (.A1(W30501), .A2(W38774), .ZN(O11875));
  NOR2X1 G3026 (.A1(I1599), .A2(W5898), .ZN(W9106));
  NOR2X1 G3027 (.A1(W2645), .A2(W14345), .ZN(O11868));
  NOR2X1 G3028 (.A1(W3079), .A2(W1764), .ZN(O11870));
  NOR2X1 G3029 (.A1(W1863), .A2(W9091), .ZN(W9103));
  NOR2X1 G3030 (.A1(W20905), .A2(W2017), .ZN(W22283));
  NOR2X1 G3031 (.A1(W7579), .A2(W41171), .ZN(O11874));
  NOR2X1 G3032 (.A1(I1339), .A2(W5876), .ZN(W9099));
  NOR2X1 G3033 (.A1(W3809), .A2(I597), .ZN(O263));
  NOR2X1 G3034 (.A1(W40320), .A2(W38346), .ZN(O11897));
  NOR2X1 G3035 (.A1(W6222), .A2(W7407), .ZN(W9096));
  NOR2X1 G3036 (.A1(W43), .A2(W7077), .ZN(W9095));
  NOR2X1 G3037 (.A1(W27374), .A2(W24028), .ZN(O4516));
  NOR2X1 G3038 (.A1(W33590), .A2(W37585), .ZN(W41820));
  NOR2X1 G3039 (.A1(W8792), .A2(W2525), .ZN(W9091));
  NOR2X1 G3040 (.A1(W26726), .A2(W11609), .ZN(O4515));
  NOR2X1 G3041 (.A1(W37626), .A2(W30252), .ZN(W41823));
  NOR2X1 G3042 (.A1(W16938), .A2(I1977), .ZN(W28457));
  NOR2X1 G3043 (.A1(I1031), .A2(I574), .ZN(W9050));
  NOR2X1 G3044 (.A1(W27314), .A2(W31851), .ZN(W41864));
  NOR2X1 G3045 (.A1(W18247), .A2(I1247), .ZN(O4513));
  NOR2X1 G3046 (.A1(W23062), .A2(W13550), .ZN(O4512));
  NOR2X1 G3047 (.A1(W23420), .A2(W32179), .ZN(O11910));
  NOR2X1 G3048 (.A1(W6632), .A2(W32402), .ZN(W41869));
  NOR2X1 G3049 (.A1(W20531), .A2(W21367), .ZN(O11912));
  NOR2X1 G3050 (.A1(W2442), .A2(W25126), .ZN(O4511));
  NOR2X1 G3051 (.A1(I1928), .A2(W718), .ZN(W9051));
  NOR2X1 G3052 (.A1(W6046), .A2(W31353), .ZN(O11916));
  NOR2X1 G3053 (.A1(W8087), .A2(W3610), .ZN(W9039));
  NOR2X1 G3054 (.A1(W2152), .A2(W543), .ZN(W9038));
  NOR2X1 G3055 (.A1(W3538), .A2(W1493), .ZN(W9037));
  NOR2X1 G3056 (.A1(W20624), .A2(W814), .ZN(O4509));
  NOR2X1 G3057 (.A1(W41827), .A2(W6811), .ZN(O11917));
  NOR2X1 G3058 (.A1(W158), .A2(W4435), .ZN(W9034));
  NOR2X1 G3059 (.A1(W5836), .A2(W13792), .ZN(O4508));
  NOR2X1 G3060 (.A1(W8460), .A2(W7584), .ZN(W9059));
  NOR2X1 G3061 (.A1(W40056), .A2(W23796), .ZN(O11898));
  NOR2X1 G3062 (.A1(W10768), .A2(W2644), .ZN(O11899));
  NOR2X1 G3063 (.A1(W8658), .A2(W1879), .ZN(W9065));
  NOR2X1 G3064 (.A1(W34412), .A2(W6670), .ZN(O11900));
  NOR2X1 G3065 (.A1(W16818), .A2(W8062), .ZN(O11901));
  NOR2X1 G3066 (.A1(I76), .A2(W4366), .ZN(W9062));
  NOR2X1 G3067 (.A1(W2953), .A2(W4777), .ZN(W9061));
  NOR2X1 G3068 (.A1(W3709), .A2(W34049), .ZN(O11902));
  NOR2X1 G3069 (.A1(W985), .A2(W5173), .ZN(W22230));
  NOR2X1 G3070 (.A1(W2225), .A2(I1188), .ZN(W28468));
  NOR2X1 G3071 (.A1(W953), .A2(W5354), .ZN(W9057));
  NOR2X1 G3072 (.A1(W39666), .A2(W37430), .ZN(O11905));
  NOR2X1 G3073 (.A1(W23648), .A2(W1359), .ZN(W28467));
  NOR2X1 G3074 (.A1(W14302), .A2(W21635), .ZN(O11907));
  NOR2X1 G3075 (.A1(W317), .A2(W5643), .ZN(W9053));
  NOR2X1 G3076 (.A1(W2532), .A2(W3862), .ZN(W9052));
  NOR2X1 G3077 (.A1(W913), .A2(W2517), .ZN(O11615));
  NOR2X1 G3078 (.A1(W1411), .A2(W5843), .ZN(W9486));
  NOR2X1 G3079 (.A1(W2039), .A2(W1653), .ZN(W9485));
  NOR2X1 G3080 (.A1(W23990), .A2(W2418), .ZN(O11605));
  NOR2X1 G3081 (.A1(W8277), .A2(W9023), .ZN(W28619));
  NOR2X1 G3082 (.A1(W18828), .A2(W7746), .ZN(W28618));
  NOR2X1 G3083 (.A1(W38340), .A2(W4097), .ZN(O11613));
  NOR2X1 G3084 (.A1(W3333), .A2(W7215), .ZN(W9477));
  NOR2X1 G3085 (.A1(W6645), .A2(W879), .ZN(W9476));
  NOR2X1 G3086 (.A1(W30135), .A2(W4937), .ZN(O11604));
  NOR2X1 G3087 (.A1(W9367), .A2(W614), .ZN(W22161));
  NOR2X1 G3088 (.A1(W28733), .A2(W21737), .ZN(O11620));
  NOR2X1 G3089 (.A1(W9785), .A2(W37376), .ZN(W41462));
  NOR2X1 G3090 (.A1(I0), .A2(W16329), .ZN(O4557));
  NOR2X1 G3091 (.A1(W4383), .A2(W7740), .ZN(W9469));
  NOR2X1 G3092 (.A1(W8902), .A2(W8762), .ZN(W9468));
  NOR2X1 G3093 (.A1(W4367), .A2(W3175), .ZN(O293));
  NOR2X1 G3094 (.A1(W25827), .A2(W22966), .ZN(O11623));
  NOR2X1 G3095 (.A1(W7194), .A2(W7930), .ZN(W9499));
  NOR2X1 G3096 (.A1(I1810), .A2(W5525), .ZN(W22141));
  NOR2X1 G3097 (.A1(W23382), .A2(W7604), .ZN(W28631));
  NOR2X1 G3098 (.A1(W26004), .A2(W20281), .ZN(W28630));
  NOR2X1 G3099 (.A1(W2031), .A2(W5438), .ZN(W9506));
  NOR2X1 G3100 (.A1(W15282), .A2(W7335), .ZN(W22145));
  NOR2X1 G3101 (.A1(W29396), .A2(W17493), .ZN(O11589));
  NOR2X1 G3102 (.A1(W6489), .A2(W3412), .ZN(W9502));
  NOR2X1 G3103 (.A1(W14537), .A2(W14272), .ZN(W22148));
  NOR2X1 G3104 (.A1(W21429), .A2(W15276), .ZN(W22164));
  NOR2X1 G3105 (.A1(W18980), .A2(W13605), .ZN(W22149));
  NOR2X1 G3106 (.A1(W5806), .A2(W3390), .ZN(O295));
  NOR2X1 G3107 (.A1(W24315), .A2(W27896), .ZN(W28627));
  NOR2X1 G3108 (.A1(W40990), .A2(I1364), .ZN(W41432));
  NOR2X1 G3109 (.A1(W121), .A2(I1190), .ZN(W28623));
  NOR2X1 G3110 (.A1(W37607), .A2(W30476), .ZN(W41434));
  NOR2X1 G3111 (.A1(W22703), .A2(W38060), .ZN(O11601));
  NOR2X1 G3112 (.A1(W6519), .A2(W1922), .ZN(O290));
  NOR2X1 G3113 (.A1(W32794), .A2(W34632), .ZN(O11636));
  NOR2X1 G3114 (.A1(W12933), .A2(W22018), .ZN(W41488));
  NOR2X1 G3115 (.A1(W9012), .A2(W3631), .ZN(O291));
  NOR2X1 G3116 (.A1(W7424), .A2(W2467), .ZN(W9443));
  NOR2X1 G3117 (.A1(W1960), .A2(W5652), .ZN(W9442));
  NOR2X1 G3118 (.A1(W22331), .A2(W18517), .ZN(O11637));
  NOR2X1 G3119 (.A1(W9364), .A2(W24172), .ZN(O11638));
  NOR2X1 G3120 (.A1(W34835), .A2(W5502), .ZN(O11641));
  NOR2X1 G3121 (.A1(W37162), .A2(W20524), .ZN(W41486));
  NOR2X1 G3122 (.A1(W14073), .A2(W24980), .ZN(W28599));
  NOR2X1 G3123 (.A1(W20614), .A2(I1110), .ZN(O2438));
  NOR2X1 G3124 (.A1(W8213), .A2(I1146), .ZN(O11644));
  NOR2X1 G3125 (.A1(W789), .A2(W996), .ZN(W9433));
  NOR2X1 G3126 (.A1(I1998), .A2(W8697), .ZN(W9432));
  NOR2X1 G3127 (.A1(W4809), .A2(W3851), .ZN(W9431));
  NOR2X1 G3128 (.A1(W38241), .A2(W30985), .ZN(O11646));
  NOR2X1 G3129 (.A1(W3058), .A2(W41134), .ZN(O11649));
  NOR2X1 G3130 (.A1(W3907), .A2(W16807), .ZN(W28601));
  NOR2X1 G3131 (.A1(W6087), .A2(W9040), .ZN(W9464));
  NOR2X1 G3132 (.A1(W8925), .A2(W25667), .ZN(O11626));
  NOR2X1 G3133 (.A1(W3941), .A2(W32566), .ZN(O11627));
  NOR2X1 G3134 (.A1(W9511), .A2(W11903), .ZN(O11628));
  NOR2X1 G3135 (.A1(W3397), .A2(W6775), .ZN(W22166));
  NOR2X1 G3136 (.A1(W17174), .A2(W39812), .ZN(O11629));
  NOR2X1 G3137 (.A1(W13390), .A2(W7111), .ZN(O2435));
  NOR2X1 G3138 (.A1(W13082), .A2(W19790), .ZN(W28602));
  NOR2X1 G3139 (.A1(W8988), .A2(W4724), .ZN(W9511));
  NOR2X1 G3140 (.A1(W6432), .A2(W5648), .ZN(O11633));
  NOR2X1 G3141 (.A1(W1082), .A2(W8827), .ZN(W9453));
  NOR2X1 G3142 (.A1(W3114), .A2(W7637), .ZN(W9452));
  NOR2X1 G3143 (.A1(W9510), .A2(W6646), .ZN(W22170));
  NOR2X1 G3144 (.A1(W1097), .A2(W6595), .ZN(W9450));
  NOR2X1 G3145 (.A1(W16110), .A2(W21491), .ZN(W41483));
  NOR2X1 G3146 (.A1(W415), .A2(W3699), .ZN(W9448));
  NOR2X1 G3147 (.A1(W5303), .A2(W9799), .ZN(O11552));
  NOR2X1 G3148 (.A1(W10548), .A2(W4773), .ZN(W22121));
  NOR2X1 G3149 (.A1(W24421), .A2(W25657), .ZN(O11545));
  NOR2X1 G3150 (.A1(W54), .A2(W3143), .ZN(W9565));
  NOR2X1 G3151 (.A1(W13690), .A2(W21587), .ZN(O11547));
  NOR2X1 G3152 (.A1(W20214), .A2(W1199), .ZN(O4569));
  NOR2X1 G3153 (.A1(W19780), .A2(W71), .ZN(W28651));
  NOR2X1 G3154 (.A1(W37546), .A2(W10327), .ZN(O11551));
  NOR2X1 G3155 (.A1(W6700), .A2(W5398), .ZN(W9560));
  NOR2X1 G3156 (.A1(W186), .A2(W3040), .ZN(W9568));
  NOR2X1 G3157 (.A1(W28608), .A2(W35726), .ZN(W41371));
  NOR2X1 G3158 (.A1(W26420), .A2(W20396), .ZN(W28649));
  NOR2X1 G3159 (.A1(W17023), .A2(W9292), .ZN(W22125));
  NOR2X1 G3160 (.A1(W35704), .A2(W16549), .ZN(W41375));
  NOR2X1 G3161 (.A1(W3119), .A2(I1629), .ZN(W9554));
  NOR2X1 G3162 (.A1(W30613), .A2(W20676), .ZN(O11556));
  NOR2X1 G3163 (.A1(W18257), .A2(W3030), .ZN(W28648));
  NOR2X1 G3164 (.A1(W8214), .A2(I1740), .ZN(W9551));
  NOR2X1 G3165 (.A1(W20073), .A2(W16333), .ZN(O2429));
  NOR2X1 G3166 (.A1(W7298), .A2(W386), .ZN(O302));
  NOR2X1 G3167 (.A1(W14726), .A2(W2481), .ZN(W22117));
  NOR2X1 G3168 (.A1(W38581), .A2(W39439), .ZN(O11531));
  NOR2X1 G3169 (.A1(W6448), .A2(I1141), .ZN(W9581));
  NOR2X1 G3170 (.A1(W20841), .A2(W30832), .ZN(O11533));
  NOR2X1 G3171 (.A1(W19591), .A2(W21725), .ZN(W22118));
  NOR2X1 G3172 (.A1(W38468), .A2(W25473), .ZN(O11534));
  NOR2X1 G3173 (.A1(W24000), .A2(W37035), .ZN(O11535));
  NOR2X1 G3174 (.A1(W4500), .A2(W16455), .ZN(W22128));
  NOR2X1 G3175 (.A1(W19475), .A2(W11695), .ZN(O2430));
  NOR2X1 G3176 (.A1(W17763), .A2(W35838), .ZN(O11538));
  NOR2X1 G3177 (.A1(W2980), .A2(W3547), .ZN(W9573));
  NOR2X1 G3178 (.A1(W3007), .A2(W35584), .ZN(O11540));
  NOR2X1 G3179 (.A1(W3560), .A2(W5725), .ZN(O300));
  NOR2X1 G3180 (.A1(W16306), .A2(I846), .ZN(O11541));
  NOR2X1 G3181 (.A1(W19496), .A2(W25040), .ZN(O11542));
  NOR2X1 G3182 (.A1(W3359), .A2(I1712), .ZN(W9521));
  NOR2X1 G3183 (.A1(I424), .A2(W4474), .ZN(W9530));
  NOR2X1 G3184 (.A1(W26649), .A2(W16677), .ZN(O11567));
  NOR2X1 G3185 (.A1(W9264), .A2(W5721), .ZN(W9528));
  NOR2X1 G3186 (.A1(I1749), .A2(W16812), .ZN(O11568));
  NOR2X1 G3187 (.A1(W14133), .A2(W11111), .ZN(W28638));
  NOR2X1 G3188 (.A1(W8623), .A2(W16977), .ZN(O4563));
  NOR2X1 G3189 (.A1(W20518), .A2(W1105), .ZN(O11570));
  NOR2X1 G3190 (.A1(W7775), .A2(W762), .ZN(W9523));
  NOR2X1 G3191 (.A1(I1328), .A2(I34), .ZN(W9531));
  NOR2X1 G3192 (.A1(W36518), .A2(W26964), .ZN(O11572));
  NOR2X1 G3193 (.A1(W37214), .A2(W17876), .ZN(O11573));
  NOR2X1 G3194 (.A1(W3202), .A2(W18034), .ZN(W22138));
  NOR2X1 G3195 (.A1(W13214), .A2(W18030), .ZN(W22139));
  NOR2X1 G3196 (.A1(W21986), .A2(W13372), .ZN(W22140));
  NOR2X1 G3197 (.A1(W23534), .A2(W15259), .ZN(O11579));
  NOR2X1 G3198 (.A1(W34615), .A2(W38824), .ZN(O11581));
  NOR2X1 G3199 (.A1(W13298), .A2(W24771), .ZN(O11583));
  NOR2X1 G3200 (.A1(W3113), .A2(W3617), .ZN(W22130));
  NOR2X1 G3201 (.A1(W38482), .A2(W29959), .ZN(W41383));
  NOR2X1 G3202 (.A1(W36362), .A2(W17784), .ZN(O11561));
  NOR2X1 G3203 (.A1(W15271), .A2(W12954), .ZN(W28645));
  NOR2X1 G3204 (.A1(I1882), .A2(W3129), .ZN(W9545));
  NOR2X1 G3205 (.A1(W8730), .A2(W556), .ZN(W9544));
  NOR2X1 G3206 (.A1(W9039), .A2(W5970), .ZN(W9543));
  NOR2X1 G3207 (.A1(W3637), .A2(W3688), .ZN(O298));
  NOR2X1 G3208 (.A1(W13883), .A2(W9131), .ZN(O11563));
  NOR2X1 G3209 (.A1(W4493), .A2(W9351), .ZN(W9428));
  NOR2X1 G3210 (.A1(W16540), .A2(W15639), .ZN(O4567));
  NOR2X1 G3211 (.A1(W5706), .A2(I294), .ZN(W9538));
  NOR2X1 G3212 (.A1(W4728), .A2(W2750), .ZN(W9536));
  NOR2X1 G3213 (.A1(W6238), .A2(W1945), .ZN(W9535));
  NOR2X1 G3214 (.A1(W12587), .A2(W33564), .ZN(O11566));
  NOR2X1 G3215 (.A1(W36931), .A2(W24632), .ZN(W41391));
  NOR2X1 G3216 (.A1(W17000), .A2(W12658), .ZN(O4566));
  NOR2X1 G3217 (.A1(W6681), .A2(W4499), .ZN(W9316));
  NOR2X1 G3218 (.A1(W16594), .A2(W22099), .ZN(W41612));
  NOR2X1 G3219 (.A1(W7919), .A2(W2168), .ZN(O282));
  NOR2X1 G3220 (.A1(W11295), .A2(W26811), .ZN(W41613));
  NOR2X1 G3221 (.A1(W134), .A2(W7392), .ZN(W9322));
  NOR2X1 G3222 (.A1(W3964), .A2(I28), .ZN(W9320));
  NOR2X1 G3223 (.A1(W4870), .A2(I1135), .ZN(W9319));
  NOR2X1 G3224 (.A1(W31197), .A2(W10428), .ZN(O11735));
  NOR2X1 G3225 (.A1(W20522), .A2(I378), .ZN(O11737));
  NOR2X1 G3226 (.A1(I1056), .A2(W1316), .ZN(O2449));
  NOR2X1 G3227 (.A1(W5285), .A2(W444), .ZN(W9315));
  NOR2X1 G3228 (.A1(W2812), .A2(W8295), .ZN(W9314));
  NOR2X1 G3229 (.A1(I1072), .A2(W18867), .ZN(O11738));
  NOR2X1 G3230 (.A1(W1484), .A2(W2787), .ZN(W9312));
  NOR2X1 G3231 (.A1(W1933), .A2(W4696), .ZN(O11739));
  NOR2X1 G3232 (.A1(W1191), .A2(W8294), .ZN(W9310));
  NOR2X1 G3233 (.A1(W3109), .A2(W6741), .ZN(O281));
  NOR2X1 G3234 (.A1(W38111), .A2(W22320), .ZN(O11742));
  NOR2X1 G3235 (.A1(W7294), .A2(W2853), .ZN(W9334));
  NOR2X1 G3236 (.A1(W32279), .A2(W20599), .ZN(O11714));
  NOR2X1 G3237 (.A1(W1867), .A2(I1087), .ZN(O11715));
  NOR2X1 G3238 (.A1(W825), .A2(W2137), .ZN(W9340));
  NOR2X1 G3239 (.A1(W18915), .A2(W13020), .ZN(W28557));
  NOR2X1 G3240 (.A1(W6665), .A2(W8364), .ZN(W22205));
  NOR2X1 G3241 (.A1(W25859), .A2(W3484), .ZN(O11720));
  NOR2X1 G3242 (.A1(W28206), .A2(W14167), .ZN(W28556));
  NOR2X1 G3243 (.A1(W17288), .A2(W6352), .ZN(O4539));
  NOR2X1 G3244 (.A1(I1250), .A2(I1008), .ZN(O280));
  NOR2X1 G3245 (.A1(I1380), .A2(W6445), .ZN(O11725));
  NOR2X1 G3246 (.A1(W7679), .A2(W1757), .ZN(W9332));
  NOR2X1 G3247 (.A1(W21766), .A2(W25090), .ZN(O11726));
  NOR2X1 G3248 (.A1(W8605), .A2(W16065), .ZN(O11727));
  NOR2X1 G3249 (.A1(W18352), .A2(W9608), .ZN(O2447));
  NOR2X1 G3250 (.A1(W20172), .A2(W19201), .ZN(O2448));
  NOR2X1 G3251 (.A1(W30341), .A2(W24045), .ZN(O11730));
  NOR2X1 G3252 (.A1(W21550), .A2(W12945), .ZN(W28534));
  NOR2X1 G3253 (.A1(W1715), .A2(W2292), .ZN(W9284));
  NOR2X1 G3254 (.A1(W19329), .A2(W1599), .ZN(O2451));
  NOR2X1 G3255 (.A1(W2749), .A2(W5253), .ZN(O279));
  NOR2X1 G3256 (.A1(W7795), .A2(W7826), .ZN(W9279));
  NOR2X1 G3257 (.A1(W5911), .A2(W5872), .ZN(W9278));
  NOR2X1 G3258 (.A1(W5392), .A2(W1112), .ZN(O2453));
  NOR2X1 G3259 (.A1(W16146), .A2(W7963), .ZN(O11762));
  NOR2X1 G3260 (.A1(W9377), .A2(W35377), .ZN(W41653));
  NOR2X1 G3261 (.A1(W23168), .A2(W35655), .ZN(W41645));
  NOR2X1 G3262 (.A1(I678), .A2(W10862), .ZN(O4532));
  NOR2X1 G3263 (.A1(W2416), .A2(W8497), .ZN(W9272));
  NOR2X1 G3264 (.A1(W8813), .A2(I740), .ZN(W9271));
  NOR2X1 G3265 (.A1(W1612), .A2(W31009), .ZN(O11765));
  NOR2X1 G3266 (.A1(W9914), .A2(W10739), .ZN(W28532));
  NOR2X1 G3267 (.A1(W6085), .A2(W2762), .ZN(W9268));
  NOR2X1 G3268 (.A1(W7959), .A2(W39015), .ZN(O11768));
  NOR2X1 G3269 (.A1(W2789), .A2(W8782), .ZN(W22229));
  NOR2X1 G3270 (.A1(W15356), .A2(W26394), .ZN(W28542));
  NOR2X1 G3271 (.A1(W21475), .A2(W2297), .ZN(W28546));
  NOR2X1 G3272 (.A1(W37889), .A2(W28359), .ZN(O11745));
  NOR2X1 G3273 (.A1(W22184), .A2(W10282), .ZN(O2450));
  NOR2X1 G3274 (.A1(W978), .A2(W12391), .ZN(W22217));
  NOR2X1 G3275 (.A1(W6810), .A2(W6803), .ZN(W9299));
  NOR2X1 G3276 (.A1(W3086), .A2(W6467), .ZN(W9298));
  NOR2X1 G3277 (.A1(W8738), .A2(W28492), .ZN(O11751));
  NOR2X1 G3278 (.A1(W8559), .A2(W7029), .ZN(W9296));
  NOR2X1 G3279 (.A1(W21234), .A2(W19144), .ZN(W22202));
  NOR2X1 G3280 (.A1(W24842), .A2(W1875), .ZN(W41637));
  NOR2X1 G3281 (.A1(W6728), .A2(W6711), .ZN(W9293));
  NOR2X1 G3282 (.A1(I1489), .A2(W6718), .ZN(W9292));
  NOR2X1 G3283 (.A1(W41526), .A2(W27336), .ZN(O11753));
  NOR2X1 G3284 (.A1(W8633), .A2(W2746), .ZN(W9289));
  NOR2X1 G3285 (.A1(W19580), .A2(W17593), .ZN(O11756));
  NOR2X1 G3286 (.A1(W38923), .A2(W22103), .ZN(O11758));
  NOR2X1 G3287 (.A1(W15606), .A2(W23070), .ZN(O4551));
  NOR2X1 G3288 (.A1(W29499), .A2(W21541), .ZN(O11666));
  NOR2X1 G3289 (.A1(W6563), .A2(W1964), .ZN(W9406));
  NOR2X1 G3290 (.A1(W31372), .A2(W26777), .ZN(O11667));
  NOR2X1 G3291 (.A1(W36881), .A2(W12903), .ZN(O11668));
  NOR2X1 G3292 (.A1(I488), .A2(W37403), .ZN(W41531));
  NOR2X1 G3293 (.A1(W1676), .A2(W1997), .ZN(W9402));
  NOR2X1 G3294 (.A1(W31994), .A2(W27596), .ZN(W41532));
  NOR2X1 G3295 (.A1(W689), .A2(W27121), .ZN(W28591));
  NOR2X1 G3296 (.A1(W32608), .A2(W40039), .ZN(O11665));
  NOR2X1 G3297 (.A1(W19804), .A2(W33447), .ZN(O11673));
  NOR2X1 G3298 (.A1(W2369), .A2(W3706), .ZN(W9397));
  NOR2X1 G3299 (.A1(W961), .A2(I570), .ZN(W9396));
  NOR2X1 G3300 (.A1(W29262), .A2(W4333), .ZN(O11674));
  NOR2X1 G3301 (.A1(W10009), .A2(W20040), .ZN(W41539));
  NOR2X1 G3302 (.A1(W2285), .A2(W17241), .ZN(O11677));
  NOR2X1 G3303 (.A1(W6835), .A2(W1636), .ZN(O286));
  NOR2X1 G3304 (.A1(W31576), .A2(W37383), .ZN(O11678));
  NOR2X1 G3305 (.A1(W34227), .A2(W8260), .ZN(W41514));
  NOR2X1 G3306 (.A1(W1162), .A2(I1373), .ZN(W9427));
  NOR2X1 G3307 (.A1(W19233), .A2(I305), .ZN(O11650));
  NOR2X1 G3308 (.A1(W7249), .A2(W5036), .ZN(W9425));
  NOR2X1 G3309 (.A1(W29989), .A2(W12976), .ZN(W41506));
  NOR2X1 G3310 (.A1(W5741), .A2(W6467), .ZN(W9423));
  NOR2X1 G3311 (.A1(W40950), .A2(W12394), .ZN(O11653));
  NOR2X1 G3312 (.A1(W7233), .A2(W6769), .ZN(W9420));
  NOR2X1 G3313 (.A1(W14136), .A2(W33377), .ZN(O11654));
  NOR2X1 G3314 (.A1(I1354), .A2(I1442), .ZN(W9390));
  NOR2X1 G3315 (.A1(W19657), .A2(W14688), .ZN(W28595));
  NOR2X1 G3316 (.A1(W35409), .A2(W33185), .ZN(O11659));
  NOR2X1 G3317 (.A1(W21823), .A2(W3688), .ZN(O11660));
  NOR2X1 G3318 (.A1(W2770), .A2(W1615), .ZN(W9413));
  NOR2X1 G3319 (.A1(W18922), .A2(W15698), .ZN(W22178));
  NOR2X1 G3320 (.A1(W2132), .A2(W36747), .ZN(O11663));
  NOR2X1 G3321 (.A1(W1106), .A2(W18715), .ZN(O4553));
  NOR2X1 G3322 (.A1(W3655), .A2(W13063), .ZN(W28569));
  NOR2X1 G3323 (.A1(W40785), .A2(W29628), .ZN(W41561));
  NOR2X1 G3324 (.A1(W19485), .A2(W22354), .ZN(O11695));
  NOR2X1 G3325 (.A1(W10023), .A2(W544), .ZN(O11698));
  NOR2X1 G3326 (.A1(W16146), .A2(W36703), .ZN(W41568));
  NOR2X1 G3327 (.A1(W4709), .A2(W4373), .ZN(W9363));
  NOR2X1 G3328 (.A1(W37783), .A2(W19082), .ZN(O11699));
  NOR2X1 G3329 (.A1(I1255), .A2(W7563), .ZN(W9361));
  NOR2X1 G3330 (.A1(W30895), .A2(W41095), .ZN(O11701));
  NOR2X1 G3331 (.A1(W37145), .A2(W3888), .ZN(O11692));
  NOR2X1 G3332 (.A1(W14667), .A2(W27647), .ZN(O11704));
  NOR2X1 G3333 (.A1(W14871), .A2(W27354), .ZN(W28565));
  NOR2X1 G3334 (.A1(W4562), .A2(W1414), .ZN(W9352));
  NOR2X1 G3335 (.A1(W540), .A2(W21183), .ZN(O4543));
  NOR2X1 G3336 (.A1(W9311), .A2(W10850), .ZN(O4542));
  NOR2X1 G3337 (.A1(W21287), .A2(W564), .ZN(O11709));
  NOR2X1 G3338 (.A1(W3518), .A2(W17372), .ZN(W22201));
  NOR2X1 G3339 (.A1(W6329), .A2(I38), .ZN(W9378));
  NOR2X1 G3340 (.A1(W3131), .A2(W34841), .ZN(W41545));
  NOR2X1 G3341 (.A1(W9371), .A2(W1619), .ZN(W41548));
  NOR2X1 G3342 (.A1(W6197), .A2(W8070), .ZN(W9384));
  NOR2X1 G3343 (.A1(W9234), .A2(W23018), .ZN(W28584));
  NOR2X1 G3344 (.A1(W39485), .A2(W7784), .ZN(O11684));
  NOR2X1 G3345 (.A1(W7403), .A2(W8624), .ZN(W9381));
  NOR2X1 G3346 (.A1(W3501), .A2(W4050), .ZN(W9380));
  NOR2X1 G3347 (.A1(W8388), .A2(W4341), .ZN(W9379));
  NOR2X1 G3348 (.A1(I1021), .A2(I1650), .ZN(W10216));
  NOR2X1 G3349 (.A1(W17392), .A2(W23677), .ZN(O11685));
  NOR2X1 G3350 (.A1(W3641), .A2(I1599), .ZN(W9376));
  NOR2X1 G3351 (.A1(W27124), .A2(W14542), .ZN(O4549));
  NOR2X1 G3352 (.A1(W6675), .A2(W3415), .ZN(W9374));
  NOR2X1 G3353 (.A1(W12241), .A2(W7277), .ZN(O11689));
  NOR2X1 G3354 (.A1(W1175), .A2(W14947), .ZN(O4548));
  NOR2X1 G3355 (.A1(W12252), .A2(W27126), .ZN(O11691));
  NOR2X1 G3356 (.A1(W4745), .A2(W1592), .ZN(W29129));
  NOR2X1 G3357 (.A1(W2929), .A2(W8347), .ZN(W11068));
  NOR2X1 G3358 (.A1(W6496), .A2(W11319), .ZN(W21663));
  NOR2X1 G3359 (.A1(W269), .A2(W1570), .ZN(W39800));
  NOR2X1 G3360 (.A1(W223), .A2(W30338), .ZN(O10457));
  NOR2X1 G3361 (.A1(W134), .A2(W4694), .ZN(W11064));
  NOR2X1 G3362 (.A1(W39256), .A2(W15346), .ZN(O10459));
  NOR2X1 G3363 (.A1(W1179), .A2(I1190), .ZN(W11062));
  NOR2X1 G3364 (.A1(W8718), .A2(W927), .ZN(W11061));
  NOR2X1 G3365 (.A1(W8823), .A2(W943), .ZN(W11069));
  NOR2X1 G3366 (.A1(W13692), .A2(W13800), .ZN(O10462));
  NOR2X1 G3367 (.A1(W21475), .A2(W7722), .ZN(W21665));
  NOR2X1 G3368 (.A1(I711), .A2(W1881), .ZN(W11057));
  NOR2X1 G3369 (.A1(W3949), .A2(I912), .ZN(W11056));
  NOR2X1 G3370 (.A1(W12653), .A2(W25294), .ZN(W29126));
  NOR2X1 G3371 (.A1(W3972), .A2(W3899), .ZN(W11053));
  NOR2X1 G3372 (.A1(W2108), .A2(W27096), .ZN(W39812));
  NOR2X1 G3373 (.A1(W5772), .A2(W3682), .ZN(W11051));
  NOR2X1 G3374 (.A1(W2982), .A2(W3589), .ZN(W11077));
  NOR2X1 G3375 (.A1(W10517), .A2(W8667), .ZN(O479));
  NOR2X1 G3376 (.A1(W10744), .A2(W7872), .ZN(W11085));
  NOR2X1 G3377 (.A1(W4094), .A2(W24530), .ZN(O10449));
  NOR2X1 G3378 (.A1(W3374), .A2(W6593), .ZN(W11083));
  NOR2X1 G3379 (.A1(W7881), .A2(W7121), .ZN(W11082));
  NOR2X1 G3380 (.A1(W10929), .A2(W7887), .ZN(O478));
  NOR2X1 G3381 (.A1(W13493), .A2(W28651), .ZN(W39791));
  NOR2X1 G3382 (.A1(W1164), .A2(W15645), .ZN(W21661));
  NOR2X1 G3383 (.A1(W4500), .A2(W4513), .ZN(O474));
  NOR2X1 G3384 (.A1(W4184), .A2(W5874), .ZN(W11076));
  NOR2X1 G3385 (.A1(W39417), .A2(W30843), .ZN(O10451));
  NOR2X1 G3386 (.A1(W7499), .A2(I112), .ZN(W11074));
  NOR2X1 G3387 (.A1(I695), .A2(W15715), .ZN(O10452));
  NOR2X1 G3388 (.A1(I578), .A2(W137), .ZN(W11072));
  NOR2X1 G3389 (.A1(W22807), .A2(W19777), .ZN(O4760));
  NOR2X1 G3390 (.A1(I1575), .A2(W10131), .ZN(W11070));
  NOR2X1 G3391 (.A1(I1392), .A2(W2562), .ZN(O4756));
  NOR2X1 G3392 (.A1(W705), .A2(I271), .ZN(O470));
  NOR2X1 G3393 (.A1(W18045), .A2(W27554), .ZN(O10480));
  NOR2X1 G3394 (.A1(W23911), .A2(W5934), .ZN(O10481));
  NOR2X1 G3395 (.A1(W25479), .A2(W36862), .ZN(O10483));
  NOR2X1 G3396 (.A1(W2184), .A2(W1403), .ZN(W11024));
  NOR2X1 G3397 (.A1(W9262), .A2(W14638), .ZN(O10485));
  NOR2X1 G3398 (.A1(W12332), .A2(W36277), .ZN(O10486));
  NOR2X1 G3399 (.A1(W5898), .A2(W38049), .ZN(O10489));
  NOR2X1 G3400 (.A1(W24090), .A2(W19282), .ZN(O10479));
  NOR2X1 G3401 (.A1(W18916), .A2(W27157), .ZN(O10490));
  NOR2X1 G3402 (.A1(W5233), .A2(W10264), .ZN(W11018));
  NOR2X1 G3403 (.A1(W10824), .A2(W3447), .ZN(O467));
  NOR2X1 G3404 (.A1(W38320), .A2(W12059), .ZN(O10491));
  NOR2X1 G3405 (.A1(W1033), .A2(W863), .ZN(O4755));
  NOR2X1 G3406 (.A1(W8028), .A2(W9342), .ZN(O466));
  NOR2X1 G3407 (.A1(W4126), .A2(W3974), .ZN(O2306));
  NOR2X1 G3408 (.A1(W26026), .A2(W20399), .ZN(W39849));
  NOR2X1 G3409 (.A1(W12812), .A2(W18991), .ZN(W21672));
  NOR2X1 G3410 (.A1(W8640), .A2(I844), .ZN(W11048));
  NOR2X1 G3411 (.A1(W7450), .A2(I371), .ZN(W21669));
  NOR2X1 G3412 (.A1(W19588), .A2(W32920), .ZN(O10468));
  NOR2X1 G3413 (.A1(W2785), .A2(W3711), .ZN(W11045));
  NOR2X1 G3414 (.A1(W1393), .A2(W7624), .ZN(W11044));
  NOR2X1 G3415 (.A1(W21144), .A2(W8817), .ZN(W39816));
  NOR2X1 G3416 (.A1(W20437), .A2(I1262), .ZN(W21670));
  NOR2X1 G3417 (.A1(W20856), .A2(I945), .ZN(W29124));
  NOR2X1 G3418 (.A1(W10686), .A2(I1121), .ZN(O2304));
  NOR2X1 G3419 (.A1(W3148), .A2(W35909), .ZN(O10473));
  NOR2X1 G3420 (.A1(W7519), .A2(W990), .ZN(W11038));
  NOR2X1 G3421 (.A1(W1602), .A2(W1785), .ZN(W11035));
  NOR2X1 G3422 (.A1(W2166), .A2(W58), .ZN(W11034));
  NOR2X1 G3423 (.A1(W6250), .A2(W8450), .ZN(O10476));
  NOR2X1 G3424 (.A1(W27292), .A2(W37111), .ZN(O10477));
  NOR2X1 G3425 (.A1(W37073), .A2(W9135), .ZN(O10478));
  NOR2X1 G3426 (.A1(W15204), .A2(W2889), .ZN(W21642));
  NOR2X1 G3427 (.A1(W10757), .A2(I103), .ZN(W11141));
  NOR2X1 G3428 (.A1(W13280), .A2(W8189), .ZN(O10403));
  NOR2X1 G3429 (.A1(W9209), .A2(W3014), .ZN(W11139));
  NOR2X1 G3430 (.A1(W22383), .A2(W16946), .ZN(W39723));
  NOR2X1 G3431 (.A1(W16917), .A2(W2878), .ZN(W29154));
  NOR2X1 G3432 (.A1(W18166), .A2(W9811), .ZN(W21639));
  NOR2X1 G3433 (.A1(W11857), .A2(W19446), .ZN(W29152));
  NOR2X1 G3434 (.A1(W979), .A2(W1218), .ZN(W21641));
  NOR2X1 G3435 (.A1(I1084), .A2(W2218), .ZN(W11143));
  NOR2X1 G3436 (.A1(W5692), .A2(W7507), .ZN(W11132));
  NOR2X1 G3437 (.A1(W3080), .A2(W8602), .ZN(O10413));
  NOR2X1 G3438 (.A1(W4713), .A2(W27083), .ZN(W29150));
  NOR2X1 G3439 (.A1(W1979), .A2(I495), .ZN(W11129));
  NOR2X1 G3440 (.A1(I1981), .A2(I1979), .ZN(W11128));
  NOR2X1 G3441 (.A1(W34891), .A2(W27959), .ZN(O10417));
  NOR2X1 G3442 (.A1(W4783), .A2(I1602), .ZN(O4767));
  NOR2X1 G3443 (.A1(I1168), .A2(W6658), .ZN(O4766));
  NOR2X1 G3444 (.A1(W18981), .A2(W17822), .ZN(O10394));
  NOR2X1 G3445 (.A1(W2198), .A2(W6460), .ZN(W11160));
  NOR2X1 G3446 (.A1(W38349), .A2(W2489), .ZN(O10390));
  NOR2X1 G3447 (.A1(W15322), .A2(W7236), .ZN(O10391));
  NOR2X1 G3448 (.A1(W1896), .A2(W1211), .ZN(W11157));
  NOR2X1 G3449 (.A1(W5670), .A2(W6513), .ZN(W11156));
  NOR2X1 G3450 (.A1(I1611), .A2(W10759), .ZN(O10392));
  NOR2X1 G3451 (.A1(W5189), .A2(W15830), .ZN(O4771));
  NOR2X1 G3452 (.A1(I726), .A2(W10413), .ZN(W11153));
  NOR2X1 G3453 (.A1(W4446), .A2(W10491), .ZN(O10420));
  NOR2X1 G3454 (.A1(I208), .A2(W2243), .ZN(W11150));
  NOR2X1 G3455 (.A1(W6116), .A2(W7060), .ZN(W11149));
  NOR2X1 G3456 (.A1(W35751), .A2(W30503), .ZN(O10396));
  NOR2X1 G3457 (.A1(W29122), .A2(W25218), .ZN(W39709));
  NOR2X1 G3458 (.A1(W7534), .A2(W20522), .ZN(O4769));
  NOR2X1 G3459 (.A1(W1228), .A2(W15765), .ZN(O2301));
  NOR2X1 G3460 (.A1(W4005), .A2(W13871), .ZN(O10400));
  NOR2X1 G3461 (.A1(W23073), .A2(W36328), .ZN(O10441));
  NOR2X1 G3462 (.A1(W34786), .A2(W14858), .ZN(W39772));
  NOR2X1 G3463 (.A1(W18229), .A2(W21865), .ZN(O4764));
  NOR2X1 G3464 (.A1(W7805), .A2(W4883), .ZN(W21653));
  NOR2X1 G3465 (.A1(W10981), .A2(W1471), .ZN(W11101));
  NOR2X1 G3466 (.A1(W10775), .A2(W10544), .ZN(O481));
  NOR2X1 G3467 (.A1(W5244), .A2(W10218), .ZN(W11099));
  NOR2X1 G3468 (.A1(W19254), .A2(W35530), .ZN(W39775));
  NOR2X1 G3469 (.A1(W7394), .A2(W10207), .ZN(W11097));
  NOR2X1 G3470 (.A1(W8663), .A2(I24), .ZN(W11105));
  NOR2X1 G3471 (.A1(W28921), .A2(W24477), .ZN(O4763));
  NOR2X1 G3472 (.A1(W3685), .A2(W7891), .ZN(W21655));
  NOR2X1 G3473 (.A1(W12746), .A2(W8788), .ZN(W39779));
  NOR2X1 G3474 (.A1(W26300), .A2(W5171), .ZN(O4762));
  NOR2X1 G3475 (.A1(W14457), .A2(W9117), .ZN(O4761));
  NOR2X1 G3476 (.A1(W6621), .A2(W23556), .ZN(W29133));
  NOR2X1 G3477 (.A1(W35815), .A2(W6514), .ZN(O10447));
  NOR2X1 G3478 (.A1(W4539), .A2(W6383), .ZN(W11088));
  NOR2X1 G3479 (.A1(W20511), .A2(W14925), .ZN(O10436));
  NOR2X1 G3480 (.A1(W3309), .A2(W6376), .ZN(W11123));
  NOR2X1 G3481 (.A1(W35604), .A2(W1349), .ZN(O10421));
  NOR2X1 G3482 (.A1(W11135), .A2(W21045), .ZN(W21647));
  NOR2X1 G3483 (.A1(W2640), .A2(W10424), .ZN(W11119));
  NOR2X1 G3484 (.A1(W10244), .A2(W4017), .ZN(W11118));
  NOR2X1 G3485 (.A1(W24984), .A2(W39541), .ZN(O10429));
  NOR2X1 G3486 (.A1(W14106), .A2(W30578), .ZN(O10431));
  NOR2X1 G3487 (.A1(W6407), .A2(W14044), .ZN(W29143));
  NOR2X1 G3488 (.A1(W32923), .A2(W5847), .ZN(O10497));
  NOR2X1 G3489 (.A1(W1763), .A2(W5203), .ZN(W11112));
  NOR2X1 G3490 (.A1(W19196), .A2(I1742), .ZN(W21650));
  NOR2X1 G3491 (.A1(W19530), .A2(W25112), .ZN(W39768));
  NOR2X1 G3492 (.A1(W22065), .A2(W14370), .ZN(W29140));
  NOR2X1 G3493 (.A1(I30), .A2(W18465), .ZN(O10438));
  NOR2X1 G3494 (.A1(W13830), .A2(W19801), .ZN(W39771));
  NOR2X1 G3495 (.A1(I1000), .A2(W5863), .ZN(W11106));
  NOR2X1 G3496 (.A1(W4504), .A2(W1039), .ZN(O452));
  NOR2X1 G3497 (.A1(W480), .A2(W24723), .ZN(O10567));
  NOR2X1 G3498 (.A1(W4475), .A2(W15331), .ZN(W39952));
  NOR2X1 G3499 (.A1(W18168), .A2(W20075), .ZN(W29094));
  NOR2X1 G3500 (.A1(W1257), .A2(W9764), .ZN(W10911));
  NOR2X1 G3501 (.A1(W39772), .A2(W16323), .ZN(O10573));
  NOR2X1 G3502 (.A1(W10245), .A2(W6119), .ZN(W10909));
  NOR2X1 G3503 (.A1(W1147), .A2(W16351), .ZN(O2316));
  NOR2X1 G3504 (.A1(W21104), .A2(W13755), .ZN(W21707));
  NOR2X1 G3505 (.A1(W10398), .A2(W5224), .ZN(W10916));
  NOR2X1 G3506 (.A1(W230), .A2(W7070), .ZN(W10904));
  NOR2X1 G3507 (.A1(W1964), .A2(W8441), .ZN(W10903));
  NOR2X1 G3508 (.A1(W17915), .A2(W10540), .ZN(W39962));
  NOR2X1 G3509 (.A1(W4253), .A2(W39525), .ZN(O10578));
  NOR2X1 G3510 (.A1(W35331), .A2(W11729), .ZN(W39965));
  NOR2X1 G3511 (.A1(W436), .A2(W8942), .ZN(W10899));
  NOR2X1 G3512 (.A1(W9078), .A2(W14146), .ZN(W29092));
  NOR2X1 G3513 (.A1(I1717), .A2(I534), .ZN(W10897));
  NOR2X1 G3514 (.A1(W10577), .A2(I541), .ZN(W10924));
  NOR2X1 G3515 (.A1(W33878), .A2(W24517), .ZN(W39922));
  NOR2X1 G3516 (.A1(W482), .A2(W394), .ZN(W39925));
  NOR2X1 G3517 (.A1(W33574), .A2(W1753), .ZN(O10552));
  NOR2X1 G3518 (.A1(W7027), .A2(W5001), .ZN(W10932));
  NOR2X1 G3519 (.A1(W7374), .A2(I701), .ZN(W10930));
  NOR2X1 G3520 (.A1(W6309), .A2(I32), .ZN(W10929));
  NOR2X1 G3521 (.A1(W9872), .A2(W1267), .ZN(O455));
  NOR2X1 G3522 (.A1(W8483), .A2(W31741), .ZN(O10557));
  NOR2X1 G3523 (.A1(W21081), .A2(I1127), .ZN(W39968));
  NOR2X1 G3524 (.A1(W22858), .A2(W22261), .ZN(O10562));
  NOR2X1 G3525 (.A1(W8586), .A2(W10812), .ZN(W10922));
  NOR2X1 G3526 (.A1(W13310), .A2(I1780), .ZN(O10563));
  NOR2X1 G3527 (.A1(W859), .A2(W13073), .ZN(O2315));
  NOR2X1 G3528 (.A1(W37409), .A2(W29977), .ZN(O10565));
  NOR2X1 G3529 (.A1(W7553), .A2(W7753), .ZN(W29096));
  NOR2X1 G3530 (.A1(W6065), .A2(W22395), .ZN(W39945));
  NOR2X1 G3531 (.A1(W14930), .A2(W20112), .ZN(W21728));
  NOR2X1 G3532 (.A1(W8354), .A2(W3342), .ZN(W10875));
  NOR2X1 G3533 (.A1(I1941), .A2(W10591), .ZN(W39992));
  NOR2X1 G3534 (.A1(W770), .A2(W27111), .ZN(W29078));
  NOR2X1 G3535 (.A1(W11231), .A2(W634), .ZN(O2318));
  NOR2X1 G3536 (.A1(W33190), .A2(W32022), .ZN(O10599));
  NOR2X1 G3537 (.A1(W680), .A2(W5461), .ZN(W10868));
  NOR2X1 G3538 (.A1(W8816), .A2(W8637), .ZN(W10865));
  NOR2X1 G3539 (.A1(W14510), .A2(W20505), .ZN(W29072));
  NOR2X1 G3540 (.A1(W10540), .A2(W9961), .ZN(O4732));
  NOR2X1 G3541 (.A1(W2158), .A2(W6328), .ZN(W10861));
  NOR2X1 G3542 (.A1(W1025), .A2(W21940), .ZN(W40007));
  NOR2X1 G3543 (.A1(W23084), .A2(W13662), .ZN(W29070));
  NOR2X1 G3544 (.A1(W10592), .A2(W2316), .ZN(W29069));
  NOR2X1 G3545 (.A1(W21975), .A2(W38590), .ZN(O10607));
  NOR2X1 G3546 (.A1(W10800), .A2(W35454), .ZN(O10609));
  NOR2X1 G3547 (.A1(W98), .A2(W28849), .ZN(O10610));
  NOR2X1 G3548 (.A1(W8935), .A2(W17038), .ZN(O10612));
  NOR2X1 G3549 (.A1(W9520), .A2(W8005), .ZN(O10587));
  NOR2X1 G3550 (.A1(W19022), .A2(W1036), .ZN(O4740));
  NOR2X1 G3551 (.A1(W12147), .A2(W19291), .ZN(W21711));
  NOR2X1 G3552 (.A1(W10292), .A2(W17053), .ZN(W21712));
  NOR2X1 G3553 (.A1(W4086), .A2(W6430), .ZN(W10892));
  NOR2X1 G3554 (.A1(W12916), .A2(W5539), .ZN(W21713));
  NOR2X1 G3555 (.A1(W16671), .A2(W10256), .ZN(O4739));
  NOR2X1 G3556 (.A1(W15903), .A2(W8896), .ZN(O4738));
  NOR2X1 G3557 (.A1(W16998), .A2(I857), .ZN(O10586));
  NOR2X1 G3558 (.A1(W98), .A2(W4657), .ZN(W10937));
  NOR2X1 G3559 (.A1(W12121), .A2(W5826), .ZN(W39980));
  NOR2X1 G3560 (.A1(W9402), .A2(W7601), .ZN(O10589));
  NOR2X1 G3561 (.A1(W26994), .A2(W12099), .ZN(O10591));
  NOR2X1 G3562 (.A1(W25165), .A2(W15264), .ZN(O10592));
  NOR2X1 G3563 (.A1(W3454), .A2(W3067), .ZN(W10879));
  NOR2X1 G3564 (.A1(W10904), .A2(W38851), .ZN(W39990));
  NOR2X1 G3565 (.A1(W10850), .A2(W8327), .ZN(W10877));
  NOR2X1 G3566 (.A1(W3785), .A2(W38855), .ZN(O10521));
  NOR2X1 G3567 (.A1(W30594), .A2(W21811), .ZN(W39877));
  NOR2X1 G3568 (.A1(W6122), .A2(W8084), .ZN(W10989));
  NOR2X1 G3569 (.A1(W10496), .A2(W23694), .ZN(O10519));
  NOR2X1 G3570 (.A1(W13001), .A2(W21375), .ZN(O2310));
  NOR2X1 G3571 (.A1(I1376), .A2(W7746), .ZN(W10986));
  NOR2X1 G3572 (.A1(W6833), .A2(W6499), .ZN(O460));
  NOR2X1 G3573 (.A1(W7563), .A2(I1120), .ZN(W10984));
  NOR2X1 G3574 (.A1(W12994), .A2(W8808), .ZN(O10520));
  NOR2X1 G3575 (.A1(W8407), .A2(W944), .ZN(W10991));
  NOR2X1 G3576 (.A1(W815), .A2(W2345), .ZN(W10981));
  NOR2X1 G3577 (.A1(W21396), .A2(I706), .ZN(W21687));
  NOR2X1 G3578 (.A1(W7459), .A2(W6957), .ZN(W10979));
  NOR2X1 G3579 (.A1(W3982), .A2(W3774), .ZN(W10978));
  NOR2X1 G3580 (.A1(W38818), .A2(W28027), .ZN(O10524));
  NOR2X1 G3581 (.A1(W6170), .A2(W1627), .ZN(W10976));
  NOR2X1 G3582 (.A1(W2114), .A2(W5697), .ZN(W10975));
  NOR2X1 G3583 (.A1(W11201), .A2(W37072), .ZN(W39887));
  NOR2X1 G3584 (.A1(W38374), .A2(W36073), .ZN(O10512));
  NOR2X1 G3585 (.A1(W4496), .A2(W9526), .ZN(O10499));
  NOR2X1 G3586 (.A1(W18861), .A2(W1485), .ZN(O2307));
  NOR2X1 G3587 (.A1(W5932), .A2(W10892), .ZN(W11008));
  NOR2X1 G3588 (.A1(W10811), .A2(W2624), .ZN(W11006));
  NOR2X1 G3589 (.A1(W5341), .A2(W28892), .ZN(O10504));
  NOR2X1 G3590 (.A1(W39854), .A2(W13576), .ZN(W39864));
  NOR2X1 G3591 (.A1(W8441), .A2(W8715), .ZN(W11002));
  NOR2X1 G3592 (.A1(W16779), .A2(W11435), .ZN(O10511));
  NOR2X1 G3593 (.A1(W25457), .A2(W3924), .ZN(O10526));
  NOR2X1 G3594 (.A1(W1522), .A2(W5940), .ZN(W10999));
  NOR2X1 G3595 (.A1(W11571), .A2(W11388), .ZN(O2309));
  NOR2X1 G3596 (.A1(W2177), .A2(W2963), .ZN(W10996));
  NOR2X1 G3597 (.A1(W16381), .A2(W16991), .ZN(O4754));
  NOR2X1 G3598 (.A1(W7239), .A2(W11947), .ZN(W21685));
  NOR2X1 G3599 (.A1(W13558), .A2(W35923), .ZN(O10518));
  NOR2X1 G3600 (.A1(W3022), .A2(W8823), .ZN(W10992));
  NOR2X1 G3601 (.A1(W8974), .A2(W21037), .ZN(W21695));
  NOR2X1 G3602 (.A1(W7408), .A2(W10166), .ZN(W10955));
  NOR2X1 G3603 (.A1(W2817), .A2(W12106), .ZN(O10534));
  NOR2X1 G3604 (.A1(W4578), .A2(I462), .ZN(O10535));
  NOR2X1 G3605 (.A1(W729), .A2(W18021), .ZN(O10536));
  NOR2X1 G3606 (.A1(W30119), .A2(W4341), .ZN(O10537));
  NOR2X1 G3607 (.A1(W3987), .A2(W9239), .ZN(W10950));
  NOR2X1 G3608 (.A1(W19364), .A2(W30045), .ZN(O10538));
  NOR2X1 G3609 (.A1(W26446), .A2(W2671), .ZN(O4748));
  NOR2X1 G3610 (.A1(W22428), .A2(W2758), .ZN(O10533));
  NOR2X1 G3611 (.A1(W14516), .A2(W6918), .ZN(O10541));
  NOR2X1 G3612 (.A1(I750), .A2(W10411), .ZN(W10945));
  NOR2X1 G3613 (.A1(W27204), .A2(W24921), .ZN(O10546));
  NOR2X1 G3614 (.A1(W10497), .A2(W976), .ZN(W10942));
  NOR2X1 G3615 (.A1(W13842), .A2(W15858), .ZN(O10547));
  NOR2X1 G3616 (.A1(W17384), .A2(W30872), .ZN(O10549));
  NOR2X1 G3617 (.A1(W10580), .A2(W9855), .ZN(W10939));
  NOR2X1 G3618 (.A1(I1462), .A2(W21096), .ZN(W29104));
  NOR2X1 G3619 (.A1(W3237), .A2(W5730), .ZN(W10964));
  NOR2X1 G3620 (.A1(W32151), .A2(W28685), .ZN(W39889));
  NOR2X1 G3621 (.A1(W2652), .A2(W7180), .ZN(O10527));
  NOR2X1 G3622 (.A1(W10581), .A2(W15149), .ZN(O4753));
  NOR2X1 G3623 (.A1(W8523), .A2(W13741), .ZN(O4752));
  NOR2X1 G3624 (.A1(I543), .A2(W4850), .ZN(W21690));
  NOR2X1 G3625 (.A1(W2062), .A2(W9385), .ZN(W10967));
  NOR2X1 G3626 (.A1(W5704), .A2(W6141), .ZN(W10966));
  NOR2X1 G3627 (.A1(W8839), .A2(W8091), .ZN(W10965));
  NOR2X1 G3628 (.A1(W5300), .A2(W4322), .ZN(W11161));
  NOR2X1 G3629 (.A1(W6630), .A2(W8620), .ZN(O456));
  NOR2X1 G3630 (.A1(W21048), .A2(W19331), .ZN(W21691));
  NOR2X1 G3631 (.A1(W16805), .A2(W7748), .ZN(O2311));
  NOR2X1 G3632 (.A1(W7466), .A2(W26701), .ZN(O4751));
  NOR2X1 G3633 (.A1(W37186), .A2(W22242), .ZN(O10532));
  NOR2X1 G3634 (.A1(I72), .A2(W10091), .ZN(W10958));
  NOR2X1 G3635 (.A1(I1148), .A2(I1006), .ZN(W10957));
  NOR2X1 G3636 (.A1(W30543), .A2(W8173), .ZN(O10257));
  NOR2X1 G3637 (.A1(W8529), .A2(W9185), .ZN(W11368));
  NOR2X1 G3638 (.A1(W11075), .A2(W937), .ZN(O10248));
  NOR2X1 G3639 (.A1(W925), .A2(W11342), .ZN(O10253));
  NOR2X1 G3640 (.A1(W5694), .A2(W5762), .ZN(W11364));
  NOR2X1 G3641 (.A1(W18556), .A2(W7690), .ZN(W39502));
  NOR2X1 G3642 (.A1(W32338), .A2(W12023), .ZN(O10255));
  NOR2X1 G3643 (.A1(W8935), .A2(W18468), .ZN(W39507));
  NOR2X1 G3644 (.A1(W5257), .A2(W2252), .ZN(W11359));
  NOR2X1 G3645 (.A1(W10178), .A2(W22267), .ZN(O10246));
  NOR2X1 G3646 (.A1(W4405), .A2(W9821), .ZN(W11357));
  NOR2X1 G3647 (.A1(W8721), .A2(I1751), .ZN(W11356));
  NOR2X1 G3648 (.A1(W8322), .A2(W7574), .ZN(W11355));
  NOR2X1 G3649 (.A1(W9918), .A2(W5176), .ZN(W11354));
  NOR2X1 G3650 (.A1(W13094), .A2(W17922), .ZN(O4789));
  NOR2X1 G3651 (.A1(W38703), .A2(W24811), .ZN(O10259));
  NOR2X1 G3652 (.A1(W2875), .A2(W410), .ZN(W21572));
  NOR2X1 G3653 (.A1(W687), .A2(W438), .ZN(W11350));
  NOR2X1 G3654 (.A1(W2532), .A2(W7321), .ZN(W11378));
  NOR2X1 G3655 (.A1(W222), .A2(W3159), .ZN(W21561));
  NOR2X1 G3656 (.A1(W5568), .A2(W5341), .ZN(W11386));
  NOR2X1 G3657 (.A1(W13762), .A2(W2967), .ZN(W21562));
  NOR2X1 G3658 (.A1(W8727), .A2(I508), .ZN(W39480));
  NOR2X1 G3659 (.A1(W11920), .A2(W7725), .ZN(W21563));
  NOR2X1 G3660 (.A1(W2191), .A2(W5312), .ZN(W11382));
  NOR2X1 G3661 (.A1(W6718), .A2(W13728), .ZN(W21564));
  NOR2X1 G3662 (.A1(W1434), .A2(W6748), .ZN(W11380));
  NOR2X1 G3663 (.A1(W18775), .A2(W1811), .ZN(W29205));
  NOR2X1 G3664 (.A1(W19210), .A2(W7931), .ZN(W21566));
  NOR2X1 G3665 (.A1(W5238), .A2(W2337), .ZN(O503));
  NOR2X1 G3666 (.A1(W32420), .A2(W37426), .ZN(W39485));
  NOR2X1 G3667 (.A1(W1912), .A2(W38913), .ZN(O10242));
  NOR2X1 G3668 (.A1(W897), .A2(W8666), .ZN(W11372));
  NOR2X1 G3669 (.A1(W22235), .A2(W3892), .ZN(W39489));
  NOR2X1 G3670 (.A1(W27094), .A2(W26361), .ZN(W29209));
  NOR2X1 G3671 (.A1(W21017), .A2(I1806), .ZN(W21581));
  NOR2X1 G3672 (.A1(W2931), .A2(W10208), .ZN(W11330));
  NOR2X1 G3673 (.A1(W2901), .A2(W5743), .ZN(W21578));
  NOR2X1 G3674 (.A1(W22519), .A2(W11262), .ZN(W29202));
  NOR2X1 G3675 (.A1(W13530), .A2(W28494), .ZN(O10280));
  NOR2X1 G3676 (.A1(W11092), .A2(W6164), .ZN(W39541));
  NOR2X1 G3677 (.A1(W6648), .A2(W9520), .ZN(W11325));
  NOR2X1 G3678 (.A1(W11663), .A2(W21265), .ZN(O10282));
  NOR2X1 G3679 (.A1(W20141), .A2(W22174), .ZN(O10284));
  NOR2X1 G3680 (.A1(W6174), .A2(I1710), .ZN(W11331));
  NOR2X1 G3681 (.A1(I1859), .A2(W13357), .ZN(W29198));
  NOR2X1 G3682 (.A1(W3740), .A2(W1124), .ZN(W11319));
  NOR2X1 G3683 (.A1(W11698), .A2(W21605), .ZN(O4786));
  NOR2X1 G3684 (.A1(W27206), .A2(W12257), .ZN(W29196));
  NOR2X1 G3685 (.A1(I1396), .A2(W2311), .ZN(W11316));
  NOR2X1 G3686 (.A1(W3828), .A2(W2255), .ZN(W21585));
  NOR2X1 G3687 (.A1(W5448), .A2(W23408), .ZN(W39556));
  NOR2X1 G3688 (.A1(W35207), .A2(W26185), .ZN(O10290));
  NOR2X1 G3689 (.A1(W36198), .A2(W3492), .ZN(O10270));
  NOR2X1 G3690 (.A1(W9834), .A2(W7620), .ZN(W11348));
  NOR2X1 G3691 (.A1(W36708), .A2(W13829), .ZN(W39516));
  NOR2X1 G3692 (.A1(W9834), .A2(W3207), .ZN(W21574));
  NOR2X1 G3693 (.A1(W25531), .A2(W18093), .ZN(O4788));
  NOR2X1 G3694 (.A1(W415), .A2(W1616), .ZN(O501));
  NOR2X1 G3695 (.A1(W6484), .A2(W2268), .ZN(O10265));
  NOR2X1 G3696 (.A1(W4748), .A2(W9753), .ZN(W11342));
  NOR2X1 G3697 (.A1(W10267), .A2(W24063), .ZN(O10267));
  NOR2X1 G3698 (.A1(W27977), .A2(W37941), .ZN(O10234));
  NOR2X1 G3699 (.A1(W10477), .A2(W36813), .ZN(W39527));
  NOR2X1 G3700 (.A1(W10379), .A2(W16998), .ZN(O2285));
  NOR2X1 G3701 (.A1(W18883), .A2(W27759), .ZN(W39530));
  NOR2X1 G3702 (.A1(W3044), .A2(W32359), .ZN(O10272));
  NOR2X1 G3703 (.A1(W27573), .A2(W14259), .ZN(O10273));
  NOR2X1 G3704 (.A1(W2855), .A2(W5247), .ZN(W11333));
  NOR2X1 G3705 (.A1(W29239), .A2(W20440), .ZN(O10276));
  NOR2X1 G3706 (.A1(W7307), .A2(W7742), .ZN(O509));
  NOR2X1 G3707 (.A1(W13543), .A2(W28834), .ZN(W39408));
  NOR2X1 G3708 (.A1(W21925), .A2(W3263), .ZN(O4797));
  NOR2X1 G3709 (.A1(W21660), .A2(W27978), .ZN(O4796));
  NOR2X1 G3710 (.A1(W1517), .A2(W10106), .ZN(W11439));
  NOR2X1 G3711 (.A1(W17553), .A2(W5487), .ZN(O4795));
  NOR2X1 G3712 (.A1(W15147), .A2(I508), .ZN(O10193));
  NOR2X1 G3713 (.A1(W33035), .A2(W39285), .ZN(O10194));
  NOR2X1 G3714 (.A1(W11716), .A2(W22900), .ZN(W29227));
  NOR2X1 G3715 (.A1(W24378), .A2(W36502), .ZN(O10185));
  NOR2X1 G3716 (.A1(W6386), .A2(W9548), .ZN(W11433));
  NOR2X1 G3717 (.A1(W18456), .A2(W22702), .ZN(W39420));
  NOR2X1 G3718 (.A1(W484), .A2(W1440), .ZN(W11431));
  NOR2X1 G3719 (.A1(W7880), .A2(W2606), .ZN(W11430));
  NOR2X1 G3720 (.A1(W21818), .A2(W1966), .ZN(W39424));
  NOR2X1 G3721 (.A1(W24190), .A2(W12764), .ZN(O10199));
  NOR2X1 G3722 (.A1(W37873), .A2(I223), .ZN(O10200));
  NOR2X1 G3723 (.A1(W30970), .A2(W19620), .ZN(O10204));
  NOR2X1 G3724 (.A1(W1521), .A2(W8080), .ZN(W11453));
  NOR2X1 G3725 (.A1(W4220), .A2(W1825), .ZN(W11463));
  NOR2X1 G3726 (.A1(W3598), .A2(W9781), .ZN(O10171));
  NOR2X1 G3727 (.A1(W215), .A2(W6998), .ZN(W11461));
  NOR2X1 G3728 (.A1(W3101), .A2(W10645), .ZN(W11460));
  NOR2X1 G3729 (.A1(W9356), .A2(W1567), .ZN(W11458));
  NOR2X1 G3730 (.A1(W15550), .A2(W24516), .ZN(O10175));
  NOR2X1 G3731 (.A1(W19574), .A2(W36148), .ZN(O10177));
  NOR2X1 G3732 (.A1(W3464), .A2(W11994), .ZN(W39394));
  NOR2X1 G3733 (.A1(W24482), .A2(W28503), .ZN(O10205));
  NOR2X1 G3734 (.A1(W27534), .A2(W23414), .ZN(O10180));
  NOR2X1 G3735 (.A1(W28637), .A2(W2413), .ZN(O10181));
  NOR2X1 G3736 (.A1(W4963), .A2(W3922), .ZN(W11450));
  NOR2X1 G3737 (.A1(W14199), .A2(W34144), .ZN(O10183));
  NOR2X1 G3738 (.A1(W619), .A2(W17688), .ZN(O4800));
  NOR2X1 G3739 (.A1(W195), .A2(W6163), .ZN(W11447));
  NOR2X1 G3740 (.A1(W5227), .A2(W36180), .ZN(O10184));
  NOR2X1 G3741 (.A1(W15603), .A2(W3384), .ZN(W21556));
  NOR2X1 G3742 (.A1(W30612), .A2(I1860), .ZN(O10218));
  NOR2X1 G3743 (.A1(W3008), .A2(W11163), .ZN(W11405));
  NOR2X1 G3744 (.A1(W6785), .A2(W519), .ZN(O10219));
  NOR2X1 G3745 (.A1(W21230), .A2(W20737), .ZN(W39454));
  NOR2X1 G3746 (.A1(W15152), .A2(W26537), .ZN(W39456));
  NOR2X1 G3747 (.A1(I316), .A2(W7824), .ZN(O4792));
  NOR2X1 G3748 (.A1(W27732), .A2(W7323), .ZN(O10223));
  NOR2X1 G3749 (.A1(W19294), .A2(W22041), .ZN(W29218));
  NOR2X1 G3750 (.A1(W28890), .A2(W2243), .ZN(W39450));
  NOR2X1 G3751 (.A1(W8437), .A2(W30282), .ZN(W39466));
  NOR2X1 G3752 (.A1(W20159), .A2(W28785), .ZN(W29217));
  NOR2X1 G3753 (.A1(W6901), .A2(W3455), .ZN(W21558));
  NOR2X1 G3754 (.A1(W33846), .A2(W28638), .ZN(O10230));
  NOR2X1 G3755 (.A1(W6946), .A2(W3729), .ZN(W11393));
  NOR2X1 G3756 (.A1(W10293), .A2(W19407), .ZN(O10231));
  NOR2X1 G3757 (.A1(I928), .A2(W1729), .ZN(W21559));
  NOR2X1 G3758 (.A1(W16221), .A2(W30724), .ZN(O10233));
  NOR2X1 G3759 (.A1(W3602), .A2(W5186), .ZN(W29220));
  NOR2X1 G3760 (.A1(W6885), .A2(W10427), .ZN(W11423));
  NOR2X1 G3761 (.A1(W10326), .A2(W10328), .ZN(O508));
  NOR2X1 G3762 (.A1(W378), .A2(W8645), .ZN(W11421));
  NOR2X1 G3763 (.A1(W12357), .A2(W23407), .ZN(W29222));
  NOR2X1 G3764 (.A1(W15274), .A2(W32568), .ZN(O10207));
  NOR2X1 G3765 (.A1(W18391), .A2(W2194), .ZN(W29221));
  NOR2X1 G3766 (.A1(W26048), .A2(W18014), .ZN(O10209));
  NOR2X1 G3767 (.A1(W32839), .A2(W18375), .ZN(O10210));
  NOR2X1 G3768 (.A1(W36738), .A2(W26503), .ZN(O10291));
  NOR2X1 G3769 (.A1(W10973), .A2(W1992), .ZN(W11414));
  NOR2X1 G3770 (.A1(W5118), .A2(W8085), .ZN(O10212));
  NOR2X1 G3771 (.A1(W5874), .A2(W5117), .ZN(W11412));
  NOR2X1 G3772 (.A1(W3240), .A2(W2923), .ZN(W11411));
  NOR2X1 G3773 (.A1(W10757), .A2(W4395), .ZN(W11410));
  NOR2X1 G3774 (.A1(W7459), .A2(W24800), .ZN(O10214));
  NOR2X1 G3775 (.A1(W13263), .A2(W4025), .ZN(O10215));
  NOR2X1 G3776 (.A1(W21639), .A2(W34089), .ZN(W39669));
  NOR2X1 G3777 (.A1(W20917), .A2(W1294), .ZN(W21618));
  NOR2X1 G3778 (.A1(W9985), .A2(W1707), .ZN(W11216));
  NOR2X1 G3779 (.A1(W8211), .A2(W17276), .ZN(O2295));
  NOR2X1 G3780 (.A1(W21824), .A2(W10603), .ZN(O4774));
  NOR2X1 G3781 (.A1(W3968), .A2(W4762), .ZN(O488));
  NOR2X1 G3782 (.A1(W19240), .A2(W2653), .ZN(W21621));
  NOR2X1 G3783 (.A1(W22337), .A2(W10583), .ZN(O10367));
  NOR2X1 G3784 (.A1(W27625), .A2(W16347), .ZN(W39667));
  NOR2X1 G3785 (.A1(W14247), .A2(W39114), .ZN(O10360));
  NOR2X1 G3786 (.A1(W14219), .A2(W18060), .ZN(O2296));
  NOR2X1 G3787 (.A1(W7265), .A2(W26811), .ZN(W39671));
  NOR2X1 G3788 (.A1(W18147), .A2(W33970), .ZN(O10371));
  NOR2X1 G3789 (.A1(W19671), .A2(W8339), .ZN(O2297));
  NOR2X1 G3790 (.A1(W10362), .A2(W17850), .ZN(W39674));
  NOR2X1 G3791 (.A1(W7365), .A2(W4314), .ZN(W11203));
  NOR2X1 G3792 (.A1(W874), .A2(W9578), .ZN(W11201));
  NOR2X1 G3793 (.A1(W3826), .A2(W17225), .ZN(O10375));
  NOR2X1 G3794 (.A1(W1276), .A2(W2420), .ZN(O4775));
  NOR2X1 G3795 (.A1(W5489), .A2(W6366), .ZN(W21616));
  NOR2X1 G3796 (.A1(W5346), .A2(W10486), .ZN(W11233));
  NOR2X1 G3797 (.A1(W23843), .A2(W18360), .ZN(W39641));
  NOR2X1 G3798 (.A1(W1952), .A2(W1275), .ZN(W11231));
  NOR2X1 G3799 (.A1(W975), .A2(W9700), .ZN(W11230));
  NOR2X1 G3800 (.A1(W20821), .A2(W20377), .ZN(O10353));
  NOR2X1 G3801 (.A1(W33568), .A2(W30712), .ZN(W39644));
  NOR2X1 G3802 (.A1(I797), .A2(W7805), .ZN(W11227));
  NOR2X1 G3803 (.A1(W11013), .A2(I338), .ZN(W11199));
  NOR2X1 G3804 (.A1(W26534), .A2(W2134), .ZN(W39646));
  NOR2X1 G3805 (.A1(W6258), .A2(W8940), .ZN(O10357));
  NOR2X1 G3806 (.A1(W3332), .A2(W1037), .ZN(W11223));
  NOR2X1 G3807 (.A1(W3985), .A2(W3136), .ZN(W11222));
  NOR2X1 G3808 (.A1(W5933), .A2(W10795), .ZN(W11221));
  NOR2X1 G3809 (.A1(W6518), .A2(W4173), .ZN(W11220));
  NOR2X1 G3810 (.A1(W11123), .A2(W29059), .ZN(W39652));
  NOR2X1 G3811 (.A1(W10731), .A2(W9410), .ZN(W21631));
  NOR2X1 G3812 (.A1(I1164), .A2(W8615), .ZN(W11180));
  NOR2X1 G3813 (.A1(W10328), .A2(W1099), .ZN(W11179));
  NOR2X1 G3814 (.A1(W9691), .A2(W7371), .ZN(W11178));
  NOR2X1 G3815 (.A1(W9856), .A2(W5473), .ZN(W11177));
  NOR2X1 G3816 (.A1(I1648), .A2(W11329), .ZN(O10384));
  NOR2X1 G3817 (.A1(W8195), .A2(W1400), .ZN(W11175));
  NOR2X1 G3818 (.A1(W3177), .A2(W2091), .ZN(O487));
  NOR2X1 G3819 (.A1(W34949), .A2(W2930), .ZN(O10385));
  NOR2X1 G3820 (.A1(W8593), .A2(W976), .ZN(W11181));
  NOR2X1 G3821 (.A1(I1621), .A2(I1357), .ZN(W11170));
  NOR2X1 G3822 (.A1(W7678), .A2(W10833), .ZN(W11169));
  NOR2X1 G3823 (.A1(W6209), .A2(W9286), .ZN(W11168));
  NOR2X1 G3824 (.A1(I1355), .A2(W2991), .ZN(W11166));
  NOR2X1 G3825 (.A1(W10236), .A2(W32990), .ZN(W39699));
  NOR2X1 G3826 (.A1(W4333), .A2(W20910), .ZN(O10389));
  NOR2X1 G3827 (.A1(W9330), .A2(W9889), .ZN(W11163));
  NOR2X1 G3828 (.A1(I566), .A2(W660), .ZN(W11162));
  NOR2X1 G3829 (.A1(W10860), .A2(W4015), .ZN(W11190));
  NOR2X1 G3830 (.A1(W37575), .A2(W38878), .ZN(O10377));
  NOR2X1 G3831 (.A1(W2527), .A2(W2879), .ZN(W11197));
  NOR2X1 G3832 (.A1(W12520), .A2(W21511), .ZN(W21625));
  NOR2X1 G3833 (.A1(W31995), .A2(W15643), .ZN(W39681));
  NOR2X1 G3834 (.A1(W3446), .A2(W7226), .ZN(W11194));
  NOR2X1 G3835 (.A1(W23472), .A2(W37341), .ZN(O10379));
  NOR2X1 G3836 (.A1(W37758), .A2(W14913), .ZN(W39684));
  NOR2X1 G3837 (.A1(W9854), .A2(I1618), .ZN(W11191));
  NOR2X1 G3838 (.A1(W13257), .A2(W18901), .ZN(W29170));
  NOR2X1 G3839 (.A1(W13823), .A2(W10263), .ZN(W29166));
  NOR2X1 G3840 (.A1(W7523), .A2(I1681), .ZN(W11188));
  NOR2X1 G3841 (.A1(W10337), .A2(W6554), .ZN(O4772));
  NOR2X1 G3842 (.A1(W32428), .A2(W37259), .ZN(W39688));
  NOR2X1 G3843 (.A1(W32033), .A2(W33402), .ZN(O10383));
  NOR2X1 G3844 (.A1(W6334), .A2(W12593), .ZN(W21629));
  NOR2X1 G3845 (.A1(W4651), .A2(W4999), .ZN(W11182));
  NOR2X1 G3846 (.A1(I1500), .A2(W9336), .ZN(W11284));
  NOR2X1 G3847 (.A1(W17633), .A2(W3523), .ZN(W21594));
  NOR2X1 G3848 (.A1(W12438), .A2(W2027), .ZN(W21595));
  NOR2X1 G3849 (.A1(W6687), .A2(W7885), .ZN(W21596));
  NOR2X1 G3850 (.A1(W18780), .A2(I386), .ZN(O10311));
  NOR2X1 G3851 (.A1(W1409), .A2(W39138), .ZN(O10312));
  NOR2X1 G3852 (.A1(W46), .A2(W8429), .ZN(W11287));
  NOR2X1 G3853 (.A1(W5971), .A2(W6561), .ZN(W11286));
  NOR2X1 G3854 (.A1(W3920), .A2(W1843), .ZN(W11285));
  NOR2X1 G3855 (.A1(W27564), .A2(W23136), .ZN(W39575));
  NOR2X1 G3856 (.A1(W3541), .A2(W24141), .ZN(W29186));
  NOR2X1 G3857 (.A1(W32061), .A2(W23051), .ZN(W39589));
  NOR2X1 G3858 (.A1(W38416), .A2(W14536), .ZN(W39590));
  NOR2X1 G3859 (.A1(W1560), .A2(W21651), .ZN(W29185));
  NOR2X1 G3860 (.A1(W17975), .A2(W9680), .ZN(W29184));
  NOR2X1 G3861 (.A1(W10904), .A2(W5822), .ZN(W11278));
  NOR2X1 G3862 (.A1(W8364), .A2(W9327), .ZN(W11277));
  NOR2X1 G3863 (.A1(W6371), .A2(W2220), .ZN(W11276));
  NOR2X1 G3864 (.A1(W3724), .A2(W23722), .ZN(O4783));
  NOR2X1 G3865 (.A1(W1061), .A2(W7216), .ZN(W11311));
  NOR2X1 G3866 (.A1(W18865), .A2(W10446), .ZN(W29194));
  NOR2X1 G3867 (.A1(W14926), .A2(W6172), .ZN(O4785));
  NOR2X1 G3868 (.A1(W3431), .A2(W3469), .ZN(W39561));
  NOR2X1 G3869 (.A1(W13880), .A2(W17520), .ZN(W21588));
  NOR2X1 G3870 (.A1(W25988), .A2(W8619), .ZN(O10295));
  NOR2X1 G3871 (.A1(W6267), .A2(W6937), .ZN(O497));
  NOR2X1 G3872 (.A1(W35660), .A2(W13178), .ZN(W39564));
  NOR2X1 G3873 (.A1(W28577), .A2(W13006), .ZN(O4780));
  NOR2X1 G3874 (.A1(W36912), .A2(W23106), .ZN(O10297));
  NOR2X1 G3875 (.A1(W18247), .A2(I1737), .ZN(W29189));
  NOR2X1 G3876 (.A1(W31950), .A2(W35853), .ZN(O10301));
  NOR2X1 G3877 (.A1(W5605), .A2(W8622), .ZN(W11298));
  NOR2X1 G3878 (.A1(W11155), .A2(W20512), .ZN(W29188));
  NOR2X1 G3879 (.A1(W37396), .A2(W28166), .ZN(O10302));
  NOR2X1 G3880 (.A1(I1815), .A2(W10368), .ZN(W21593));
  NOR2X1 G3881 (.A1(W420), .A2(W18974), .ZN(W21613));
  NOR2X1 G3882 (.A1(W16526), .A2(W12818), .ZN(O10331));
  NOR2X1 G3883 (.A1(W7637), .A2(W11035), .ZN(O493));
  NOR2X1 G3884 (.A1(W10075), .A2(W33110), .ZN(O10333));
  NOR2X1 G3885 (.A1(W4778), .A2(W5467), .ZN(O2294));
  NOR2X1 G3886 (.A1(W14299), .A2(W11804), .ZN(O10336));
  NOR2X1 G3887 (.A1(I398), .A2(W33104), .ZN(O10338));
  NOR2X1 G3888 (.A1(W38333), .A2(W7366), .ZN(O10339));
  NOR2X1 G3889 (.A1(W31674), .A2(W3208), .ZN(O10340));
  NOR2X1 G3890 (.A1(W3488), .A2(W19345), .ZN(O4778));
  NOR2X1 G3891 (.A1(I38), .A2(W7374), .ZN(W11243));
  NOR2X1 G3892 (.A1(W15579), .A2(W32253), .ZN(O10341));
  NOR2X1 G3893 (.A1(W3038), .A2(W1472), .ZN(O491));
  NOR2X1 G3894 (.A1(W3485), .A2(W5600), .ZN(O10342));
  NOR2X1 G3895 (.A1(W1156), .A2(W37692), .ZN(O10344));
  NOR2X1 G3896 (.A1(W38593), .A2(W18487), .ZN(O10347));
  NOR2X1 G3897 (.A1(W4036), .A2(I806), .ZN(W11236));
  NOR2X1 G3898 (.A1(W684), .A2(W3176), .ZN(W21602));
  NOR2X1 G3899 (.A1(W38542), .A2(W34187), .ZN(O10318));
  NOR2X1 G3900 (.A1(W15959), .A2(W39009), .ZN(O10321));
  NOR2X1 G3901 (.A1(W1762), .A2(W2876), .ZN(W11272));
  NOR2X1 G3902 (.A1(W11662), .A2(W3909), .ZN(W39599));
  NOR2X1 G3903 (.A1(W10121), .A2(I232), .ZN(W11270));
  NOR2X1 G3904 (.A1(W8233), .A2(W8415), .ZN(W11269));
  NOR2X1 G3905 (.A1(W29070), .A2(W8803), .ZN(W39600));
  NOR2X1 G3906 (.A1(W6137), .A2(I1859), .ZN(W11267));
  NOR2X1 G3907 (.A1(W23345), .A2(W30110), .ZN(W40016));
  NOR2X1 G3908 (.A1(I549), .A2(W1380), .ZN(O10323));
  NOR2X1 G3909 (.A1(W34447), .A2(W34082), .ZN(O10324));
  NOR2X1 G3910 (.A1(W33409), .A2(W33843), .ZN(O10325));
  NOR2X1 G3911 (.A1(W18875), .A2(W20179), .ZN(O2291));
  NOR2X1 G3912 (.A1(W18616), .A2(W15112), .ZN(W29180));
  NOR2X1 G3913 (.A1(W8900), .A2(W717), .ZN(W11259));
  NOR2X1 G3914 (.A1(I612), .A2(W16123), .ZN(O2292));
  NOR2X1 G3915 (.A1(W23610), .A2(W26552), .ZN(O10919));
  NOR2X1 G3916 (.A1(W3712), .A2(W7277), .ZN(O10905));
  NOR2X1 G3917 (.A1(W26353), .A2(W9393), .ZN(O10907));
  NOR2X1 G3918 (.A1(W7472), .A2(W28646), .ZN(W40451));
  NOR2X1 G3919 (.A1(W26170), .A2(W16886), .ZN(O10914));
  NOR2X1 G3920 (.A1(W19226), .A2(W25476), .ZN(O10915));
  NOR2X1 G3921 (.A1(W18424), .A2(W2782), .ZN(W40460));
  NOR2X1 G3922 (.A1(W2774), .A2(W16954), .ZN(O2354));
  NOR2X1 G3923 (.A1(W5840), .A2(W5146), .ZN(O10917));
  NOR2X1 G3924 (.A1(W8512), .A2(W4174), .ZN(W10437));
  NOR2X1 G3925 (.A1(W18154), .A2(W8123), .ZN(O10921));
  NOR2X1 G3926 (.A1(W9524), .A2(W5810), .ZN(W10424));
  NOR2X1 G3927 (.A1(W33184), .A2(W38735), .ZN(O10922));
  NOR2X1 G3928 (.A1(I402), .A2(I1763), .ZN(W10422));
  NOR2X1 G3929 (.A1(W15872), .A2(W10237), .ZN(W21863));
  NOR2X1 G3930 (.A1(W24302), .A2(W21176), .ZN(W28922));
  NOR2X1 G3931 (.A1(W710), .A2(W5600), .ZN(W10419));
  NOR2X1 G3932 (.A1(W20008), .A2(W20291), .ZN(W21865));
  NOR2X1 G3933 (.A1(W3055), .A2(W8686), .ZN(W10445));
  NOR2X1 G3934 (.A1(I317), .A2(W2892), .ZN(W10453));
  NOR2X1 G3935 (.A1(W9092), .A2(W343), .ZN(W10452));
  NOR2X1 G3936 (.A1(W9845), .A2(W5637), .ZN(W10451));
  NOR2X1 G3937 (.A1(W22315), .A2(W11799), .ZN(O10892));
  NOR2X1 G3938 (.A1(W4991), .A2(W33385), .ZN(O10893));
  NOR2X1 G3939 (.A1(I80), .A2(W29077), .ZN(O10894));
  NOR2X1 G3940 (.A1(W7148), .A2(W4866), .ZN(W10447));
  NOR2X1 G3941 (.A1(W35802), .A2(W27861), .ZN(O10896));
  NOR2X1 G3942 (.A1(I115), .A2(I389), .ZN(W10417));
  NOR2X1 G3943 (.A1(W9923), .A2(W2617), .ZN(W10444));
  NOR2X1 G3944 (.A1(W12525), .A2(I457), .ZN(O10897));
  NOR2X1 G3945 (.A1(W5866), .A2(W1327), .ZN(W10442));
  NOR2X1 G3946 (.A1(W7236), .A2(W3380), .ZN(O10901));
  NOR2X1 G3947 (.A1(W6556), .A2(W6619), .ZN(O390));
  NOR2X1 G3948 (.A1(W17750), .A2(W20241), .ZN(O10902));
  NOR2X1 G3949 (.A1(W23831), .A2(I454), .ZN(O4669));
  NOR2X1 G3950 (.A1(W4875), .A2(W29647), .ZN(O10955));
  NOR2X1 G3951 (.A1(W36302), .A2(I1402), .ZN(O10938));
  NOR2X1 G3952 (.A1(W13161), .A2(W11340), .ZN(W28913));
  NOR2X1 G3953 (.A1(W10342), .A2(W20643), .ZN(O10941));
  NOR2X1 G3954 (.A1(W30047), .A2(W28159), .ZN(W40500));
  NOR2X1 G3955 (.A1(W6918), .A2(W4096), .ZN(O2361));
  NOR2X1 G3956 (.A1(W36335), .A2(W10562), .ZN(O10949));
  NOR2X1 G3957 (.A1(W4978), .A2(W23577), .ZN(W28908));
  NOR2X1 G3958 (.A1(W17220), .A2(W14087), .ZN(O10954));
  NOR2X1 G3959 (.A1(I924), .A2(W2062), .ZN(O10935));
  NOR2X1 G3960 (.A1(W6860), .A2(W18673), .ZN(O2363));
  NOR2X1 G3961 (.A1(I1247), .A2(W19478), .ZN(W28906));
  NOR2X1 G3962 (.A1(W603), .A2(W10843), .ZN(W28902));
  NOR2X1 G3963 (.A1(W5454), .A2(W8216), .ZN(O2364));
  NOR2X1 G3964 (.A1(W37704), .A2(W4303), .ZN(O10958));
  NOR2X1 G3965 (.A1(W15048), .A2(W1556), .ZN(O4660));
  NOR2X1 G3966 (.A1(W10962), .A2(W12223), .ZN(O4659));
  NOR2X1 G3967 (.A1(W11280), .A2(W10600), .ZN(O4656));
  NOR2X1 G3968 (.A1(W33952), .A2(W4465), .ZN(O10930));
  NOR2X1 G3969 (.A1(W7769), .A2(W1707), .ZN(W10415));
  NOR2X1 G3970 (.A1(W15367), .A2(W9570), .ZN(O10927));
  NOR2X1 G3971 (.A1(W19940), .A2(W3966), .ZN(W28918));
  NOR2X1 G3972 (.A1(W15263), .A2(W33371), .ZN(W40477));
  NOR2X1 G3973 (.A1(W14260), .A2(W27450), .ZN(O4666));
  NOR2X1 G3974 (.A1(I1394), .A2(W6299), .ZN(W10410));
  NOR2X1 G3975 (.A1(W28520), .A2(W27281), .ZN(O4665));
  NOR2X1 G3976 (.A1(W32451), .A2(W22961), .ZN(O10929));
  NOR2X1 G3977 (.A1(W5779), .A2(W2484), .ZN(W10454));
  NOR2X1 G3978 (.A1(W8004), .A2(W5153), .ZN(W28914));
  NOR2X1 G3979 (.A1(W35808), .A2(W30041), .ZN(O10933));
  NOR2X1 G3980 (.A1(I1415), .A2(W7146), .ZN(W10403));
  NOR2X1 G3981 (.A1(W871), .A2(W9772), .ZN(W10402));
  NOR2X1 G3982 (.A1(W692), .A2(W9590), .ZN(W10401));
  NOR2X1 G3983 (.A1(W5494), .A2(W6829), .ZN(W10400));
  NOR2X1 G3984 (.A1(W16776), .A2(W2718), .ZN(W40486));
  NOR2X1 G3985 (.A1(W1317), .A2(W1083), .ZN(W10505));
  NOR2X1 G3986 (.A1(W2129), .A2(W4801), .ZN(W10515));
  NOR2X1 G3987 (.A1(W37258), .A2(W5347), .ZN(W40368));
  NOR2X1 G3988 (.A1(W14832), .A2(W14557), .ZN(W21841));
  NOR2X1 G3989 (.A1(W32633), .A2(W39669), .ZN(W40372));
  NOR2X1 G3990 (.A1(W23567), .A2(W2618), .ZN(O4676));
  NOR2X1 G3991 (.A1(W4614), .A2(W3017), .ZN(W10508));
  NOR2X1 G3992 (.A1(W2843), .A2(I181), .ZN(O4675));
  NOR2X1 G3993 (.A1(I1739), .A2(W32815), .ZN(W40378));
  NOR2X1 G3994 (.A1(W5221), .A2(W13571), .ZN(W21839));
  NOR2X1 G3995 (.A1(W11850), .A2(W29372), .ZN(O10849));
  NOR2X1 G3996 (.A1(W2561), .A2(W5006), .ZN(W10503));
  NOR2X1 G3997 (.A1(W6697), .A2(W2433), .ZN(O400));
  NOR2X1 G3998 (.A1(W33333), .A2(W11963), .ZN(O10850));
  NOR2X1 G3999 (.A1(W1317), .A2(W5445), .ZN(W21846));
  NOR2X1 G4000 (.A1(W5968), .A2(W5265), .ZN(O399));
  NOR2X1 G4001 (.A1(W307), .A2(W14630), .ZN(W21848));
  NOR2X1 G4002 (.A1(W15630), .A2(W343), .ZN(O10858));
  NOR2X1 G4003 (.A1(W38282), .A2(W30822), .ZN(O10833));
  NOR2X1 G4004 (.A1(W16484), .A2(W9870), .ZN(O10821));
  NOR2X1 G4005 (.A1(W5476), .A2(W12711), .ZN(W21829));
  NOR2X1 G4006 (.A1(W1272), .A2(W16115), .ZN(O10824));
  NOR2X1 G4007 (.A1(W1997), .A2(W10643), .ZN(W21831));
  NOR2X1 G4008 (.A1(W22107), .A2(W28002), .ZN(W28962));
  NOR2X1 G4009 (.A1(W3953), .A2(W706), .ZN(W10531));
  NOR2X1 G4010 (.A1(W33678), .A2(W34728), .ZN(W40348));
  NOR2X1 G4011 (.A1(W3988), .A2(W21459), .ZN(O10832));
  NOR2X1 G4012 (.A1(I1675), .A2(I1952), .ZN(O398));
  NOR2X1 G4013 (.A1(W4207), .A2(W8195), .ZN(W10526));
  NOR2X1 G4014 (.A1(W21567), .A2(W18752), .ZN(O10834));
  NOR2X1 G4015 (.A1(W9679), .A2(W3562), .ZN(W10524));
  NOR2X1 G4016 (.A1(W9595), .A2(W8942), .ZN(O10836));
  NOR2X1 G4017 (.A1(W25203), .A2(W30461), .ZN(O10837));
  NOR2X1 G4018 (.A1(W29), .A2(W31120), .ZN(O10838));
  NOR2X1 G4019 (.A1(W22973), .A2(W21631), .ZN(O4680));
  NOR2X1 G4020 (.A1(W5199), .A2(W2828), .ZN(W21857));
  NOR2X1 G4021 (.A1(W5299), .A2(W851), .ZN(O10879));
  NOR2X1 G4022 (.A1(W14173), .A2(W38157), .ZN(O10880));
  NOR2X1 G4023 (.A1(W1200), .A2(W3706), .ZN(W10470));
  NOR2X1 G4024 (.A1(W3070), .A2(W9679), .ZN(W10469));
  NOR2X1 G4025 (.A1(I1831), .A2(W446), .ZN(W10468));
  NOR2X1 G4026 (.A1(W10296), .A2(W8387), .ZN(O396));
  NOR2X1 G4027 (.A1(W12413), .A2(W16901), .ZN(W40421));
  NOR2X1 G4028 (.A1(W14960), .A2(W1284), .ZN(O10884));
  NOR2X1 G4029 (.A1(W11887), .A2(W26757), .ZN(W28936));
  NOR2X1 G4030 (.A1(W22688), .A2(W1700), .ZN(O10887));
  NOR2X1 G4031 (.A1(W15184), .A2(W15646), .ZN(O2353));
  NOR2X1 G4032 (.A1(W8996), .A2(W4324), .ZN(O392));
  NOR2X1 G4033 (.A1(W5848), .A2(W1212), .ZN(W10459));
  NOR2X1 G4034 (.A1(W3712), .A2(W8009), .ZN(W10458));
  NOR2X1 G4035 (.A1(W4151), .A2(W3056), .ZN(W10457));
  NOR2X1 G4036 (.A1(W26263), .A2(W5168), .ZN(O10889));
  NOR2X1 G4037 (.A1(W18926), .A2(W11449), .ZN(O10891));
  NOR2X1 G4038 (.A1(I811), .A2(W18669), .ZN(O10868));
  NOR2X1 G4039 (.A1(W18889), .A2(W17583), .ZN(O2352));
  NOR2X1 G4040 (.A1(W11772), .A2(W35247), .ZN(O10861));
  NOR2X1 G4041 (.A1(W8577), .A2(W1652), .ZN(W10491));
  NOR2X1 G4042 (.A1(W9593), .A2(W9108), .ZN(W10490));
  NOR2X1 G4043 (.A1(W20470), .A2(W1646), .ZN(W40396));
  NOR2X1 G4044 (.A1(W37763), .A2(W21932), .ZN(O10864));
  NOR2X1 G4045 (.A1(W1995), .A2(W1554), .ZN(O10865));
  NOR2X1 G4046 (.A1(W11893), .A2(W38060), .ZN(W40400));
  NOR2X1 G4047 (.A1(I217), .A2(I671), .ZN(W10375));
  NOR2X1 G4048 (.A1(W6503), .A2(W8998), .ZN(W10482));
  NOR2X1 G4049 (.A1(W6565), .A2(W6465), .ZN(W21852));
  NOR2X1 G4050 (.A1(W9263), .A2(I1119), .ZN(W10480));
  NOR2X1 G4051 (.A1(W10221), .A2(W21124), .ZN(W40408));
  NOR2X1 G4052 (.A1(I61), .A2(I1944), .ZN(O10873));
  NOR2X1 G4053 (.A1(I1690), .A2(W35571), .ZN(O10874));
  NOR2X1 G4054 (.A1(W34620), .A2(W26276), .ZN(O10875));
  NOR2X1 G4055 (.A1(W3293), .A2(W7472), .ZN(W10269));
  NOR2X1 G4056 (.A1(W3205), .A2(W28541), .ZN(O11013));
  NOR2X1 G4057 (.A1(W25312), .A2(W16529), .ZN(W40601));
  NOR2X1 G4058 (.A1(W1196), .A2(W979), .ZN(O11016));
  NOR2X1 G4059 (.A1(W2309), .A2(W6275), .ZN(W10275));
  NOR2X1 G4060 (.A1(W12173), .A2(W24418), .ZN(O11020));
  NOR2X1 G4061 (.A1(W19700), .A2(W9747), .ZN(O2373));
  NOR2X1 G4062 (.A1(W3966), .A2(W6451), .ZN(O11023));
  NOR2X1 G4063 (.A1(W3117), .A2(W6112), .ZN(W10270));
  NOR2X1 G4064 (.A1(I284), .A2(W25807), .ZN(O4650));
  NOR2X1 G4065 (.A1(W19965), .A2(W28853), .ZN(O11024));
  NOR2X1 G4066 (.A1(W19825), .A2(W1179), .ZN(O11025));
  NOR2X1 G4067 (.A1(W26573), .A2(W17133), .ZN(W40614));
  NOR2X1 G4068 (.A1(W5695), .A2(W9012), .ZN(W10265));
  NOR2X1 G4069 (.A1(W4110), .A2(W21051), .ZN(W21909));
  NOR2X1 G4070 (.A1(W9303), .A2(W8856), .ZN(W10263));
  NOR2X1 G4071 (.A1(W2504), .A2(W10975), .ZN(O11027));
  NOR2X1 G4072 (.A1(W19667), .A2(W16781), .ZN(W28871));
  NOR2X1 G4073 (.A1(W36060), .A2(W29107), .ZN(O11009));
  NOR2X1 G4074 (.A1(W25880), .A2(W32992), .ZN(O11001));
  NOR2X1 G4075 (.A1(W37612), .A2(W3646), .ZN(W40587));
  NOR2X1 G4076 (.A1(W8247), .A2(W23077), .ZN(O11004));
  NOR2X1 G4077 (.A1(W4902), .A2(I1894), .ZN(W10294));
  NOR2X1 G4078 (.A1(W3240), .A2(I1043), .ZN(W10293));
  NOR2X1 G4079 (.A1(W30331), .A2(W995), .ZN(O11005));
  NOR2X1 G4080 (.A1(W30291), .A2(W22327), .ZN(O11006));
  NOR2X1 G4081 (.A1(W21596), .A2(I1123), .ZN(O11008));
  NOR2X1 G4082 (.A1(W9495), .A2(W18438), .ZN(W28868));
  NOR2X1 G4083 (.A1(W4102), .A2(I195), .ZN(O377));
  NOR2X1 G4084 (.A1(W4020), .A2(W267), .ZN(W10287));
  NOR2X1 G4085 (.A1(W7563), .A2(W2031), .ZN(W10286));
  NOR2X1 G4086 (.A1(W4871), .A2(W8965), .ZN(W10285));
  NOR2X1 G4087 (.A1(W31049), .A2(I828), .ZN(O11010));
  NOR2X1 G4088 (.A1(W8687), .A2(W1009), .ZN(W10283));
  NOR2X1 G4089 (.A1(W33379), .A2(W16114), .ZN(O11011));
  NOR2X1 G4090 (.A1(W5556), .A2(W8072), .ZN(W10225));
  NOR2X1 G4091 (.A1(W5678), .A2(W7144), .ZN(W10237));
  NOR2X1 G4092 (.A1(I1510), .A2(W32750), .ZN(O11045));
  NOR2X1 G4093 (.A1(W13011), .A2(W8885), .ZN(W40640));
  NOR2X1 G4094 (.A1(W4690), .A2(W1076), .ZN(O11046));
  NOR2X1 G4095 (.A1(W6517), .A2(W6115), .ZN(W10232));
  NOR2X1 G4096 (.A1(W7061), .A2(W26548), .ZN(O11048));
  NOR2X1 G4097 (.A1(W35707), .A2(I1036), .ZN(O11052));
  NOR2X1 G4098 (.A1(W13793), .A2(W9026), .ZN(O11053));
  NOR2X1 G4099 (.A1(W28515), .A2(W1984), .ZN(O11043));
  NOR2X1 G4100 (.A1(W8329), .A2(W6387), .ZN(W10224));
  NOR2X1 G4101 (.A1(I147), .A2(W9759), .ZN(W10223));
  NOR2X1 G4102 (.A1(I499), .A2(W945), .ZN(W10222));
  NOR2X1 G4103 (.A1(W16725), .A2(W13751), .ZN(O11054));
  NOR2X1 G4104 (.A1(W1127), .A2(W1115), .ZN(W40654));
  NOR2X1 G4105 (.A1(W31146), .A2(W529), .ZN(W40655));
  NOR2X1 G4106 (.A1(W9987), .A2(W2555), .ZN(W21921));
  NOR2X1 G4107 (.A1(W10003), .A2(W3729), .ZN(W10217));
  NOR2X1 G4108 (.A1(W33925), .A2(W11276), .ZN(O11034));
  NOR2X1 G4109 (.A1(W505), .A2(W8713), .ZN(W10259));
  NOR2X1 G4110 (.A1(I1710), .A2(W2685), .ZN(W10258));
  NOR2X1 G4111 (.A1(W8768), .A2(W9622), .ZN(W10257));
  NOR2X1 G4112 (.A1(W5687), .A2(W3609), .ZN(W10256));
  NOR2X1 G4113 (.A1(W1663), .A2(W132), .ZN(W10254));
  NOR2X1 G4114 (.A1(W7946), .A2(W7112), .ZN(W10253));
  NOR2X1 G4115 (.A1(W10441), .A2(W12963), .ZN(O11033));
  NOR2X1 G4116 (.A1(W8941), .A2(W1775), .ZN(O373));
  NOR2X1 G4117 (.A1(W20554), .A2(W10140), .ZN(O11000));
  NOR2X1 G4118 (.A1(W7992), .A2(W30538), .ZN(O11035));
  NOR2X1 G4119 (.A1(W29658), .A2(W34355), .ZN(O11038));
  NOR2X1 G4120 (.A1(W3676), .A2(W5365), .ZN(W10244));
  NOR2X1 G4121 (.A1(W561), .A2(W119), .ZN(W10243));
  NOR2X1 G4122 (.A1(W8680), .A2(W9616), .ZN(W10241));
  NOR2X1 G4123 (.A1(W25570), .A2(W694), .ZN(O11040));
  NOR2X1 G4124 (.A1(W22315), .A2(W19984), .ZN(O11041));
  NOR2X1 G4125 (.A1(W10776), .A2(W4317), .ZN(O4652));
  NOR2X1 G4126 (.A1(I936), .A2(I412), .ZN(W10355));
  NOR2X1 G4127 (.A1(W10222), .A2(W7837), .ZN(W10354));
  NOR2X1 G4128 (.A1(W1693), .A2(W2657), .ZN(W10353));
  NOR2X1 G4129 (.A1(W7476), .A2(W17706), .ZN(W40537));
  NOR2X1 G4130 (.A1(W26473), .A2(W14657), .ZN(O10970));
  NOR2X1 G4131 (.A1(W18078), .A2(W636), .ZN(W21892));
  NOR2X1 G4132 (.A1(W31844), .A2(W27157), .ZN(O10972));
  NOR2X1 G4133 (.A1(W32753), .A2(W5003), .ZN(W40542));
  NOR2X1 G4134 (.A1(W33477), .A2(W18963), .ZN(O10969));
  NOR2X1 G4135 (.A1(I1888), .A2(W5611), .ZN(W10346));
  NOR2X1 G4136 (.A1(W4004), .A2(I1096), .ZN(W10344));
  NOR2X1 G4137 (.A1(W3553), .A2(I1104), .ZN(W10343));
  NOR2X1 G4138 (.A1(W27990), .A2(I1104), .ZN(O10976));
  NOR2X1 G4139 (.A1(W40354), .A2(W36843), .ZN(O10977));
  NOR2X1 G4140 (.A1(I1325), .A2(W18019), .ZN(O10978));
  NOR2X1 G4141 (.A1(W7360), .A2(W5744), .ZN(W10339));
  NOR2X1 G4142 (.A1(W2803), .A2(I74), .ZN(W10338));
  NOR2X1 G4143 (.A1(W9054), .A2(W2367), .ZN(O10965));
  NOR2X1 G4144 (.A1(W7408), .A2(W795), .ZN(W10374));
  NOR2X1 G4145 (.A1(W39417), .A2(I564), .ZN(O10962));
  NOR2X1 G4146 (.A1(W1493), .A2(W9896), .ZN(W10372));
  NOR2X1 G4147 (.A1(W5831), .A2(W6528), .ZN(W10370));
  NOR2X1 G4148 (.A1(W3265), .A2(W7385), .ZN(W10369));
  NOR2X1 G4149 (.A1(I1308), .A2(W18087), .ZN(W21888));
  NOR2X1 G4150 (.A1(W10093), .A2(W1782), .ZN(W10367));
  NOR2X1 G4151 (.A1(W3695), .A2(W8688), .ZN(W10366));
  NOR2X1 G4152 (.A1(W1301), .A2(W4335), .ZN(W10337));
  NOR2X1 G4153 (.A1(W2335), .A2(W3588), .ZN(W10364));
  NOR2X1 G4154 (.A1(W18555), .A2(W15619), .ZN(W21889));
  NOR2X1 G4155 (.A1(W8094), .A2(W4576), .ZN(W10362));
  NOR2X1 G4156 (.A1(W2458), .A2(W1014), .ZN(O4653));
  NOR2X1 G4157 (.A1(W7487), .A2(W7915), .ZN(W10360));
  NOR2X1 G4158 (.A1(W22986), .A2(W1486), .ZN(O10967));
  NOR2X1 G4159 (.A1(W8783), .A2(W3363), .ZN(O383));
  NOR2X1 G4160 (.A1(W36041), .A2(W28851), .ZN(O10994));
  NOR2X1 G4161 (.A1(W8756), .A2(W3918), .ZN(W10315));
  NOR2X1 G4162 (.A1(W14641), .A2(W4909), .ZN(O10990));
  NOR2X1 G4163 (.A1(W28412), .A2(W36618), .ZN(W40568));
  NOR2X1 G4164 (.A1(W35167), .A2(W29660), .ZN(W40569));
  NOR2X1 G4165 (.A1(W23453), .A2(I1059), .ZN(O10991));
  NOR2X1 G4166 (.A1(W8956), .A2(W14886), .ZN(W21901));
  NOR2X1 G4167 (.A1(W25938), .A2(W7783), .ZN(O10993));
  NOR2X1 G4168 (.A1(W9572), .A2(W5776), .ZN(W10308));
  NOR2X1 G4169 (.A1(W4973), .A2(I797), .ZN(W10316));
  NOR2X1 G4170 (.A1(W24203), .A2(W23108), .ZN(W40575));
  NOR2X1 G4171 (.A1(W904), .A2(W5414), .ZN(W10305));
  NOR2X1 G4172 (.A1(W18193), .A2(W16831), .ZN(O2371));
  NOR2X1 G4173 (.A1(W27738), .A2(W3647), .ZN(O4651));
  NOR2X1 G4174 (.A1(W33810), .A2(W13249), .ZN(O10996));
  NOR2X1 G4175 (.A1(W20402), .A2(W29198), .ZN(O10998));
  NOR2X1 G4176 (.A1(W36890), .A2(W8142), .ZN(W40582));
  NOR2X1 G4177 (.A1(W126), .A2(W4823), .ZN(W10299));
  NOR2X1 G4178 (.A1(W2053), .A2(W18233), .ZN(W40558));
  NOR2X1 G4179 (.A1(W5520), .A2(W918), .ZN(W10336));
  NOR2X1 G4180 (.A1(W3827), .A2(W1484), .ZN(W10335));
  NOR2X1 G4181 (.A1(W1342), .A2(W5136), .ZN(W10334));
  NOR2X1 G4182 (.A1(W5704), .A2(W7628), .ZN(W10333));
  NOR2X1 G4183 (.A1(W5271), .A2(W8065), .ZN(W10331));
  NOR2X1 G4184 (.A1(W3084), .A2(W9290), .ZN(W10330));
  NOR2X1 G4185 (.A1(W9341), .A2(W6678), .ZN(W10328));
  NOR2X1 G4186 (.A1(W32022), .A2(W2293), .ZN(O10983));
  NOR2X1 G4187 (.A1(W20900), .A2(W27856), .ZN(W40339));
  NOR2X1 G4188 (.A1(I1888), .A2(W3620), .ZN(W10324));
  NOR2X1 G4189 (.A1(W334), .A2(W6031), .ZN(W10323));
  NOR2X1 G4190 (.A1(I364), .A2(W1615), .ZN(W10321));
  NOR2X1 G4191 (.A1(W1706), .A2(W25605), .ZN(W28882));
  NOR2X1 G4192 (.A1(W2189), .A2(I1429), .ZN(W10319));
  NOR2X1 G4193 (.A1(W9511), .A2(W18966), .ZN(W21900));
  NOR2X1 G4194 (.A1(W3928), .A2(W3861), .ZN(W10317));
  NOR2X1 G4195 (.A1(W5822), .A2(W3267), .ZN(W10746));
  NOR2X1 G4196 (.A1(I693), .A2(W10650), .ZN(W10754));
  NOR2X1 G4197 (.A1(W30053), .A2(W3258), .ZN(W40108));
  NOR2X1 G4198 (.A1(W20135), .A2(W38789), .ZN(O10678));
  NOR2X1 G4199 (.A1(W10184), .A2(W58), .ZN(O430));
  NOR2X1 G4200 (.A1(W643), .A2(W17614), .ZN(O10679));
  NOR2X1 G4201 (.A1(W34187), .A2(W37812), .ZN(O10680));
  NOR2X1 G4202 (.A1(I1261), .A2(W7533), .ZN(O10682));
  NOR2X1 G4203 (.A1(W8592), .A2(W8089), .ZN(O2328));
  NOR2X1 G4204 (.A1(I1486), .A2(W134), .ZN(W10755));
  NOR2X1 G4205 (.A1(W27746), .A2(W26992), .ZN(W40124));
  NOR2X1 G4206 (.A1(W21278), .A2(W9674), .ZN(O4716));
  NOR2X1 G4207 (.A1(W3480), .A2(W4637), .ZN(O429));
  NOR2X1 G4208 (.A1(W721), .A2(W9386), .ZN(W10739));
  NOR2X1 G4209 (.A1(W9328), .A2(W3026), .ZN(W10738));
  NOR2X1 G4210 (.A1(W36872), .A2(W39012), .ZN(W40133));
  NOR2X1 G4211 (.A1(W8544), .A2(W303), .ZN(W10735));
  NOR2X1 G4212 (.A1(W35512), .A2(W12132), .ZN(W40134));
  NOR2X1 G4213 (.A1(W33325), .A2(W24201), .ZN(O10672));
  NOR2X1 G4214 (.A1(W4825), .A2(W1251), .ZN(O433));
  NOR2X1 G4215 (.A1(W7552), .A2(W32458), .ZN(O10663));
  NOR2X1 G4216 (.A1(W9279), .A2(W2628), .ZN(W10769));
  NOR2X1 G4217 (.A1(W9426), .A2(I1088), .ZN(W10768));
  NOR2X1 G4218 (.A1(W16766), .A2(I1659), .ZN(W21759));
  NOR2X1 G4219 (.A1(I1104), .A2(W17396), .ZN(W40100));
  NOR2X1 G4220 (.A1(W23520), .A2(W26476), .ZN(O10670));
  NOR2X1 G4221 (.A1(W19651), .A2(W32577), .ZN(O10671));
  NOR2X1 G4222 (.A1(W1718), .A2(W1434), .ZN(O428));
  NOR2X1 G4223 (.A1(W2584), .A2(I1281), .ZN(W10762));
  NOR2X1 G4224 (.A1(W10254), .A2(W625), .ZN(W10761));
  NOR2X1 G4225 (.A1(W2416), .A2(I1546), .ZN(W10760));
  NOR2X1 G4226 (.A1(W35839), .A2(W12140), .ZN(O10673));
  NOR2X1 G4227 (.A1(W10561), .A2(W8570), .ZN(O431));
  NOR2X1 G4228 (.A1(W8822), .A2(W17837), .ZN(W29041));
  NOR2X1 G4229 (.A1(W17209), .A2(W29126), .ZN(W40107));
  NOR2X1 G4230 (.A1(W22459), .A2(W20423), .ZN(W29024));
  NOR2X1 G4231 (.A1(W1134), .A2(W19853), .ZN(W40154));
  NOR2X1 G4232 (.A1(W5892), .A2(W6508), .ZN(W10713));
  NOR2X1 G4233 (.A1(W14609), .A2(W21164), .ZN(O10710));
  NOR2X1 G4234 (.A1(W10704), .A2(W7443), .ZN(W10711));
  NOR2X1 G4235 (.A1(W17077), .A2(W13055), .ZN(O4710));
  NOR2X1 G4236 (.A1(W2869), .A2(W2191), .ZN(W10709));
  NOR2X1 G4237 (.A1(W6518), .A2(W9158), .ZN(W10708));
  NOR2X1 G4238 (.A1(W28614), .A2(W22986), .ZN(O4709));
  NOR2X1 G4239 (.A1(W23980), .A2(W5825), .ZN(O10709));
  NOR2X1 G4240 (.A1(W7742), .A2(W2302), .ZN(W10705));
  NOR2X1 G4241 (.A1(W24644), .A2(W23956), .ZN(W29023));
  NOR2X1 G4242 (.A1(W2376), .A2(W19905), .ZN(O10714));
  NOR2X1 G4243 (.A1(W10377), .A2(I1076), .ZN(W10702));
  NOR2X1 G4244 (.A1(W454), .A2(W36353), .ZN(O10716));
  NOR2X1 G4245 (.A1(W5860), .A2(W2900), .ZN(W10700));
  NOR2X1 G4246 (.A1(W29126), .A2(W15410), .ZN(W40171));
  NOR2X1 G4247 (.A1(W9796), .A2(W1737), .ZN(W10697));
  NOR2X1 G4248 (.A1(W2907), .A2(I1824), .ZN(O426));
  NOR2X1 G4249 (.A1(W20237), .A2(W30373), .ZN(O10695));
  NOR2X1 G4250 (.A1(W8096), .A2(W7317), .ZN(W10731));
  NOR2X1 G4251 (.A1(W23750), .A2(W39298), .ZN(O10697));
  NOR2X1 G4252 (.A1(W11473), .A2(W6210), .ZN(O10699));
  NOR2X1 G4253 (.A1(W27277), .A2(W17429), .ZN(W40142));
  NOR2X1 G4254 (.A1(W21838), .A2(W36348), .ZN(O10701));
  NOR2X1 G4255 (.A1(W5403), .A2(I923), .ZN(W10726));
  NOR2X1 G4256 (.A1(W4255), .A2(I944), .ZN(O10704));
  NOR2X1 G4257 (.A1(I1270), .A2(W28632), .ZN(W29047));
  NOR2X1 G4258 (.A1(W26486), .A2(W8943), .ZN(O10705));
  NOR2X1 G4259 (.A1(W12241), .A2(W15740), .ZN(O10706));
  NOR2X1 G4260 (.A1(W4494), .A2(W21461), .ZN(W29029));
  NOR2X1 G4261 (.A1(W757), .A2(W10127), .ZN(W10719));
  NOR2X1 G4262 (.A1(W39336), .A2(W21889), .ZN(O10708));
  NOR2X1 G4263 (.A1(W53), .A2(W4569), .ZN(W10717));
  NOR2X1 G4264 (.A1(W145), .A2(I774), .ZN(W10716));
  NOR2X1 G4265 (.A1(W1973), .A2(W7061), .ZN(W10822));
  NOR2X1 G4266 (.A1(W10446), .A2(W3388), .ZN(W10833));
  NOR2X1 G4267 (.A1(W5908), .A2(W2319), .ZN(W10832));
  NOR2X1 G4268 (.A1(W31629), .A2(W20811), .ZN(O10627));
  NOR2X1 G4269 (.A1(W10212), .A2(W19904), .ZN(W40038));
  NOR2X1 G4270 (.A1(I1686), .A2(W20043), .ZN(O10631));
  NOR2X1 G4271 (.A1(W8956), .A2(W9972), .ZN(W29063));
  NOR2X1 G4272 (.A1(W7360), .A2(W12962), .ZN(O10633));
  NOR2X1 G4273 (.A1(W1013), .A2(W10512), .ZN(W10824));
  NOR2X1 G4274 (.A1(W4487), .A2(W10299), .ZN(W10834));
  NOR2X1 G4275 (.A1(W39086), .A2(I1302), .ZN(W40049));
  NOR2X1 G4276 (.A1(W7453), .A2(W595), .ZN(W10820));
  NOR2X1 G4277 (.A1(W4759), .A2(W765), .ZN(W10819));
  NOR2X1 G4278 (.A1(W405), .A2(I269), .ZN(W10817));
  NOR2X1 G4279 (.A1(W3364), .A2(W7001), .ZN(W10816));
  NOR2X1 G4280 (.A1(W21300), .A2(W39527), .ZN(W40052));
  NOR2X1 G4281 (.A1(W16010), .A2(W160), .ZN(W21742));
  NOR2X1 G4282 (.A1(W2746), .A2(W5668), .ZN(O10637));
  NOR2X1 G4283 (.A1(W9165), .A2(W8573), .ZN(W10843));
  NOR2X1 G4284 (.A1(W21128), .A2(W6317), .ZN(W21732));
  NOR2X1 G4285 (.A1(W3763), .A2(W8515), .ZN(O10614));
  NOR2X1 G4286 (.A1(W2758), .A2(W8993), .ZN(W10849));
  NOR2X1 G4287 (.A1(W24560), .A2(I1299), .ZN(O10618));
  NOR2X1 G4288 (.A1(W15714), .A2(W33396), .ZN(W40025));
  NOR2X1 G4289 (.A1(W17944), .A2(I698), .ZN(O2319));
  NOR2X1 G4290 (.A1(W5428), .A2(W11543), .ZN(W29067));
  NOR2X1 G4291 (.A1(W19561), .A2(W33746), .ZN(O10620));
  NOR2X1 G4292 (.A1(W34457), .A2(W12577), .ZN(W40056));
  NOR2X1 G4293 (.A1(W21402), .A2(W22308), .ZN(O10622));
  NOR2X1 G4294 (.A1(I559), .A2(W9344), .ZN(W10840));
  NOR2X1 G4295 (.A1(W13422), .A2(W6631), .ZN(W21736));
  NOR2X1 G4296 (.A1(W5875), .A2(W15450), .ZN(O10623));
  NOR2X1 G4297 (.A1(W32892), .A2(W2923), .ZN(O10624));
  NOR2X1 G4298 (.A1(W104), .A2(I902), .ZN(W10836));
  NOR2X1 G4299 (.A1(W8536), .A2(W8973), .ZN(W10835));
  NOR2X1 G4300 (.A1(I153), .A2(W30253), .ZN(O10655));
  NOR2X1 G4301 (.A1(W8805), .A2(W20797), .ZN(O4723));
  NOR2X1 G4302 (.A1(W4590), .A2(W10608), .ZN(W10791));
  NOR2X1 G4303 (.A1(W6062), .A2(W9041), .ZN(O435));
  NOR2X1 G4304 (.A1(W3989), .A2(W249), .ZN(W21749));
  NOR2X1 G4305 (.A1(I1996), .A2(W20998), .ZN(W21750));
  NOR2X1 G4306 (.A1(W4925), .A2(W5799), .ZN(W10786));
  NOR2X1 G4307 (.A1(W31465), .A2(I1872), .ZN(O10653));
  NOR2X1 G4308 (.A1(I1632), .A2(W4706), .ZN(W10784));
  NOR2X1 G4309 (.A1(W34911), .A2(W34941), .ZN(W40076));
  NOR2X1 G4310 (.A1(W4776), .A2(W7686), .ZN(W10782));
  NOR2X1 G4311 (.A1(W8808), .A2(W7075), .ZN(W10781));
  NOR2X1 G4312 (.A1(W17352), .A2(W10133), .ZN(W21751));
  NOR2X1 G4313 (.A1(W678), .A2(W19817), .ZN(W21753));
  NOR2X1 G4314 (.A1(W29225), .A2(W2407), .ZN(W40089));
  NOR2X1 G4315 (.A1(W8471), .A2(W9953), .ZN(O4721));
  NOR2X1 G4316 (.A1(W138), .A2(W10334), .ZN(O4720));
  NOR2X1 G4317 (.A1(W17607), .A2(W5582), .ZN(W21756));
  NOR2X1 G4318 (.A1(I940), .A2(W1696), .ZN(O437));
  NOR2X1 G4319 (.A1(W8236), .A2(W9580), .ZN(W10811));
  NOR2X1 G4320 (.A1(W36633), .A2(W14124), .ZN(O10638));
  NOR2X1 G4321 (.A1(W4262), .A2(W20126), .ZN(O10640));
  NOR2X1 G4322 (.A1(W19927), .A2(W5052), .ZN(O10641));
  NOR2X1 G4323 (.A1(W11684), .A2(W8219), .ZN(W29058));
  NOR2X1 G4324 (.A1(W35993), .A2(W31088), .ZN(O10645));
  NOR2X1 G4325 (.A1(W15610), .A2(W11869), .ZN(W40066));
  NOR2X1 G4326 (.A1(W5852), .A2(W13811), .ZN(W40067));
  NOR2X1 G4327 (.A1(W5448), .A2(W7780), .ZN(W10696));
  NOR2X1 G4328 (.A1(I551), .A2(W5746), .ZN(O10646));
  NOR2X1 G4329 (.A1(W37455), .A2(W2507), .ZN(W40071));
  NOR2X1 G4330 (.A1(W26592), .A2(W4652), .ZN(O10648));
  NOR2X1 G4331 (.A1(W8128), .A2(W8671), .ZN(W10797));
  NOR2X1 G4332 (.A1(W17953), .A2(I232), .ZN(W21746));
  NOR2X1 G4333 (.A1(W5823), .A2(W34475), .ZN(O10650));
  NOR2X1 G4334 (.A1(W28879), .A2(W16096), .ZN(O10651));
  NOR2X1 G4335 (.A1(W39528), .A2(W14498), .ZN(W40281));
  NOR2X1 G4336 (.A1(I1409), .A2(W5581), .ZN(W10596));
  NOR2X1 G4337 (.A1(W1469), .A2(W23053), .ZN(O10785));
  NOR2X1 G4338 (.A1(W22689), .A2(W2947), .ZN(O10787));
  NOR2X1 G4339 (.A1(W23388), .A2(W10086), .ZN(W40275));
  NOR2X1 G4340 (.A1(W37554), .A2(I1334), .ZN(W40276));
  NOR2X1 G4341 (.A1(W3945), .A2(W60), .ZN(W10591));
  NOR2X1 G4342 (.A1(W6329), .A2(W11111), .ZN(W21808));
  NOR2X1 G4343 (.A1(W4755), .A2(W628), .ZN(W21809));
  NOR2X1 G4344 (.A1(W37726), .A2(W5236), .ZN(O10784));
  NOR2X1 G4345 (.A1(W23185), .A2(W24290), .ZN(W28983));
  NOR2X1 G4346 (.A1(W1515), .A2(W5834), .ZN(W10584));
  NOR2X1 G4347 (.A1(W18459), .A2(W15237), .ZN(O4691));
  NOR2X1 G4348 (.A1(W31952), .A2(W6161), .ZN(O10795));
  NOR2X1 G4349 (.A1(W5671), .A2(W4004), .ZN(O10797));
  NOR2X1 G4350 (.A1(W8239), .A2(W3581), .ZN(W10578));
  NOR2X1 G4351 (.A1(W1078), .A2(W4381), .ZN(W10577));
  NOR2X1 G4352 (.A1(W14623), .A2(W20993), .ZN(O2342));
  NOR2X1 G4353 (.A1(W9985), .A2(W16453), .ZN(W40263));
  NOR2X1 G4354 (.A1(W10401), .A2(W7125), .ZN(O410));
  NOR2X1 G4355 (.A1(W7727), .A2(W5841), .ZN(W10612));
  NOR2X1 G4356 (.A1(W10364), .A2(W6931), .ZN(O4694));
  NOR2X1 G4357 (.A1(W8296), .A2(W4484), .ZN(W10610));
  NOR2X1 G4358 (.A1(W4920), .A2(W8984), .ZN(W21803));
  NOR2X1 G4359 (.A1(W4562), .A2(W26203), .ZN(W28986));
  NOR2X1 G4360 (.A1(W27525), .A2(W4638), .ZN(W28985));
  NOR2X1 G4361 (.A1(I1512), .A2(W17944), .ZN(W21806));
  NOR2X1 G4362 (.A1(W36194), .A2(W4170), .ZN(W40296));
  NOR2X1 G4363 (.A1(W27889), .A2(W10323), .ZN(W40264));
  NOR2X1 G4364 (.A1(W10207), .A2(W23919), .ZN(O10781));
  NOR2X1 G4365 (.A1(W6774), .A2(W13299), .ZN(W21807));
  NOR2X1 G4366 (.A1(W2783), .A2(W23068), .ZN(O10782));
  NOR2X1 G4367 (.A1(W1557), .A2(W5588), .ZN(W10600));
  NOR2X1 G4368 (.A1(W8084), .A2(W7550), .ZN(W10599));
  NOR2X1 G4369 (.A1(W27015), .A2(W1072), .ZN(O10783));
  NOR2X1 G4370 (.A1(W9939), .A2(W3637), .ZN(O10816));
  NOR2X1 G4371 (.A1(W19460), .A2(W15250), .ZN(O4686));
  NOR2X1 G4372 (.A1(I1465), .A2(W8560), .ZN(W10555));
  NOR2X1 G4373 (.A1(W14591), .A2(W12759), .ZN(W40323));
  NOR2X1 G4374 (.A1(W17910), .A2(W11748), .ZN(W21825));
  NOR2X1 G4375 (.A1(W17774), .A2(W3313), .ZN(O4685));
  NOR2X1 G4376 (.A1(W24102), .A2(W32345), .ZN(W40327));
  NOR2X1 G4377 (.A1(W2020), .A2(W4043), .ZN(W10550));
  NOR2X1 G4378 (.A1(W40178), .A2(W34205), .ZN(O10814));
  NOR2X1 G4379 (.A1(W6850), .A2(W35923), .ZN(O10812));
  NOR2X1 G4380 (.A1(W17174), .A2(W19910), .ZN(W28967));
  NOR2X1 G4381 (.A1(W26206), .A2(W17331), .ZN(W40335));
  NOR2X1 G4382 (.A1(W36), .A2(W10397), .ZN(W21828));
  NOR2X1 G4383 (.A1(W6676), .A2(W2957), .ZN(W10544));
  NOR2X1 G4384 (.A1(W8083), .A2(W6873), .ZN(W10543));
  NOR2X1 G4385 (.A1(I1477), .A2(W16890), .ZN(O10820));
  NOR2X1 G4386 (.A1(W29409), .A2(W26024), .ZN(W40338));
  NOR2X1 G4387 (.A1(W9230), .A2(W7505), .ZN(W10540));
  NOR2X1 G4388 (.A1(W10220), .A2(W3624), .ZN(W10565));
  NOR2X1 G4389 (.A1(W8025), .A2(W441), .ZN(O407));
  NOR2X1 G4390 (.A1(W26596), .A2(W29928), .ZN(O10804));
  NOR2X1 G4391 (.A1(W11039), .A2(W13809), .ZN(W21818));
  NOR2X1 G4392 (.A1(W322), .A2(W3423), .ZN(O406));
  NOR2X1 G4393 (.A1(W30432), .A2(W38139), .ZN(W40304));
  NOR2X1 G4394 (.A1(W10829), .A2(W15678), .ZN(O2343));
  NOR2X1 G4395 (.A1(W1998), .A2(W4343), .ZN(W10567));
  NOR2X1 G4396 (.A1(W12513), .A2(I892), .ZN(W28973));
  NOR2X1 G4397 (.A1(W1393), .A2(W7695), .ZN(W10615));
  NOR2X1 G4398 (.A1(W37405), .A2(W23877), .ZN(O10809));
  NOR2X1 G4399 (.A1(W2869), .A2(W26870), .ZN(W28972));
  NOR2X1 G4400 (.A1(W5563), .A2(W9782), .ZN(W10562));
  NOR2X1 G4401 (.A1(W23967), .A2(W22721), .ZN(W40317));
  NOR2X1 G4402 (.A1(W4275), .A2(W5925), .ZN(W10560));
  NOR2X1 G4403 (.A1(W14447), .A2(I1197), .ZN(W28971));
  NOR2X1 G4404 (.A1(W4234), .A2(I1113), .ZN(W21823));
  NOR2X1 G4405 (.A1(W1525), .A2(W8677), .ZN(W10664));
  NOR2X1 G4406 (.A1(W5863), .A2(W2326), .ZN(W10673));
  NOR2X1 G4407 (.A1(W34196), .A2(W9745), .ZN(W40200));
  NOR2X1 G4408 (.A1(W11428), .A2(W13341), .ZN(O10737));
  NOR2X1 G4409 (.A1(W33253), .A2(W29661), .ZN(O10738));
  NOR2X1 G4410 (.A1(W8815), .A2(W4515), .ZN(O419));
  NOR2X1 G4411 (.A1(W34812), .A2(W1619), .ZN(O10741));
  NOR2X1 G4412 (.A1(W1423), .A2(W27886), .ZN(O10743));
  NOR2X1 G4413 (.A1(W35482), .A2(W710), .ZN(O10744));
  NOR2X1 G4414 (.A1(W4065), .A2(W5205), .ZN(W10674));
  NOR2X1 G4415 (.A1(W11055), .A2(W30869), .ZN(O10745));
  NOR2X1 G4416 (.A1(W19823), .A2(W15237), .ZN(W40211));
  NOR2X1 G4417 (.A1(W6779), .A2(W3473), .ZN(W10661));
  NOR2X1 G4418 (.A1(W2776), .A2(W4562), .ZN(O418));
  NOR2X1 G4419 (.A1(I1003), .A2(W10509), .ZN(W10659));
  NOR2X1 G4420 (.A1(W37103), .A2(W34206), .ZN(W40212));
  NOR2X1 G4421 (.A1(W7128), .A2(W9018), .ZN(W10657));
  NOR2X1 G4422 (.A1(W17431), .A2(W8874), .ZN(W40215));
  NOR2X1 G4423 (.A1(W15907), .A2(W11695), .ZN(W21782));
  NOR2X1 G4424 (.A1(W7604), .A2(W6315), .ZN(O4705));
  NOR2X1 G4425 (.A1(W24739), .A2(W2849), .ZN(W29018));
  NOR2X1 G4426 (.A1(W22659), .A2(W7250), .ZN(O10723));
  NOR2X1 G4427 (.A1(W6481), .A2(W3996), .ZN(W10690));
  NOR2X1 G4428 (.A1(W9021), .A2(W12685), .ZN(W21779));
  NOR2X1 G4429 (.A1(W27), .A2(W23918), .ZN(W29015));
  NOR2X1 G4430 (.A1(W38877), .A2(I1367), .ZN(O10730));
  NOR2X1 G4431 (.A1(W19475), .A2(W17699), .ZN(W21781));
  NOR2X1 G4432 (.A1(W7928), .A2(W5392), .ZN(W10654));
  NOR2X1 G4433 (.A1(W21412), .A2(W39229), .ZN(W40192));
  NOR2X1 G4434 (.A1(W3537), .A2(I483), .ZN(O423));
  NOR2X1 G4435 (.A1(W28348), .A2(W11817), .ZN(O4703));
  NOR2X1 G4436 (.A1(W2683), .A2(W7009), .ZN(W29011));
  NOR2X1 G4437 (.A1(W4581), .A2(W23120), .ZN(O4700));
  NOR2X1 G4438 (.A1(W2091), .A2(W5641), .ZN(O4699));
  NOR2X1 G4439 (.A1(W8214), .A2(W4514), .ZN(W10675));
  NOR2X1 G4440 (.A1(W9737), .A2(W8005), .ZN(W10623));
  NOR2X1 G4441 (.A1(W4865), .A2(W31899), .ZN(O10765));
  NOR2X1 G4442 (.A1(W14282), .A2(I932), .ZN(W28994));
  NOR2X1 G4443 (.A1(W39421), .A2(W22332), .ZN(O10768));
  NOR2X1 G4444 (.A1(W5934), .A2(W3371), .ZN(W10630));
  NOR2X1 G4445 (.A1(W8750), .A2(W2434), .ZN(W10629));
  NOR2X1 G4446 (.A1(W7074), .A2(W4033), .ZN(W10627));
  NOR2X1 G4447 (.A1(W12512), .A2(W13172), .ZN(O4696));
  NOR2X1 G4448 (.A1(W1814), .A2(W536), .ZN(W10624));
  NOR2X1 G4449 (.A1(W9091), .A2(W8764), .ZN(W10634));
  NOR2X1 G4450 (.A1(W1041), .A2(W16738), .ZN(O10772));
  NOR2X1 G4451 (.A1(W9017), .A2(W3778), .ZN(W10621));
  NOR2X1 G4452 (.A1(W173), .A2(I1856), .ZN(O10775));
  NOR2X1 G4453 (.A1(W11239), .A2(W13515), .ZN(W28990));
  NOR2X1 G4454 (.A1(W806), .A2(W7686), .ZN(W10618));
  NOR2X1 G4455 (.A1(W7902), .A2(I36), .ZN(W10617));
  NOR2X1 G4456 (.A1(W5416), .A2(W3128), .ZN(W10616));
  NOR2X1 G4457 (.A1(W35125), .A2(W11898), .ZN(O10754));
  NOR2X1 G4458 (.A1(W1328), .A2(W6507), .ZN(W10652));
  NOR2X1 G4459 (.A1(W17139), .A2(W34767), .ZN(O10749));
  NOR2X1 G4460 (.A1(W11921), .A2(W6004), .ZN(O10751));
  NOR2X1 G4461 (.A1(W2356), .A2(W4591), .ZN(W10649));
  NOR2X1 G4462 (.A1(W18867), .A2(W14068), .ZN(W21792));
  NOR2X1 G4463 (.A1(W6935), .A2(W9381), .ZN(O416));
  NOR2X1 G4464 (.A1(W8391), .A2(W1727), .ZN(W40222));
  NOR2X1 G4465 (.A1(W14866), .A2(W16653), .ZN(O10753));
  NOR2X1 G4466 (.A1(W19250), .A2(W11844), .ZN(O2066));
  NOR2X1 G4467 (.A1(W28933), .A2(W11044), .ZN(W28999));
  NOR2X1 G4468 (.A1(W31435), .A2(W28574), .ZN(O10755));
  NOR2X1 G4469 (.A1(W5444), .A2(W8116), .ZN(W10641));
  NOR2X1 G4470 (.A1(W8279), .A2(W3161), .ZN(W10638));
  NOR2X1 G4471 (.A1(W31743), .A2(W34255), .ZN(W40234));
  NOR2X1 G4472 (.A1(W16701), .A2(W12393), .ZN(O10762));
  NOR2X1 G4473 (.A1(W38130), .A2(I227), .ZN(W40238));
  NOR2X1 G4474 (.A1(W16616), .A2(W116), .ZN(W19579));
  NOR2X1 G4475 (.A1(W26475), .A2(W4224), .ZN(W33541));
  NOR2X1 G4476 (.A1(W26612), .A2(W30842), .ZN(O6751));
  NOR2X1 G4477 (.A1(W17827), .A2(W1661), .ZN(O5711));
  NOR2X1 G4478 (.A1(W1885), .A2(W6858), .ZN(W19574));
  NOR2X1 G4479 (.A1(W1185), .A2(I1128), .ZN(W19575));
  NOR2X1 G4480 (.A1(W9396), .A2(W15507), .ZN(W19577));
  NOR2X1 G4481 (.A1(W2985), .A2(I1763), .ZN(W31260));
  NOR2X1 G4482 (.A1(W8789), .A2(W31609), .ZN(W33553));
  NOR2X1 G4483 (.A1(W10524), .A2(W9188), .ZN(W19571));
  NOR2X1 G4484 (.A1(W17227), .A2(W15797), .ZN(O1374));
  NOR2X1 G4485 (.A1(I945), .A2(W12828), .ZN(W17336));
  NOR2X1 G4486 (.A1(W22897), .A2(W24566), .ZN(W31255));
  NOR2X1 G4487 (.A1(W10699), .A2(W13219), .ZN(W33560));
  NOR2X1 G4488 (.A1(W21057), .A2(W22625), .ZN(O6761));
  NOR2X1 G4489 (.A1(W24983), .A2(W23766), .ZN(O6762));
  NOR2X1 G4490 (.A1(W15062), .A2(W5044), .ZN(W33563));
  NOR2X1 G4491 (.A1(W18658), .A2(W23361), .ZN(W33570));
  NOR2X1 G4492 (.A1(W4756), .A2(W1594), .ZN(W19570));
  NOR2X1 G4493 (.A1(W5845), .A2(W17149), .ZN(W17367));
  NOR2X1 G4494 (.A1(W6305), .A2(W5110), .ZN(W17366));
  NOR2X1 G4495 (.A1(W12453), .A2(W16289), .ZN(W17365));
  NOR2X1 G4496 (.A1(W7865), .A2(W9400), .ZN(W17364));
  NOR2X1 G4497 (.A1(W984), .A2(W212), .ZN(W31265));
  NOR2X1 G4498 (.A1(W171), .A2(W18790), .ZN(O6745));
  NOR2X1 G4499 (.A1(W25193), .A2(W29095), .ZN(W33532));
  NOR2X1 G4500 (.A1(W4116), .A2(W17452), .ZN(W19569));
  NOR2X1 G4501 (.A1(W28693), .A2(W12622), .ZN(W33572));
  NOR2X1 G4502 (.A1(I1303), .A2(W5972), .ZN(W17358));
  NOR2X1 G4503 (.A1(W7286), .A2(W6181), .ZN(W17357));
  NOR2X1 G4504 (.A1(W6450), .A2(W13857), .ZN(W17356));
  NOR2X1 G4505 (.A1(W26838), .A2(I1385), .ZN(W33536));
  NOR2X1 G4506 (.A1(W11420), .A2(W30097), .ZN(O6748));
  NOR2X1 G4507 (.A1(W15834), .A2(W10515), .ZN(W33538));
  NOR2X1 G4508 (.A1(I150), .A2(W12441), .ZN(W17352));
  NOR2X1 G4509 (.A1(W6648), .A2(W5962), .ZN(W19594));
  NOR2X1 G4510 (.A1(W23295), .A2(W4130), .ZN(W33591));
  NOR2X1 G4511 (.A1(W14929), .A2(W13749), .ZN(O6774));
  NOR2X1 G4512 (.A1(W728), .A2(W4703), .ZN(O1367));
  NOR2X1 G4513 (.A1(W1485), .A2(I309), .ZN(O6776));
  NOR2X1 G4514 (.A1(W13418), .A2(W2023), .ZN(W17303));
  NOR2X1 G4515 (.A1(W12973), .A2(W9789), .ZN(O6777));
  NOR2X1 G4516 (.A1(W25219), .A2(W24350), .ZN(W31243));
  NOR2X1 G4517 (.A1(W17293), .A2(W14417), .ZN(O1364));
  NOR2X1 G4518 (.A1(W2780), .A2(W10402), .ZN(O1368));
  NOR2X1 G4519 (.A1(W9792), .A2(W24058), .ZN(W33604));
  NOR2X1 G4520 (.A1(W11296), .A2(W13699), .ZN(W17297));
  NOR2X1 G4521 (.A1(W4607), .A2(I1339), .ZN(W17295));
  NOR2X1 G4522 (.A1(W16249), .A2(W10697), .ZN(O1362));
  NOR2X1 G4523 (.A1(W33149), .A2(W5319), .ZN(W33607));
  NOR2X1 G4524 (.A1(W12783), .A2(W10255), .ZN(W17292));
  NOR2X1 G4525 (.A1(W22784), .A2(W29078), .ZN(W33608));
  NOR2X1 G4526 (.A1(W2460), .A2(W16906), .ZN(W19596));
  NOR2X1 G4527 (.A1(W13626), .A2(W25804), .ZN(O5709));
  NOR2X1 G4528 (.A1(W13324), .A2(W5507), .ZN(W19584));
  NOR2X1 G4529 (.A1(W1700), .A2(W6141), .ZN(W17326));
  NOR2X1 G4530 (.A1(W13510), .A2(W10866), .ZN(W17324));
  NOR2X1 G4531 (.A1(W5698), .A2(W31108), .ZN(W33576));
  NOR2X1 G4532 (.A1(W7702), .A2(W944), .ZN(W17322));
  NOR2X1 G4533 (.A1(W6363), .A2(W3495), .ZN(O1803));
  NOR2X1 G4534 (.A1(W17355), .A2(W9480), .ZN(W33578));
  NOR2X1 G4535 (.A1(W3911), .A2(W2175), .ZN(O6767));
  NOR2X1 G4536 (.A1(W26136), .A2(W632), .ZN(W31266));
  NOR2X1 G4537 (.A1(W12679), .A2(W7781), .ZN(W33581));
  NOR2X1 G4538 (.A1(W31513), .A2(W19321), .ZN(W33583));
  NOR2X1 G4539 (.A1(W25297), .A2(W15902), .ZN(W31249));
  NOR2X1 G4540 (.A1(W8508), .A2(W24355), .ZN(W31248));
  NOR2X1 G4541 (.A1(W9981), .A2(W3868), .ZN(W17312));
  NOR2X1 G4542 (.A1(W26108), .A2(W9472), .ZN(W31246));
  NOR2X1 G4543 (.A1(W1533), .A2(W6809), .ZN(W17310));
  NOR2X1 G4544 (.A1(W25379), .A2(W17262), .ZN(W33477));
  NOR2X1 G4545 (.A1(W8819), .A2(W26062), .ZN(O6719));
  NOR2X1 G4546 (.A1(W1992), .A2(W4531), .ZN(W17423));
  NOR2X1 G4547 (.A1(W1938), .A2(I1273), .ZN(W17422));
  NOR2X1 G4548 (.A1(W28096), .A2(W21606), .ZN(W33473));
  NOR2X1 G4549 (.A1(W7174), .A2(W33257), .ZN(O6720));
  NOR2X1 G4550 (.A1(I947), .A2(W10427), .ZN(W17419));
  NOR2X1 G4551 (.A1(W5771), .A2(W14288), .ZN(O6721));
  NOR2X1 G4552 (.A1(W3663), .A2(W12925), .ZN(W17417));
  NOR2X1 G4553 (.A1(W9336), .A2(W671), .ZN(W33470));
  NOR2X1 G4554 (.A1(W17690), .A2(W1108), .ZN(W19550));
  NOR2X1 G4555 (.A1(W7169), .A2(W6447), .ZN(O6724));
  NOR2X1 G4556 (.A1(W7847), .A2(W3899), .ZN(W19551));
  NOR2X1 G4557 (.A1(W1946), .A2(W13056), .ZN(O1384));
  NOR2X1 G4558 (.A1(W2003), .A2(W3208), .ZN(W33483));
  NOR2X1 G4559 (.A1(W8156), .A2(I1483), .ZN(W17410));
  NOR2X1 G4560 (.A1(W6979), .A2(W14320), .ZN(W17409));
  NOR2X1 G4561 (.A1(W5425), .A2(W20474), .ZN(W31279));
  NOR2X1 G4562 (.A1(W2893), .A2(W28331), .ZN(W31286));
  NOR2X1 G4563 (.A1(W9252), .A2(W14529), .ZN(W17442));
  NOR2X1 G4564 (.A1(W15931), .A2(W6827), .ZN(W19543));
  NOR2X1 G4565 (.A1(W7250), .A2(W8303), .ZN(W17440));
  NOR2X1 G4566 (.A1(W6013), .A2(W7715), .ZN(O1390));
  NOR2X1 G4567 (.A1(W6173), .A2(W7358), .ZN(W31287));
  NOR2X1 G4568 (.A1(W2673), .A2(W13612), .ZN(W19545));
  NOR2X1 G4569 (.A1(W2941), .A2(W23418), .ZN(O6715));
  NOR2X1 G4570 (.A1(W7454), .A2(W8547), .ZN(W17435));
  NOR2X1 G4571 (.A1(W20875), .A2(W6820), .ZN(W31277));
  NOR2X1 G4572 (.A1(W14860), .A2(W19506), .ZN(O5720));
  NOR2X1 G4573 (.A1(W15185), .A2(I623), .ZN(W17432));
  NOR2X1 G4574 (.A1(W4600), .A2(W25886), .ZN(W31283));
  NOR2X1 G4575 (.A1(I1386), .A2(W24427), .ZN(W33469));
  NOR2X1 G4576 (.A1(I1031), .A2(I713), .ZN(W17429));
  NOR2X1 G4577 (.A1(W7280), .A2(W130), .ZN(O1387));
  NOR2X1 G4578 (.A1(I1670), .A2(W2761), .ZN(W17427));
  NOR2X1 G4579 (.A1(W2320), .A2(W15782), .ZN(W17378));
  NOR2X1 G4580 (.A1(I904), .A2(W12735), .ZN(W33505));
  NOR2X1 G4581 (.A1(W15168), .A2(W7399), .ZN(W19561));
  NOR2X1 G4582 (.A1(W6768), .A2(W9275), .ZN(W17385));
  NOR2X1 G4583 (.A1(W14129), .A2(W6050), .ZN(W17384));
  NOR2X1 G4584 (.A1(W6274), .A2(W6780), .ZN(W19563));
  NOR2X1 G4585 (.A1(W22063), .A2(W20745), .ZN(W33515));
  NOR2X1 G4586 (.A1(I968), .A2(W534), .ZN(W17380));
  NOR2X1 G4587 (.A1(I1725), .A2(W6881), .ZN(W19564));
  NOR2X1 G4588 (.A1(W29262), .A2(W22445), .ZN(O6734));
  NOR2X1 G4589 (.A1(W2591), .A2(W32592), .ZN(W33519));
  NOR2X1 G4590 (.A1(W17966), .A2(W10734), .ZN(W33521));
  NOR2X1 G4591 (.A1(W23772), .A2(W27544), .ZN(O6743));
  NOR2X1 G4592 (.A1(W2053), .A2(W17151), .ZN(W17373));
  NOR2X1 G4593 (.A1(W14304), .A2(W15220), .ZN(W17372));
  NOR2X1 G4594 (.A1(W4547), .A2(W11450), .ZN(W33524));
  NOR2X1 G4595 (.A1(W13495), .A2(W8776), .ZN(O5712));
  NOR2X1 G4596 (.A1(W12109), .A2(W9318), .ZN(O1379));
  NOR2X1 G4597 (.A1(W13163), .A2(W11640), .ZN(W19556));
  NOR2X1 G4598 (.A1(W5010), .A2(W5766), .ZN(W31275));
  NOR2X1 G4599 (.A1(W13943), .A2(W5293), .ZN(O1383));
  NOR2X1 G4600 (.A1(W16035), .A2(W26063), .ZN(W33492));
  NOR2X1 G4601 (.A1(W16876), .A2(W30412), .ZN(O6730));
  NOR2X1 G4602 (.A1(W15679), .A2(W16650), .ZN(O6731));
  NOR2X1 G4603 (.A1(W15122), .A2(W481), .ZN(W17400));
  NOR2X1 G4604 (.A1(W14456), .A2(W14258), .ZN(W17399));
  NOR2X1 G4605 (.A1(W4225), .A2(W6088), .ZN(W17398));
  NOR2X1 G4606 (.A1(W24356), .A2(W17200), .ZN(O6783));
  NOR2X1 G4607 (.A1(W5623), .A2(W11619), .ZN(W17395));
  NOR2X1 G4608 (.A1(W258), .A2(W10640), .ZN(W19558));
  NOR2X1 G4609 (.A1(W7507), .A2(I1542), .ZN(W17393));
  NOR2X1 G4610 (.A1(W713), .A2(W4283), .ZN(W17392));
  NOR2X1 G4611 (.A1(W17077), .A2(W7776), .ZN(O5714));
  NOR2X1 G4612 (.A1(W30900), .A2(W6600), .ZN(W33500));
  NOR2X1 G4613 (.A1(W6560), .A2(W12646), .ZN(O1799));
  NOR2X1 G4614 (.A1(W12133), .A2(I1835), .ZN(W33721));
  NOR2X1 G4615 (.A1(W3506), .A2(W15786), .ZN(O1812));
  NOR2X1 G4616 (.A1(W9010), .A2(W8073), .ZN(O1341));
  NOR2X1 G4617 (.A1(W4198), .A2(W8935), .ZN(W17184));
  NOR2X1 G4618 (.A1(W15375), .A2(W3391), .ZN(W17183));
  NOR2X1 G4619 (.A1(W4409), .A2(W410), .ZN(W17182));
  NOR2X1 G4620 (.A1(W439), .A2(W19161), .ZN(O1813));
  NOR2X1 G4621 (.A1(W11058), .A2(W8507), .ZN(W17180));
  NOR2X1 G4622 (.A1(W2333), .A2(W2284), .ZN(W31194));
  NOR2X1 G4623 (.A1(W13780), .A2(I1266), .ZN(W17187));
  NOR2X1 G4624 (.A1(W19563), .A2(W12919), .ZN(W19637));
  NOR2X1 G4625 (.A1(W3481), .A2(I1865), .ZN(W17176));
  NOR2X1 G4626 (.A1(I1106), .A2(W10086), .ZN(W19638));
  NOR2X1 G4627 (.A1(W9070), .A2(W9336), .ZN(W17174));
  NOR2X1 G4628 (.A1(W13461), .A2(W14556), .ZN(W17173));
  NOR2X1 G4629 (.A1(W10622), .A2(W4479), .ZN(W17172));
  NOR2X1 G4630 (.A1(W30077), .A2(W8835), .ZN(W33724));
  NOR2X1 G4631 (.A1(W5045), .A2(W12328), .ZN(O1338));
  NOR2X1 G4632 (.A1(W16213), .A2(W256), .ZN(W17198));
  NOR2X1 G4633 (.A1(W15698), .A2(W15209), .ZN(W17208));
  NOR2X1 G4634 (.A1(W1570), .A2(W11477), .ZN(W17207));
  NOR2X1 G4635 (.A1(W13394), .A2(W30759), .ZN(O6839));
  NOR2X1 G4636 (.A1(W5901), .A2(W12011), .ZN(W19627));
  NOR2X1 G4637 (.A1(W15470), .A2(W2693), .ZN(O5689));
  NOR2X1 G4638 (.A1(W28081), .A2(W1474), .ZN(W31205));
  NOR2X1 G4639 (.A1(W3767), .A2(W1316), .ZN(W17200));
  NOR2X1 G4640 (.A1(W3779), .A2(W20283), .ZN(O6842));
  NOR2X1 G4641 (.A1(W13519), .A2(I212), .ZN(W17169));
  NOR2X1 G4642 (.A1(W16285), .A2(W3609), .ZN(W17197));
  NOR2X1 G4643 (.A1(W8807), .A2(W14149), .ZN(W17196));
  NOR2X1 G4644 (.A1(W17574), .A2(W7232), .ZN(W31197));
  NOR2X1 G4645 (.A1(W11567), .A2(W4620), .ZN(W17192));
  NOR2X1 G4646 (.A1(W15285), .A2(W7051), .ZN(W17190));
  NOR2X1 G4647 (.A1(W10402), .A2(W16446), .ZN(W17189));
  NOR2X1 G4648 (.A1(W13285), .A2(W7293), .ZN(W33715));
  NOR2X1 G4649 (.A1(W12309), .A2(W9215), .ZN(W19652));
  NOR2X1 G4650 (.A1(W15310), .A2(I423), .ZN(W33748));
  NOR2X1 G4651 (.A1(W6548), .A2(W8625), .ZN(W19650));
  NOR2X1 G4652 (.A1(W7508), .A2(W11401), .ZN(O1333));
  NOR2X1 G4653 (.A1(W22792), .A2(W24045), .ZN(W33756));
  NOR2X1 G4654 (.A1(W7091), .A2(W28837), .ZN(W33760));
  NOR2X1 G4655 (.A1(W7777), .A2(W14236), .ZN(W19651));
  NOR2X1 G4656 (.A1(I317), .A2(W302), .ZN(W17142));
  NOR2X1 G4657 (.A1(W9694), .A2(W3520), .ZN(O1331));
  NOR2X1 G4658 (.A1(W11321), .A2(W2571), .ZN(W19647));
  NOR2X1 G4659 (.A1(W12298), .A2(W7290), .ZN(W19653));
  NOR2X1 G4660 (.A1(W9864), .A2(W9424), .ZN(O6869));
  NOR2X1 G4661 (.A1(W7417), .A2(W4413), .ZN(W33766));
  NOR2X1 G4662 (.A1(W4369), .A2(W6715), .ZN(W33769));
  NOR2X1 G4663 (.A1(W7142), .A2(W10042), .ZN(O1815));
  NOR2X1 G4664 (.A1(W11373), .A2(W14159), .ZN(O1330));
  NOR2X1 G4665 (.A1(I257), .A2(W5038), .ZN(W19655));
  NOR2X1 G4666 (.A1(W23829), .A2(W7697), .ZN(W33773));
  NOR2X1 G4667 (.A1(W2414), .A2(W74), .ZN(W31191));
  NOR2X1 G4668 (.A1(W2720), .A2(W753), .ZN(W17168));
  NOR2X1 G4669 (.A1(W9721), .A2(W9696), .ZN(W19639));
  NOR2X1 G4670 (.A1(W57), .A2(I1861), .ZN(W17166));
  NOR2X1 G4671 (.A1(W14543), .A2(W14827), .ZN(O5681));
  NOR2X1 G4672 (.A1(W9447), .A2(W4858), .ZN(W17164));
  NOR2X1 G4673 (.A1(W5354), .A2(W25823), .ZN(O5680));
  NOR2X1 G4674 (.A1(W17725), .A2(W931), .ZN(W19642));
  NOR2X1 G4675 (.A1(W10781), .A2(W1452), .ZN(W33734));
  NOR2X1 G4676 (.A1(W4657), .A2(I1330), .ZN(W17209));
  NOR2X1 G4677 (.A1(W15701), .A2(W8176), .ZN(W17159));
  NOR2X1 G4678 (.A1(W19601), .A2(W18064), .ZN(W31186));
  NOR2X1 G4679 (.A1(W12067), .A2(W19658), .ZN(O5675));
  NOR2X1 G4680 (.A1(W9670), .A2(W11699), .ZN(W33743));
  NOR2X1 G4681 (.A1(W8333), .A2(W6156), .ZN(W17154));
  NOR2X1 G4682 (.A1(W7011), .A2(I86), .ZN(W17153));
  NOR2X1 G4683 (.A1(W10811), .A2(W23575), .ZN(O6863));
  NOR2X1 G4684 (.A1(W25208), .A2(W16097), .ZN(O5700));
  NOR2X1 G4685 (.A1(W21058), .A2(W474), .ZN(W31233));
  NOR2X1 G4686 (.A1(W25700), .A2(W9300), .ZN(O6803));
  NOR2X1 G4687 (.A1(W2380), .A2(W16816), .ZN(O5702));
  NOR2X1 G4688 (.A1(W17563), .A2(W25217), .ZN(O6805));
  NOR2X1 G4689 (.A1(W2516), .A2(W11392), .ZN(W17263));
  NOR2X1 G4690 (.A1(W10822), .A2(W11129), .ZN(W17262));
  NOR2X1 G4691 (.A1(W21191), .A2(I1577), .ZN(W33643));
  NOR2X1 G4692 (.A1(W4435), .A2(W14695), .ZN(W19606));
  NOR2X1 G4693 (.A1(W2780), .A2(W11859), .ZN(O6798));
  NOR2X1 G4694 (.A1(I856), .A2(W3336), .ZN(O1358));
  NOR2X1 G4695 (.A1(W6055), .A2(W8489), .ZN(W31227));
  NOR2X1 G4696 (.A1(W3810), .A2(W2521), .ZN(W17256));
  NOR2X1 G4697 (.A1(W29778), .A2(W9822), .ZN(O6810));
  NOR2X1 G4698 (.A1(W22886), .A2(W32909), .ZN(W33651));
  NOR2X1 G4699 (.A1(W18243), .A2(W17157), .ZN(W33653));
  NOR2X1 G4700 (.A1(W13906), .A2(W3073), .ZN(O6812));
  NOR2X1 G4701 (.A1(W1124), .A2(W4587), .ZN(O6813));
  NOR2X1 G4702 (.A1(W26338), .A2(W28508), .ZN(O6789));
  NOR2X1 G4703 (.A1(W6898), .A2(W20997), .ZN(W31241));
  NOR2X1 G4704 (.A1(W16006), .A2(W21838), .ZN(O6785));
  NOR2X1 G4705 (.A1(I1566), .A2(W26034), .ZN(O6787));
  NOR2X1 G4706 (.A1(W6492), .A2(W7124), .ZN(W17283));
  NOR2X1 G4707 (.A1(W14767), .A2(W7180), .ZN(W17282));
  NOR2X1 G4708 (.A1(W1736), .A2(W11911), .ZN(W17281));
  NOR2X1 G4709 (.A1(I673), .A2(W18776), .ZN(W19600));
  NOR2X1 G4710 (.A1(W10368), .A2(W4351), .ZN(O1361));
  NOR2X1 G4711 (.A1(I953), .A2(I771), .ZN(W19611));
  NOR2X1 G4712 (.A1(W20035), .A2(W29163), .ZN(O6790));
  NOR2X1 G4713 (.A1(W26065), .A2(W6105), .ZN(O6791));
  NOR2X1 G4714 (.A1(W2650), .A2(W6388), .ZN(O5704));
  NOR2X1 G4715 (.A1(I439), .A2(W1743), .ZN(O1360));
  NOR2X1 G4716 (.A1(W20588), .A2(W1200), .ZN(O6793));
  NOR2X1 G4717 (.A1(W8130), .A2(W29389), .ZN(O6795));
  NOR2X1 G4718 (.A1(W3780), .A2(W9166), .ZN(W17269));
  NOR2X1 G4719 (.A1(W14251), .A2(W11024), .ZN(W17218));
  NOR2X1 G4720 (.A1(W6229), .A2(W8299), .ZN(W17226));
  NOR2X1 G4721 (.A1(W29808), .A2(W3258), .ZN(W33681));
  NOR2X1 G4722 (.A1(W29882), .A2(W1025), .ZN(O6831));
  NOR2X1 G4723 (.A1(W10257), .A2(W13681), .ZN(O1810));
  NOR2X1 G4724 (.A1(W16556), .A2(W747), .ZN(W19622));
  NOR2X1 G4725 (.A1(W1833), .A2(W5425), .ZN(W17221));
  NOR2X1 G4726 (.A1(W8662), .A2(W23660), .ZN(W33691));
  NOR2X1 G4727 (.A1(W4348), .A2(W13446), .ZN(W17219));
  NOR2X1 G4728 (.A1(I1992), .A2(W16468), .ZN(W17227));
  NOR2X1 G4729 (.A1(W29145), .A2(W27948), .ZN(W33694));
  NOR2X1 G4730 (.A1(I626), .A2(W2953), .ZN(O1350));
  NOR2X1 G4731 (.A1(W789), .A2(W21811), .ZN(O5690));
  NOR2X1 G4732 (.A1(W15383), .A2(W16173), .ZN(O1349));
  NOR2X1 G4733 (.A1(W5304), .A2(W2551), .ZN(W17213));
  NOR2X1 G4734 (.A1(W9704), .A2(W15157), .ZN(W17212));
  NOR2X1 G4735 (.A1(W25579), .A2(W20270), .ZN(W33698));
  NOR2X1 G4736 (.A1(W365), .A2(W13914), .ZN(W19624));
  NOR2X1 G4737 (.A1(W11392), .A2(W13123), .ZN(W17236));
  NOR2X1 G4738 (.A1(W19055), .A2(W3766), .ZN(W31219));
  NOR2X1 G4739 (.A1(W792), .A2(W8554), .ZN(W17245));
  NOR2X1 G4740 (.A1(W21640), .A2(W18100), .ZN(O6818));
  NOR2X1 G4741 (.A1(W7128), .A2(W9881), .ZN(O1352));
  NOR2X1 G4742 (.A1(W16141), .A2(W7781), .ZN(O5694));
  NOR2X1 G4743 (.A1(W174), .A2(I1939), .ZN(W17240));
  NOR2X1 G4744 (.A1(W31123), .A2(W30298), .ZN(W33667));
  NOR2X1 G4745 (.A1(W19041), .A2(W10995), .ZN(W19616));
  NOR2X1 G4746 (.A1(W10203), .A2(W8004), .ZN(W17443));
  NOR2X1 G4747 (.A1(W1817), .A2(W11421), .ZN(W17235));
  NOR2X1 G4748 (.A1(W16724), .A2(W17366), .ZN(W19618));
  NOR2X1 G4749 (.A1(W24225), .A2(W15870), .ZN(O6824));
  NOR2X1 G4750 (.A1(W27035), .A2(W25807), .ZN(O6828));
  NOR2X1 G4751 (.A1(W3738), .A2(W2014), .ZN(W17230));
  NOR2X1 G4752 (.A1(W962), .A2(W13950), .ZN(W33679));
  NOR2X1 G4753 (.A1(I1818), .A2(W7999), .ZN(W19620));
  NOR2X1 G4754 (.A1(W12758), .A2(W17603), .ZN(W17657));
  NOR2X1 G4755 (.A1(W3497), .A2(W18990), .ZN(W33216));
  NOR2X1 G4756 (.A1(W17808), .A2(W31334), .ZN(W33218));
  NOR2X1 G4757 (.A1(W4370), .A2(W22508), .ZN(O6600));
  NOR2X1 G4758 (.A1(W11478), .A2(W4787), .ZN(W33221));
  NOR2X1 G4759 (.A1(W16569), .A2(I358), .ZN(W17662));
  NOR2X1 G4760 (.A1(W16814), .A2(W6719), .ZN(W33224));
  NOR2X1 G4761 (.A1(W17067), .A2(W12621), .ZN(W17659));
  NOR2X1 G4762 (.A1(W16611), .A2(W15976), .ZN(O1425));
  NOR2X1 G4763 (.A1(W10239), .A2(W20074), .ZN(O6598));
  NOR2X1 G4764 (.A1(W7993), .A2(W13023), .ZN(W33226));
  NOR2X1 G4765 (.A1(W3836), .A2(W11522), .ZN(W19463));
  NOR2X1 G4766 (.A1(W6087), .A2(I1912), .ZN(W19464));
  NOR2X1 G4767 (.A1(W25797), .A2(W13763), .ZN(O6606));
  NOR2X1 G4768 (.A1(W1612), .A2(W20875), .ZN(W33231));
  NOR2X1 G4769 (.A1(W14312), .A2(W16733), .ZN(W19465));
  NOR2X1 G4770 (.A1(W32258), .A2(W5986), .ZN(O6609));
  NOR2X1 G4771 (.A1(W15098), .A2(W18552), .ZN(W19466));
  NOR2X1 G4772 (.A1(W22365), .A2(W625), .ZN(W33201));
  NOR2X1 G4773 (.A1(W782), .A2(W23225), .ZN(W33184));
  NOR2X1 G4774 (.A1(W1389), .A2(W27551), .ZN(O6584));
  NOR2X1 G4775 (.A1(W27637), .A2(W17220), .ZN(W33188));
  NOR2X1 G4776 (.A1(W7171), .A2(W5413), .ZN(W17682));
  NOR2X1 G4777 (.A1(W27556), .A2(W18360), .ZN(O6585));
  NOR2X1 G4778 (.A1(W23576), .A2(W15798), .ZN(O6588));
  NOR2X1 G4779 (.A1(W23819), .A2(W26405), .ZN(O6589));
  NOR2X1 G4780 (.A1(W27589), .A2(I1483), .ZN(W31372));
  NOR2X1 G4781 (.A1(I546), .A2(W832), .ZN(O1421));
  NOR2X1 G4782 (.A1(W3806), .A2(W11782), .ZN(O1428));
  NOR2X1 G4783 (.A1(W2589), .A2(W1238), .ZN(O6592));
  NOR2X1 G4784 (.A1(W26325), .A2(W8022), .ZN(O6596));
  NOR2X1 G4785 (.A1(W28960), .A2(W3935), .ZN(O6597));
  NOR2X1 G4786 (.A1(W11765), .A2(W11111), .ZN(W19461));
  NOR2X1 G4787 (.A1(W17559), .A2(W22570), .ZN(W33212));
  NOR2X1 G4788 (.A1(W31544), .A2(W30151), .ZN(W33213));
  NOR2X1 G4789 (.A1(W689), .A2(W4702), .ZN(W33275));
  NOR2X1 G4790 (.A1(W781), .A2(W15756), .ZN(W31354));
  NOR2X1 G4791 (.A1(W5114), .A2(W13686), .ZN(W17624));
  NOR2X1 G4792 (.A1(W10327), .A2(W14265), .ZN(W17622));
  NOR2X1 G4793 (.A1(W1581), .A2(I421), .ZN(W17620));
  NOR2X1 G4794 (.A1(W2064), .A2(W4352), .ZN(W17619));
  NOR2X1 G4795 (.A1(W23161), .A2(W23565), .ZN(W31350));
  NOR2X1 G4796 (.A1(W12018), .A2(I941), .ZN(W17617));
  NOR2X1 G4797 (.A1(W31128), .A2(W20969), .ZN(W31349));
  NOR2X1 G4798 (.A1(W8803), .A2(W503), .ZN(O5750));
  NOR2X1 G4799 (.A1(W14063), .A2(W16236), .ZN(W19482));
  NOR2X1 G4800 (.A1(W10317), .A2(W8592), .ZN(W17612));
  NOR2X1 G4801 (.A1(W9983), .A2(W16905), .ZN(W17611));
  NOR2X1 G4802 (.A1(W11711), .A2(I956), .ZN(W17610));
  NOR2X1 G4803 (.A1(W17363), .A2(W16179), .ZN(W17609));
  NOR2X1 G4804 (.A1(W27311), .A2(W30140), .ZN(W33278));
  NOR2X1 G4805 (.A1(W5076), .A2(W8712), .ZN(W19486));
  NOR2X1 G4806 (.A1(W6174), .A2(W15521), .ZN(W17604));
  NOR2X1 G4807 (.A1(W6908), .A2(W32621), .ZN(O6623));
  NOR2X1 G4808 (.A1(W5463), .A2(W15287), .ZN(W17647));
  NOR2X1 G4809 (.A1(W10317), .A2(W15001), .ZN(W17645));
  NOR2X1 G4810 (.A1(W33153), .A2(W23832), .ZN(O6621));
  NOR2X1 G4811 (.A1(W11226), .A2(W6457), .ZN(W17642));
  NOR2X1 G4812 (.A1(W6990), .A2(W21401), .ZN(W33252));
  NOR2X1 G4813 (.A1(W23210), .A2(W23502), .ZN(W31361));
  NOR2X1 G4814 (.A1(W848), .A2(W5999), .ZN(W19471));
  NOR2X1 G4815 (.A1(I859), .A2(W7628), .ZN(W17637));
  NOR2X1 G4816 (.A1(W15804), .A2(W15003), .ZN(W17687));
  NOR2X1 G4817 (.A1(W18369), .A2(W8812), .ZN(W19472));
  NOR2X1 G4818 (.A1(I9), .A2(W1700), .ZN(W17634));
  NOR2X1 G4819 (.A1(W11670), .A2(W6454), .ZN(W17632));
  NOR2X1 G4820 (.A1(W5163), .A2(W5756), .ZN(W33263));
  NOR2X1 G4821 (.A1(W14326), .A2(W15481), .ZN(W19475));
  NOR2X1 G4822 (.A1(W25548), .A2(W17696), .ZN(W33265));
  NOR2X1 G4823 (.A1(W19792), .A2(W16098), .ZN(O6627));
  NOR2X1 G4824 (.A1(W17307), .A2(W2429), .ZN(W17735));
  NOR2X1 G4825 (.A1(W30710), .A2(W8964), .ZN(W33126));
  NOR2X1 G4826 (.A1(W12965), .A2(I304), .ZN(W19438));
  NOR2X1 G4827 (.A1(W16884), .A2(W748), .ZN(W19439));
  NOR2X1 G4828 (.A1(W1305), .A2(W1578), .ZN(W17740));
  NOR2X1 G4829 (.A1(W2890), .A2(W1714), .ZN(W17739));
  NOR2X1 G4830 (.A1(W29857), .A2(W15356), .ZN(O6560));
  NOR2X1 G4831 (.A1(W9262), .A2(W26136), .ZN(W33132));
  NOR2X1 G4832 (.A1(W20728), .A2(W191), .ZN(O5765));
  NOR2X1 G4833 (.A1(W17946), .A2(W987), .ZN(O6557));
  NOR2X1 G4834 (.A1(W1050), .A2(I1875), .ZN(W17734));
  NOR2X1 G4835 (.A1(W31963), .A2(W2691), .ZN(O6561));
  NOR2X1 G4836 (.A1(W10842), .A2(W9874), .ZN(W17731));
  NOR2X1 G4837 (.A1(W27414), .A2(W27482), .ZN(O6563));
  NOR2X1 G4838 (.A1(W9712), .A2(W12479), .ZN(W17729));
  NOR2X1 G4839 (.A1(W11351), .A2(W30499), .ZN(W31388));
  NOR2X1 G4840 (.A1(W13454), .A2(W19114), .ZN(W19443));
  NOR2X1 G4841 (.A1(W29243), .A2(W16058), .ZN(W33140));
  NOR2X1 G4842 (.A1(W7490), .A2(W16138), .ZN(W17752));
  NOR2X1 G4843 (.A1(W31474), .A2(W32790), .ZN(O6549));
  NOR2X1 G4844 (.A1(W23571), .A2(W28477), .ZN(O6550));
  NOR2X1 G4845 (.A1(W26404), .A2(W28503), .ZN(O6551));
  NOR2X1 G4846 (.A1(I928), .A2(W429), .ZN(W17757));
  NOR2X1 G4847 (.A1(W9649), .A2(W13939), .ZN(W19434));
  NOR2X1 G4848 (.A1(I11), .A2(W445), .ZN(W17755));
  NOR2X1 G4849 (.A1(W8191), .A2(I1364), .ZN(W19435));
  NOR2X1 G4850 (.A1(W2419), .A2(W4735), .ZN(O6553));
  NOR2X1 G4851 (.A1(I315), .A2(I1550), .ZN(W17725));
  NOR2X1 G4852 (.A1(W14722), .A2(W7465), .ZN(W31394));
  NOR2X1 G4853 (.A1(W5938), .A2(W4974), .ZN(W17750));
  NOR2X1 G4854 (.A1(W3524), .A2(W1730), .ZN(W17749));
  NOR2X1 G4855 (.A1(W25692), .A2(W4112), .ZN(W33121));
  NOR2X1 G4856 (.A1(W7911), .A2(W175), .ZN(W17747));
  NOR2X1 G4857 (.A1(W13334), .A2(W12111), .ZN(W17746));
  NOR2X1 G4858 (.A1(W27404), .A2(W30630), .ZN(W31392));
  NOR2X1 G4859 (.A1(W29561), .A2(W19551), .ZN(W33175));
  NOR2X1 G4860 (.A1(W2095), .A2(W4407), .ZN(W17707));
  NOR2X1 G4861 (.A1(W942), .A2(W9826), .ZN(W17706));
  NOR2X1 G4862 (.A1(W30753), .A2(W1575), .ZN(O5761));
  NOR2X1 G4863 (.A1(W10421), .A2(I992), .ZN(W17703));
  NOR2X1 G4864 (.A1(W4846), .A2(W26328), .ZN(O5760));
  NOR2X1 G4865 (.A1(W20830), .A2(W32526), .ZN(W33169));
  NOR2X1 G4866 (.A1(W10526), .A2(W13749), .ZN(W19454));
  NOR2X1 G4867 (.A1(W7519), .A2(W24352), .ZN(W31378));
  NOR2X1 G4868 (.A1(W15094), .A2(I418), .ZN(W19449));
  NOR2X1 G4869 (.A1(W12368), .A2(W2642), .ZN(W17696));
  NOR2X1 G4870 (.A1(W7445), .A2(W7520), .ZN(W17695));
  NOR2X1 G4871 (.A1(W25103), .A2(W1866), .ZN(O6579));
  NOR2X1 G4872 (.A1(W12065), .A2(I1442), .ZN(O6580));
  NOR2X1 G4873 (.A1(W17766), .A2(W6101), .ZN(O6581));
  NOR2X1 G4874 (.A1(I1650), .A2(W32688), .ZN(O6582));
  NOR2X1 G4875 (.A1(W20902), .A2(W30547), .ZN(W33182));
  NOR2X1 G4876 (.A1(W28811), .A2(W21593), .ZN(O6583));
  NOR2X1 G4877 (.A1(W16329), .A2(W10562), .ZN(O1777));
  NOR2X1 G4878 (.A1(W28212), .A2(W15785), .ZN(O6565));
  NOR2X1 G4879 (.A1(W24258), .A2(W21509), .ZN(W33146));
  NOR2X1 G4880 (.A1(W6316), .A2(W15820), .ZN(O1776));
  NOR2X1 G4881 (.A1(W21016), .A2(W28627), .ZN(W33148));
  NOR2X1 G4882 (.A1(I1853), .A2(W18), .ZN(W17720));
  NOR2X1 G4883 (.A1(W8035), .A2(W12665), .ZN(O1435));
  NOR2X1 G4884 (.A1(W12673), .A2(W32250), .ZN(W33149));
  NOR2X1 G4885 (.A1(W8989), .A2(W14090), .ZN(W17717));
  NOR2X1 G4886 (.A1(W27119), .A2(W16017), .ZN(W31342));
  NOR2X1 G4887 (.A1(W6350), .A2(W13017), .ZN(W17715));
  NOR2X1 G4888 (.A1(W4361), .A2(W22177), .ZN(O5762));
  NOR2X1 G4889 (.A1(W28565), .A2(W22155), .ZN(W33153));
  NOR2X1 G4890 (.A1(W14287), .A2(W10672), .ZN(W31385));
  NOR2X1 G4891 (.A1(W11536), .A2(I1925), .ZN(W19448));
  NOR2X1 G4892 (.A1(W13484), .A2(W9711), .ZN(O1434));
  NOR2X1 G4893 (.A1(W9015), .A2(W22418), .ZN(W33157));
  NOR2X1 G4894 (.A1(W2899), .A2(W7010), .ZN(W17490));
  NOR2X1 G4895 (.A1(W27663), .A2(W20528), .ZN(W31307));
  NOR2X1 G4896 (.A1(W18634), .A2(I1482), .ZN(O5731));
  NOR2X1 G4897 (.A1(W2398), .A2(W10765), .ZN(O1402));
  NOR2X1 G4898 (.A1(W33338), .A2(W22928), .ZN(W33403));
  NOR2X1 G4899 (.A1(W662), .A2(W15313), .ZN(W33405));
  NOR2X1 G4900 (.A1(W16460), .A2(W6862), .ZN(W33406));
  NOR2X1 G4901 (.A1(W3459), .A2(W5630), .ZN(W31303));
  NOR2X1 G4902 (.A1(W5709), .A2(W9760), .ZN(W19528));
  NOR2X1 G4903 (.A1(W28975), .A2(W5191), .ZN(W33397));
  NOR2X1 G4904 (.A1(W3306), .A2(I1138), .ZN(W17489));
  NOR2X1 G4905 (.A1(W9722), .A2(W20607), .ZN(O5728));
  NOR2X1 G4906 (.A1(W21483), .A2(I1204), .ZN(W33413));
  NOR2X1 G4907 (.A1(I989), .A2(W8780), .ZN(W17486));
  NOR2X1 G4908 (.A1(W2242), .A2(W1096), .ZN(W17485));
  NOR2X1 G4909 (.A1(W13686), .A2(W27382), .ZN(O6688));
  NOR2X1 G4910 (.A1(W21600), .A2(W20380), .ZN(W33419));
  NOR2X1 G4911 (.A1(W18697), .A2(W24520), .ZN(O6691));
  NOR2X1 G4912 (.A1(W16386), .A2(W13990), .ZN(W19518));
  NOR2X1 G4913 (.A1(W12101), .A2(W16258), .ZN(O1407));
  NOR2X1 G4914 (.A1(W12374), .A2(I264), .ZN(O6673));
  NOR2X1 G4915 (.A1(W16630), .A2(W3459), .ZN(W17520));
  NOR2X1 G4916 (.A1(W11896), .A2(W7834), .ZN(W17519));
  NOR2X1 G4917 (.A1(W10829), .A2(W29098), .ZN(O6674));
  NOR2X1 G4918 (.A1(W32972), .A2(W29846), .ZN(W33371));
  NOR2X1 G4919 (.A1(W11412), .A2(W5068), .ZN(O1406));
  NOR2X1 G4920 (.A1(W9819), .A2(W15809), .ZN(O6675));
  NOR2X1 G4921 (.A1(W7766), .A2(W24679), .ZN(W31300));
  NOR2X1 G4922 (.A1(W18133), .A2(W27921), .ZN(W33377));
  NOR2X1 G4923 (.A1(I1144), .A2(W23638), .ZN(O6676));
  NOR2X1 G4924 (.A1(W29241), .A2(W6817), .ZN(W31314));
  NOR2X1 G4925 (.A1(W23201), .A2(I1724), .ZN(O6678));
  NOR2X1 G4926 (.A1(W6144), .A2(W13009), .ZN(O1404));
  NOR2X1 G4927 (.A1(W6329), .A2(W1416), .ZN(W33384));
  NOR2X1 G4928 (.A1(W26192), .A2(W25878), .ZN(W33387));
  NOR2X1 G4929 (.A1(W12816), .A2(W6554), .ZN(W17453));
  NOR2X1 G4930 (.A1(W19563), .A2(W7674), .ZN(W33444));
  NOR2X1 G4931 (.A1(W4421), .A2(I1769), .ZN(W31293));
  NOR2X1 G4932 (.A1(W9156), .A2(W2934), .ZN(W17459));
  NOR2X1 G4933 (.A1(W12168), .A2(W675), .ZN(W19538));
  NOR2X1 G4934 (.A1(W13460), .A2(W16975), .ZN(O5723));
  NOR2X1 G4935 (.A1(W10862), .A2(W22769), .ZN(O6704));
  NOR2X1 G4936 (.A1(W15734), .A2(W11937), .ZN(W17455));
  NOR2X1 G4937 (.A1(W13392), .A2(W11304), .ZN(O6706));
  NOR2X1 G4938 (.A1(W13098), .A2(W4802), .ZN(O6702));
  NOR2X1 G4939 (.A1(W11845), .A2(W1161), .ZN(W17452));
  NOR2X1 G4940 (.A1(W4931), .A2(W30343), .ZN(O6708));
  NOR2X1 G4941 (.A1(W29303), .A2(W8793), .ZN(W33455));
  NOR2X1 G4942 (.A1(W28544), .A2(W32454), .ZN(O6709));
  NOR2X1 G4943 (.A1(W23498), .A2(W26990), .ZN(W31288));
  NOR2X1 G4944 (.A1(W955), .A2(W6989), .ZN(W17446));
  NOR2X1 G4945 (.A1(W11499), .A2(W28835), .ZN(O6711));
  NOR2X1 G4946 (.A1(W8413), .A2(W159), .ZN(W19542));
  NOR2X1 G4947 (.A1(W472), .A2(W10392), .ZN(W17471));
  NOR2X1 G4948 (.A1(W13362), .A2(I1586), .ZN(O1400));
  NOR2X1 G4949 (.A1(W3166), .A2(W784), .ZN(W19532));
  NOR2X1 G4950 (.A1(W2346), .A2(W16808), .ZN(W19533));
  NOR2X1 G4951 (.A1(W15562), .A2(W4147), .ZN(W17476));
  NOR2X1 G4952 (.A1(W21301), .A2(W9606), .ZN(O6695));
  NOR2X1 G4953 (.A1(W11854), .A2(W11304), .ZN(O1397));
  NOR2X1 G4954 (.A1(W18441), .A2(W23534), .ZN(W33429));
  NOR2X1 G4955 (.A1(W15802), .A2(W8827), .ZN(O1396));
  NOR2X1 G4956 (.A1(W15659), .A2(W32823), .ZN(W33367));
  NOR2X1 G4957 (.A1(W8901), .A2(W6876), .ZN(W17470));
  NOR2X1 G4958 (.A1(W8831), .A2(W24142), .ZN(O6697));
  NOR2X1 G4959 (.A1(W32430), .A2(I250), .ZN(W33435));
  NOR2X1 G4960 (.A1(W13781), .A2(W4428), .ZN(W19534));
  NOR2X1 G4961 (.A1(W6377), .A2(W27823), .ZN(W33437));
  NOR2X1 G4962 (.A1(W4786), .A2(W30719), .ZN(W33439));
  NOR2X1 G4963 (.A1(W2367), .A2(W10744), .ZN(O5724));
  NOR2X1 G4964 (.A1(W15353), .A2(W3372), .ZN(W19498));
  NOR2X1 G4965 (.A1(W9243), .A2(W12884), .ZN(W17582));
  NOR2X1 G4966 (.A1(W6266), .A2(W12131), .ZN(W17581));
  NOR2X1 G4967 (.A1(W1692), .A2(W2586), .ZN(W31335));
  NOR2X1 G4968 (.A1(W32871), .A2(W19156), .ZN(W33306));
  NOR2X1 G4969 (.A1(W31888), .A2(W22879), .ZN(W33307));
  NOR2X1 G4970 (.A1(W3449), .A2(I1267), .ZN(W17577));
  NOR2X1 G4971 (.A1(W16847), .A2(W6682), .ZN(W19497));
  NOR2X1 G4972 (.A1(W28136), .A2(W20345), .ZN(W33309));
  NOR2X1 G4973 (.A1(W15662), .A2(W17221), .ZN(O6639));
  NOR2X1 G4974 (.A1(W858), .A2(W11347), .ZN(W17573));
  NOR2X1 G4975 (.A1(W9405), .A2(W16463), .ZN(W19499));
  NOR2X1 G4976 (.A1(W8308), .A2(W3016), .ZN(W31334));
  NOR2X1 G4977 (.A1(W17260), .A2(W12716), .ZN(W17570));
  NOR2X1 G4978 (.A1(W12995), .A2(W3355), .ZN(O1411));
  NOR2X1 G4979 (.A1(W33053), .A2(I1195), .ZN(W33316));
  NOR2X1 G4980 (.A1(W16941), .A2(W8303), .ZN(W17565));
  NOR2X1 G4981 (.A1(W1456), .A2(W7702), .ZN(W17564));
  NOR2X1 G4982 (.A1(W16964), .A2(W6862), .ZN(W33295));
  NOR2X1 G4983 (.A1(W31708), .A2(W1863), .ZN(W33287));
  NOR2X1 G4984 (.A1(W1346), .A2(I1314), .ZN(W19490));
  NOR2X1 G4985 (.A1(W6547), .A2(W15380), .ZN(W33289));
  NOR2X1 G4986 (.A1(I1273), .A2(W32292), .ZN(W33290));
  NOR2X1 G4987 (.A1(W14225), .A2(W4218), .ZN(W17596));
  NOR2X1 G4988 (.A1(W13754), .A2(W28015), .ZN(O5744));
  NOR2X1 G4989 (.A1(W7602), .A2(W31417), .ZN(W33292));
  NOR2X1 G4990 (.A1(W15774), .A2(W13693), .ZN(W17593));
  NOR2X1 G4991 (.A1(W18465), .A2(W13501), .ZN(W33325));
  NOR2X1 G4992 (.A1(W9530), .A2(W10653), .ZN(W33296));
  NOR2X1 G4993 (.A1(W15395), .A2(W14597), .ZN(W17590));
  NOR2X1 G4994 (.A1(I1847), .A2(W20343), .ZN(O6637));
  NOR2X1 G4995 (.A1(W6329), .A2(W11026), .ZN(O1784));
  NOR2X1 G4996 (.A1(W10499), .A2(W14785), .ZN(O5742));
  NOR2X1 G4997 (.A1(W11019), .A2(W1941), .ZN(W17585));
  NOR2X1 G4998 (.A1(W8158), .A2(W4623), .ZN(O1785));
  NOR2X1 G4999 (.A1(W28016), .A2(W23875), .ZN(W33355));
  NOR2X1 G5000 (.A1(W15896), .A2(W18624), .ZN(W19509));
  NOR2X1 G5001 (.A1(W11923), .A2(W2644), .ZN(W17540));
  NOR2X1 G5002 (.A1(W13617), .A2(W18021), .ZN(W33346));
  NOR2X1 G5003 (.A1(W8080), .A2(W9917), .ZN(W33347));
  NOR2X1 G5004 (.A1(W18715), .A2(W12577), .ZN(O1787));
  NOR2X1 G5005 (.A1(W30804), .A2(W1842), .ZN(W31322));
  NOR2X1 G5006 (.A1(W13697), .A2(W6200), .ZN(O5734));
  NOR2X1 G5007 (.A1(I308), .A2(W20863), .ZN(W33354));
  NOR2X1 G5008 (.A1(W4338), .A2(W8455), .ZN(W17542));
  NOR2X1 G5009 (.A1(W24206), .A2(W25428), .ZN(O6667));
  NOR2X1 G5010 (.A1(W5870), .A2(W549), .ZN(W17530));
  NOR2X1 G5011 (.A1(W32779), .A2(W9809), .ZN(O6668));
  NOR2X1 G5012 (.A1(W2109), .A2(W4499), .ZN(W17528));
  NOR2X1 G5013 (.A1(W10850), .A2(W28983), .ZN(O6670));
  NOR2X1 G5014 (.A1(W26897), .A2(I458), .ZN(O6671));
  NOR2X1 G5015 (.A1(W17991), .A2(W27132), .ZN(O5733));
  NOR2X1 G5016 (.A1(W3784), .A2(W17838), .ZN(W19515));
  NOR2X1 G5017 (.A1(W15352), .A2(W4563), .ZN(W17552));
  NOR2X1 G5018 (.A1(I606), .A2(W6201), .ZN(W17560));
  NOR2X1 G5019 (.A1(W24507), .A2(W21655), .ZN(W33327));
  NOR2X1 G5020 (.A1(W4879), .A2(W12855), .ZN(W17558));
  NOR2X1 G5021 (.A1(W1414), .A2(W21903), .ZN(W31327));
  NOR2X1 G5022 (.A1(W26307), .A2(W26562), .ZN(O6652));
  NOR2X1 G5023 (.A1(W4426), .A2(W26410), .ZN(W33332));
  NOR2X1 G5024 (.A1(W8194), .A2(W21918), .ZN(W33333));
  NOR2X1 G5025 (.A1(W7403), .A2(I622), .ZN(W19506));
  NOR2X1 G5026 (.A1(I1800), .A2(W448), .ZN(O1328));
  NOR2X1 G5027 (.A1(W23728), .A2(W25418), .ZN(O6655));
  NOR2X1 G5028 (.A1(W15747), .A2(W14108), .ZN(W17549));
  NOR2X1 G5029 (.A1(W1093), .A2(W12453), .ZN(W17548));
  NOR2X1 G5030 (.A1(W10328), .A2(W16837), .ZN(W17547));
  NOR2X1 G5031 (.A1(W11143), .A2(W12680), .ZN(W17546));
  NOR2X1 G5032 (.A1(W12856), .A2(W29355), .ZN(O6658));
  NOR2X1 G5033 (.A1(W18149), .A2(W26509), .ZN(O6661));
  NOR2X1 G5034 (.A1(W11767), .A2(W2298), .ZN(W16708));
  NOR2X1 G5035 (.A1(W3267), .A2(W23226), .ZN(O7107));
  NOR2X1 G5036 (.A1(I1165), .A2(W15615), .ZN(W34177));
  NOR2X1 G5037 (.A1(W28484), .A2(W11596), .ZN(O7111));
  NOR2X1 G5038 (.A1(W16612), .A2(W4816), .ZN(O1236));
  NOR2X1 G5039 (.A1(W5887), .A2(W30127), .ZN(O7112));
  NOR2X1 G5040 (.A1(W1124), .A2(W946), .ZN(O1235));
  NOR2X1 G5041 (.A1(W24906), .A2(W28623), .ZN(O5612));
  NOR2X1 G5042 (.A1(W10075), .A2(W15130), .ZN(W16709));
  NOR2X1 G5043 (.A1(W15312), .A2(W7081), .ZN(O7106));
  NOR2X1 G5044 (.A1(W24028), .A2(W21788), .ZN(O7114));
  NOR2X1 G5045 (.A1(W11854), .A2(W13927), .ZN(W34187));
  NOR2X1 G5046 (.A1(W19722), .A2(W7251), .ZN(W34190));
  NOR2X1 G5047 (.A1(W3777), .A2(W22667), .ZN(W34191));
  NOR2X1 G5048 (.A1(W5974), .A2(W13171), .ZN(W16702));
  NOR2X1 G5049 (.A1(W5399), .A2(W15321), .ZN(W16701));
  NOR2X1 G5050 (.A1(W7322), .A2(W7775), .ZN(W34192));
  NOR2X1 G5051 (.A1(W31058), .A2(W22213), .ZN(O7116));
  NOR2X1 G5052 (.A1(I410), .A2(W8212), .ZN(O1241));
  NOR2X1 G5053 (.A1(W4904), .A2(W12544), .ZN(W16739));
  NOR2X1 G5054 (.A1(W14443), .A2(W11049), .ZN(O5621));
  NOR2X1 G5055 (.A1(I936), .A2(W8750), .ZN(O7096));
  NOR2X1 G5056 (.A1(W14862), .A2(W18005), .ZN(O7098));
  NOR2X1 G5057 (.A1(W3018), .A2(W5637), .ZN(O7099));
  NOR2X1 G5058 (.A1(W1636), .A2(W4551), .ZN(W19793));
  NOR2X1 G5059 (.A1(W8028), .A2(I1509), .ZN(O5619));
  NOR2X1 G5060 (.A1(W5955), .A2(W15834), .ZN(W34166));
  NOR2X1 G5061 (.A1(W7491), .A2(W26346), .ZN(O5607));
  NOR2X1 G5062 (.A1(W9382), .A2(W11153), .ZN(W16729));
  NOR2X1 G5063 (.A1(W8538), .A2(I1948), .ZN(O1240));
  NOR2X1 G5064 (.A1(W12823), .A2(W8571), .ZN(O1855));
  NOR2X1 G5065 (.A1(W11753), .A2(W5135), .ZN(O5618));
  NOR2X1 G5066 (.A1(W15556), .A2(W19742), .ZN(O5615));
  NOR2X1 G5067 (.A1(W10016), .A2(W7898), .ZN(W16722));
  NOR2X1 G5068 (.A1(W8065), .A2(W6571), .ZN(O1239));
  NOR2X1 G5069 (.A1(W12262), .A2(W5720), .ZN(W16666));
  NOR2X1 G5070 (.A1(W10578), .A2(W15176), .ZN(O1861));
  NOR2X1 G5071 (.A1(I1519), .A2(W11796), .ZN(O1225));
  NOR2X1 G5072 (.A1(W6164), .A2(W6253), .ZN(O1862));
  NOR2X1 G5073 (.A1(I1263), .A2(W13511), .ZN(W19817));
  NOR2X1 G5074 (.A1(W3638), .A2(W9477), .ZN(W16671));
  NOR2X1 G5075 (.A1(W11058), .A2(W15083), .ZN(W16670));
  NOR2X1 G5076 (.A1(W1698), .A2(W3665), .ZN(W16668));
  NOR2X1 G5077 (.A1(W24779), .A2(W22687), .ZN(O7137));
  NOR2X1 G5078 (.A1(W17581), .A2(W719), .ZN(W19813));
  NOR2X1 G5079 (.A1(W15060), .A2(W13493), .ZN(W16665));
  NOR2X1 G5080 (.A1(W32552), .A2(W3076), .ZN(O7138));
  NOR2X1 G5081 (.A1(W1027), .A2(W18081), .ZN(W19819));
  NOR2X1 G5082 (.A1(W16783), .A2(W17284), .ZN(W19820));
  NOR2X1 G5083 (.A1(W7041), .A2(W2093), .ZN(W16661));
  NOR2X1 G5084 (.A1(W253), .A2(W12749), .ZN(O1223));
  NOR2X1 G5085 (.A1(W4183), .A2(W1280), .ZN(W34232));
  NOR2X1 G5086 (.A1(I987), .A2(W12178), .ZN(W16658));
  NOR2X1 G5087 (.A1(W27535), .A2(W28709), .ZN(O7126));
  NOR2X1 G5088 (.A1(I286), .A2(W15650), .ZN(W16695));
  NOR2X1 G5089 (.A1(W641), .A2(W1575), .ZN(O1231));
  NOR2X1 G5090 (.A1(W30426), .A2(W6719), .ZN(O7122));
  NOR2X1 G5091 (.A1(W566), .A2(W9700), .ZN(O1229));
  NOR2X1 G5092 (.A1(W12720), .A2(W16318), .ZN(W34206));
  NOR2X1 G5093 (.A1(W29636), .A2(W12148), .ZN(O5604));
  NOR2X1 G5094 (.A1(W6729), .A2(W6823), .ZN(W16687));
  NOR2X1 G5095 (.A1(W17862), .A2(I90), .ZN(O5603));
  NOR2X1 G5096 (.A1(W10084), .A2(W18536), .ZN(O7091));
  NOR2X1 G5097 (.A1(W14967), .A2(W26792), .ZN(O7127));
  NOR2X1 G5098 (.A1(W24066), .A2(W7285), .ZN(W31010));
  NOR2X1 G5099 (.A1(W15831), .A2(W11867), .ZN(W16682));
  NOR2X1 G5100 (.A1(W10799), .A2(W13092), .ZN(W16681));
  NOR2X1 G5101 (.A1(W18492), .A2(W9026), .ZN(W34217));
  NOR2X1 G5102 (.A1(W28040), .A2(W10551), .ZN(O7130));
  NOR2X1 G5103 (.A1(W6866), .A2(W2033), .ZN(W16678));
  NOR2X1 G5104 (.A1(W9527), .A2(W8029), .ZN(W16787));
  NOR2X1 G5105 (.A1(W3799), .A2(W8455), .ZN(O1264));
  NOR2X1 G5106 (.A1(W2814), .A2(W10371), .ZN(W19775));
  NOR2X1 G5107 (.A1(W3527), .A2(W11488), .ZN(W19776));
  NOR2X1 G5108 (.A1(W7157), .A2(W4139), .ZN(W19777));
  NOR2X1 G5109 (.A1(W13101), .A2(W17453), .ZN(W19779));
  NOR2X1 G5110 (.A1(I562), .A2(W16164), .ZN(W16790));
  NOR2X1 G5111 (.A1(W12756), .A2(W8781), .ZN(W34109));
  NOR2X1 G5112 (.A1(I904), .A2(W3891), .ZN(W16788));
  NOR2X1 G5113 (.A1(W19520), .A2(W21769), .ZN(O7065));
  NOR2X1 G5114 (.A1(W12271), .A2(W11120), .ZN(O1260));
  NOR2X1 G5115 (.A1(W32095), .A2(W19229), .ZN(O7071));
  NOR2X1 G5116 (.A1(W7854), .A2(W2724), .ZN(W16784));
  NOR2X1 G5117 (.A1(W10869), .A2(W190), .ZN(W34111));
  NOR2X1 G5118 (.A1(W6591), .A2(W525), .ZN(W16782));
  NOR2X1 G5119 (.A1(W26577), .A2(W8610), .ZN(O7072));
  NOR2X1 G5120 (.A1(W30995), .A2(W24937), .ZN(W34114));
  NOR2X1 G5121 (.A1(W2425), .A2(W7252), .ZN(W16779));
  NOR2X1 G5122 (.A1(W9524), .A2(W14748), .ZN(O5629));
  NOR2X1 G5123 (.A1(W26721), .A2(W33124), .ZN(W34082));
  NOR2X1 G5124 (.A1(W4808), .A2(W23178), .ZN(W31067));
  NOR2X1 G5125 (.A1(W3422), .A2(W9582), .ZN(W34084));
  NOR2X1 G5126 (.A1(W30361), .A2(W1367), .ZN(O7059));
  NOR2X1 G5127 (.A1(W15971), .A2(W13831), .ZN(O1848));
  NOR2X1 G5128 (.A1(I1675), .A2(W8985), .ZN(W16809));
  NOR2X1 G5129 (.A1(W3353), .A2(W14991), .ZN(W19769));
  NOR2X1 G5130 (.A1(W18150), .A2(I54), .ZN(W31066));
  NOR2X1 G5131 (.A1(W15783), .A2(I1990), .ZN(W31059));
  NOR2X1 G5132 (.A1(W15819), .A2(W4078), .ZN(W16805));
  NOR2X1 G5133 (.A1(W7704), .A2(W27140), .ZN(W31064));
  NOR2X1 G5134 (.A1(W2210), .A2(W1189), .ZN(W16803));
  NOR2X1 G5135 (.A1(W11748), .A2(W21595), .ZN(W31062));
  NOR2X1 G5136 (.A1(W3697), .A2(W18778), .ZN(W19774));
  NOR2X1 G5137 (.A1(W28408), .A2(W33026), .ZN(W34097));
  NOR2X1 G5138 (.A1(W11261), .A2(W9885), .ZN(O1265));
  NOR2X1 G5139 (.A1(W8639), .A2(W8172), .ZN(O1853));
  NOR2X1 G5140 (.A1(I501), .A2(W22314), .ZN(W34133));
  NOR2X1 G5141 (.A1(W12779), .A2(W16116), .ZN(W16758));
  NOR2X1 G5142 (.A1(W6284), .A2(W3563), .ZN(W16757));
  NOR2X1 G5143 (.A1(W8518), .A2(W5155), .ZN(W16756));
  NOR2X1 G5144 (.A1(W13061), .A2(W14837), .ZN(W16754));
  NOR2X1 G5145 (.A1(W3078), .A2(W25066), .ZN(W34135));
  NOR2X1 G5146 (.A1(W4821), .A2(W10766), .ZN(O1252));
  NOR2X1 G5147 (.A1(W3702), .A2(W29779), .ZN(O5625));
  NOR2X1 G5148 (.A1(W15154), .A2(W6983), .ZN(W16760));
  NOR2X1 G5149 (.A1(W11295), .A2(W8828), .ZN(W16749));
  NOR2X1 G5150 (.A1(W22062), .A2(W22531), .ZN(W31049));
  NOR2X1 G5151 (.A1(W18778), .A2(W1445), .ZN(W34142));
  NOR2X1 G5152 (.A1(W31898), .A2(W3381), .ZN(W34143));
  NOR2X1 G5153 (.A1(W14599), .A2(W11938), .ZN(W16745));
  NOR2X1 G5154 (.A1(I1160), .A2(I1547), .ZN(W16743));
  NOR2X1 G5155 (.A1(W2571), .A2(W5921), .ZN(O1246));
  NOR2X1 G5156 (.A1(W11486), .A2(W23576), .ZN(O7089));
  NOR2X1 G5157 (.A1(W13393), .A2(I1002), .ZN(O1256));
  NOR2X1 G5158 (.A1(W7868), .A2(W2627), .ZN(W34117));
  NOR2X1 G5159 (.A1(W31906), .A2(W14024), .ZN(O7075));
  NOR2X1 G5160 (.A1(I233), .A2(W16851), .ZN(O7076));
  NOR2X1 G5161 (.A1(W23123), .A2(W29163), .ZN(W31057));
  NOR2X1 G5162 (.A1(W13705), .A2(W2228), .ZN(W16773));
  NOR2X1 G5163 (.A1(W29947), .A2(W19145), .ZN(O7077));
  NOR2X1 G5164 (.A1(W23136), .A2(W23688), .ZN(O7078));
  NOR2X1 G5165 (.A1(W33686), .A2(W20413), .ZN(O7080));
  NOR2X1 G5166 (.A1(W7230), .A2(W15992), .ZN(W16657));
  NOR2X1 G5167 (.A1(W16290), .A2(W1984), .ZN(W16768));
  NOR2X1 G5168 (.A1(W4084), .A2(W7839), .ZN(W16767));
  NOR2X1 G5169 (.A1(W29867), .A2(W29141), .ZN(O7081));
  NOR2X1 G5170 (.A1(W14599), .A2(W16717), .ZN(W34127));
  NOR2X1 G5171 (.A1(W16262), .A2(W14472), .ZN(W19783));
  NOR2X1 G5172 (.A1(W10967), .A2(I1165), .ZN(W16762));
  NOR2X1 G5173 (.A1(W10649), .A2(W11394), .ZN(O5626));
  NOR2X1 G5174 (.A1(W6938), .A2(W16111), .ZN(W16544));
  NOR2X1 G5175 (.A1(W5133), .A2(W12355), .ZN(W16553));
  NOR2X1 G5176 (.A1(W15017), .A2(W30306), .ZN(W34336));
  NOR2X1 G5177 (.A1(W22857), .A2(I1377), .ZN(W34337));
  NOR2X1 G5178 (.A1(W33583), .A2(W12181), .ZN(O7201));
  NOR2X1 G5179 (.A1(W353), .A2(W6477), .ZN(O1869));
  NOR2X1 G5180 (.A1(W20898), .A2(W17828), .ZN(W34340));
  NOR2X1 G5181 (.A1(W15733), .A2(W12778), .ZN(W34342));
  NOR2X1 G5182 (.A1(W27138), .A2(W8558), .ZN(W30965));
  NOR2X1 G5183 (.A1(W1461), .A2(W15899), .ZN(W16554));
  NOR2X1 G5184 (.A1(W13012), .A2(W5322), .ZN(W16543));
  NOR2X1 G5185 (.A1(W25904), .A2(W27182), .ZN(W30963));
  NOR2X1 G5186 (.A1(I214), .A2(W13486), .ZN(O1196));
  NOR2X1 G5187 (.A1(W5412), .A2(W1029), .ZN(W34346));
  NOR2X1 G5188 (.A1(W1692), .A2(W4035), .ZN(W16539));
  NOR2X1 G5189 (.A1(W3300), .A2(W12491), .ZN(O7205));
  NOR2X1 G5190 (.A1(W8195), .A2(W5668), .ZN(W16537));
  NOR2X1 G5191 (.A1(W18596), .A2(W13303), .ZN(W34349));
  NOR2X1 G5192 (.A1(W6126), .A2(W16953), .ZN(W19857));
  NOR2X1 G5193 (.A1(I1523), .A2(W23587), .ZN(W30971));
  NOR2X1 G5194 (.A1(W15904), .A2(W9120), .ZN(W19855));
  NOR2X1 G5195 (.A1(W7282), .A2(W9250), .ZN(W16569));
  NOR2X1 G5196 (.A1(W21648), .A2(W6611), .ZN(O7195));
  NOR2X1 G5197 (.A1(W23838), .A2(W8780), .ZN(W34324));
  NOR2X1 G5198 (.A1(W20833), .A2(W1967), .ZN(W34328));
  NOR2X1 G5199 (.A1(W34136), .A2(W30663), .ZN(O7197));
  NOR2X1 G5200 (.A1(W15373), .A2(W10172), .ZN(W16563));
  NOR2X1 G5201 (.A1(W13835), .A2(W12582), .ZN(W16535));
  NOR2X1 G5202 (.A1(W488), .A2(W7274), .ZN(O5579));
  NOR2X1 G5203 (.A1(W15090), .A2(W19616), .ZN(O7199));
  NOR2X1 G5204 (.A1(W1456), .A2(W13209), .ZN(W16559));
  NOR2X1 G5205 (.A1(W29590), .A2(W7913), .ZN(O7200));
  NOR2X1 G5206 (.A1(W15775), .A2(W1277), .ZN(W16557));
  NOR2X1 G5207 (.A1(I486), .A2(W5265), .ZN(W16556));
  NOR2X1 G5208 (.A1(W22674), .A2(W10645), .ZN(W34335));
  NOR2X1 G5209 (.A1(W2946), .A2(W30461), .ZN(W34378));
  NOR2X1 G5210 (.A1(W30597), .A2(W17221), .ZN(W34367));
  NOR2X1 G5211 (.A1(W21081), .A2(I1198), .ZN(O5571));
  NOR2X1 G5212 (.A1(W14716), .A2(I661), .ZN(W16510));
  NOR2X1 G5213 (.A1(W4295), .A2(W11565), .ZN(W16509));
  NOR2X1 G5214 (.A1(I512), .A2(W363), .ZN(W16507));
  NOR2X1 G5215 (.A1(W22937), .A2(W2412), .ZN(W30953));
  NOR2X1 G5216 (.A1(W2945), .A2(W16885), .ZN(W19874));
  NOR2X1 G5217 (.A1(W17384), .A2(W14105), .ZN(O1874));
  NOR2X1 G5218 (.A1(W10700), .A2(W6120), .ZN(W16514));
  NOR2X1 G5219 (.A1(W14449), .A2(W6385), .ZN(O5568));
  NOR2X1 G5220 (.A1(W14539), .A2(W7598), .ZN(O1875));
  NOR2X1 G5221 (.A1(W31930), .A2(W3585), .ZN(O7221));
  NOR2X1 G5222 (.A1(W2847), .A2(I1758), .ZN(W16499));
  NOR2X1 G5223 (.A1(W14271), .A2(I29), .ZN(W16498));
  NOR2X1 G5224 (.A1(W12983), .A2(W9955), .ZN(W19878));
  NOR2X1 G5225 (.A1(W18174), .A2(W13204), .ZN(O5567));
  NOR2X1 G5226 (.A1(W8567), .A2(W8), .ZN(O1186));
  NOR2X1 G5227 (.A1(W8944), .A2(W4889), .ZN(W16524));
  NOR2X1 G5228 (.A1(W96), .A2(W9873), .ZN(W16533));
  NOR2X1 G5229 (.A1(W28725), .A2(W13148), .ZN(O7208));
  NOR2X1 G5230 (.A1(W3458), .A2(W7609), .ZN(W16531));
  NOR2X1 G5231 (.A1(W1460), .A2(W7884), .ZN(O7209));
  NOR2X1 G5232 (.A1(I1836), .A2(W29733), .ZN(W34354));
  NOR2X1 G5233 (.A1(I1272), .A2(W22664), .ZN(W30961));
  NOR2X1 G5234 (.A1(W2890), .A2(W23680), .ZN(W30960));
  NOR2X1 G5235 (.A1(I490), .A2(W18371), .ZN(W19866));
  NOR2X1 G5236 (.A1(W9330), .A2(W5063), .ZN(W19852));
  NOR2X1 G5237 (.A1(W11144), .A2(W7972), .ZN(O1191));
  NOR2X1 G5238 (.A1(W31981), .A2(W28750), .ZN(O7212));
  NOR2X1 G5239 (.A1(W15101), .A2(I1841), .ZN(W16521));
  NOR2X1 G5240 (.A1(W7593), .A2(W9770), .ZN(W16519));
  NOR2X1 G5241 (.A1(W4228), .A2(W17476), .ZN(W34363));
  NOR2X1 G5242 (.A1(W14889), .A2(W5046), .ZN(W16517));
  NOR2X1 G5243 (.A1(W2357), .A2(W11179), .ZN(O7213));
  NOR2X1 G5244 (.A1(W6467), .A2(W2114), .ZN(W34265));
  NOR2X1 G5245 (.A1(W9150), .A2(W16509), .ZN(W16636));
  NOR2X1 G5246 (.A1(W13971), .A2(W15325), .ZN(W16634));
  NOR2X1 G5247 (.A1(W12972), .A2(W3277), .ZN(W19830));
  NOR2X1 G5248 (.A1(W31400), .A2(W29858), .ZN(W34258));
  NOR2X1 G5249 (.A1(W15206), .A2(W6637), .ZN(W19831));
  NOR2X1 G5250 (.A1(W10666), .A2(W4919), .ZN(W16630));
  NOR2X1 G5251 (.A1(W7977), .A2(W20895), .ZN(W34262));
  NOR2X1 G5252 (.A1(W14011), .A2(W17939), .ZN(W19833));
  NOR2X1 G5253 (.A1(W18956), .A2(W7399), .ZN(W31005));
  NOR2X1 G5254 (.A1(W1612), .A2(W15744), .ZN(W16624));
  NOR2X1 G5255 (.A1(W5129), .A2(W15445), .ZN(W16623));
  NOR2X1 G5256 (.A1(W3860), .A2(W12837), .ZN(W16622));
  NOR2X1 G5257 (.A1(W15164), .A2(W3598), .ZN(O1215));
  NOR2X1 G5258 (.A1(W32962), .A2(W7596), .ZN(W34268));
  NOR2X1 G5259 (.A1(W7044), .A2(W15188), .ZN(O1214));
  NOR2X1 G5260 (.A1(W22005), .A2(W29734), .ZN(W34272));
  NOR2X1 G5261 (.A1(W8008), .A2(W12303), .ZN(W19836));
  NOR2X1 G5262 (.A1(W30119), .A2(W15274), .ZN(W34239));
  NOR2X1 G5263 (.A1(W15688), .A2(W5791), .ZN(W16655));
  NOR2X1 G5264 (.A1(W15217), .A2(W8768), .ZN(W16654));
  NOR2X1 G5265 (.A1(W25798), .A2(W23933), .ZN(W34236));
  NOR2X1 G5266 (.A1(W4540), .A2(W8354), .ZN(W16652));
  NOR2X1 G5267 (.A1(W27047), .A2(W23399), .ZN(W34237));
  NOR2X1 G5268 (.A1(W764), .A2(W17753), .ZN(O1864));
  NOR2X1 G5269 (.A1(W14337), .A2(W7627), .ZN(O1220));
  NOR2X1 G5270 (.A1(W14582), .A2(W16333), .ZN(W16648));
  NOR2X1 G5271 (.A1(W2063), .A2(W1199), .ZN(W16615));
  NOR2X1 G5272 (.A1(W12144), .A2(W5513), .ZN(W16646));
  NOR2X1 G5273 (.A1(W10185), .A2(W7704), .ZN(O1219));
  NOR2X1 G5274 (.A1(W15834), .A2(W9279), .ZN(O7148));
  NOR2X1 G5275 (.A1(W2838), .A2(W19281), .ZN(W19824));
  NOR2X1 G5276 (.A1(W7633), .A2(I1959), .ZN(W19825));
  NOR2X1 G5277 (.A1(W3664), .A2(W23043), .ZN(O7151));
  NOR2X1 G5278 (.A1(W5217), .A2(W2928), .ZN(W19826));
  NOR2X1 G5279 (.A1(W3498), .A2(W16549), .ZN(W16582));
  NOR2X1 G5280 (.A1(W4209), .A2(I504), .ZN(O1209));
  NOR2X1 G5281 (.A1(W1721), .A2(W8692), .ZN(W16593));
  NOR2X1 G5282 (.A1(W16000), .A2(I1122), .ZN(O5587));
  NOR2X1 G5283 (.A1(W10208), .A2(W8584), .ZN(W16590));
  NOR2X1 G5284 (.A1(W12843), .A2(W9353), .ZN(W16589));
  NOR2X1 G5285 (.A1(W22330), .A2(W12256), .ZN(W30978));
  NOR2X1 G5286 (.A1(W2423), .A2(W17531), .ZN(W19847));
  NOR2X1 G5287 (.A1(W5116), .A2(W11796), .ZN(W16583));
  NOR2X1 G5288 (.A1(W5839), .A2(W2963), .ZN(O7180));
  NOR2X1 G5289 (.A1(I642), .A2(W8494), .ZN(W16581));
  NOR2X1 G5290 (.A1(I567), .A2(W58), .ZN(O1207));
  NOR2X1 G5291 (.A1(W27991), .A2(W22155), .ZN(W34311));
  NOR2X1 G5292 (.A1(W13584), .A2(W14893), .ZN(O7188));
  NOR2X1 G5293 (.A1(I1200), .A2(W23960), .ZN(O7189));
  NOR2X1 G5294 (.A1(W34111), .A2(W31176), .ZN(O7191));
  NOR2X1 G5295 (.A1(W17441), .A2(W30922), .ZN(W30973));
  NOR2X1 G5296 (.A1(W3434), .A2(W6692), .ZN(O1206));
  NOR2X1 G5297 (.A1(W17353), .A2(W18303), .ZN(O7165));
  NOR2X1 G5298 (.A1(W11101), .A2(W2462), .ZN(W16614));
  NOR2X1 G5299 (.A1(W19322), .A2(W3523), .ZN(W30995));
  NOR2X1 G5300 (.A1(W10541), .A2(W2477), .ZN(W34275));
  NOR2X1 G5301 (.A1(W9299), .A2(W18134), .ZN(W19838));
  NOR2X1 G5302 (.A1(W11129), .A2(W14546), .ZN(O7162));
  NOR2X1 G5303 (.A1(W20160), .A2(W10761), .ZN(O7163));
  NOR2X1 G5304 (.A1(W12337), .A2(W2753), .ZN(O1213));
  NOR2X1 G5305 (.A1(W10775), .A2(W10926), .ZN(W16607));
  NOR2X1 G5306 (.A1(W9369), .A2(W3975), .ZN(W16816));
  NOR2X1 G5307 (.A1(W18316), .A2(W18777), .ZN(W19839));
  NOR2X1 G5308 (.A1(W12680), .A2(W16914), .ZN(O5593));
  NOR2X1 G5309 (.A1(I1909), .A2(W5333), .ZN(W16602));
  NOR2X1 G5310 (.A1(W18008), .A2(W21824), .ZN(O7174));
  NOR2X1 G5311 (.A1(W23702), .A2(W26146), .ZN(O7175));
  NOR2X1 G5312 (.A1(W10085), .A2(W684), .ZN(O1211));
  NOR2X1 G5313 (.A1(W17551), .A2(W6061), .ZN(O7176));
  NOR2X1 G5314 (.A1(W7328), .A2(W11743), .ZN(O6938));
  NOR2X1 G5315 (.A1(W28355), .A2(W33), .ZN(O5658));
  NOR2X1 G5316 (.A1(W2384), .A2(W6411), .ZN(W17027));
  NOR2X1 G5317 (.A1(W12116), .A2(W18957), .ZN(W33888));
  NOR2X1 G5318 (.A1(W8505), .A2(W2283), .ZN(W17025));
  NOR2X1 G5319 (.A1(W5981), .A2(W7132), .ZN(W17024));
  NOR2X1 G5320 (.A1(W16466), .A2(I1021), .ZN(W17023));
  NOR2X1 G5321 (.A1(W14147), .A2(W1375), .ZN(O6937));
  NOR2X1 G5322 (.A1(W31683), .A2(W28842), .ZN(W33890));
  NOR2X1 G5323 (.A1(W19447), .A2(W22235), .ZN(O6935));
  NOR2X1 G5324 (.A1(W25202), .A2(W21262), .ZN(W33893));
  NOR2X1 G5325 (.A1(W1320), .A2(W14340), .ZN(W17017));
  NOR2X1 G5326 (.A1(W18130), .A2(W10774), .ZN(W19697));
  NOR2X1 G5327 (.A1(W5278), .A2(W2035), .ZN(W33900));
  NOR2X1 G5328 (.A1(W2504), .A2(W32533), .ZN(O6945));
  NOR2X1 G5329 (.A1(W19408), .A2(W12939), .ZN(W33902));
  NOR2X1 G5330 (.A1(W13581), .A2(W6143), .ZN(W17010));
  NOR2X1 G5331 (.A1(W16377), .A2(W7501), .ZN(W19699));
  NOR2X1 G5332 (.A1(W22245), .A2(W26633), .ZN(O6929));
  NOR2X1 G5333 (.A1(W16738), .A2(W17803), .ZN(O1822));
  NOR2X1 G5334 (.A1(W32784), .A2(W23228), .ZN(W33869));
  NOR2X1 G5335 (.A1(W14218), .A2(W15364), .ZN(W17043));
  NOR2X1 G5336 (.A1(W6146), .A2(W8620), .ZN(W19686));
  NOR2X1 G5337 (.A1(W15982), .A2(W18108), .ZN(O5663));
  NOR2X1 G5338 (.A1(W14322), .A2(W11018), .ZN(W17040));
  NOR2X1 G5339 (.A1(I1509), .A2(W549), .ZN(W17039));
  NOR2X1 G5340 (.A1(W8510), .A2(W11731), .ZN(W19688));
  NOR2X1 G5341 (.A1(W4949), .A2(W3922), .ZN(O6946));
  NOR2X1 G5342 (.A1(W9167), .A2(W1236), .ZN(O5662));
  NOR2X1 G5343 (.A1(W1287), .A2(W490), .ZN(W17035));
  NOR2X1 G5344 (.A1(W8177), .A2(W7511), .ZN(W19690));
  NOR2X1 G5345 (.A1(W10761), .A2(W15643), .ZN(W33880));
  NOR2X1 G5346 (.A1(W2083), .A2(W10958), .ZN(W19691));
  NOR2X1 G5347 (.A1(W13712), .A2(W1413), .ZN(W31146));
  NOR2X1 G5348 (.A1(W13405), .A2(W22629), .ZN(O5660));
  NOR2X1 G5349 (.A1(W2780), .A2(W5881), .ZN(W16980));
  NOR2X1 G5350 (.A1(W6706), .A2(W6689), .ZN(O1295));
  NOR2X1 G5351 (.A1(W13936), .A2(W5908), .ZN(W19706));
  NOR2X1 G5352 (.A1(W21314), .A2(W4554), .ZN(O6960));
  NOR2X1 G5353 (.A1(W5226), .A2(W10303), .ZN(O1293));
  NOR2X1 G5354 (.A1(W10503), .A2(W7737), .ZN(W16984));
  NOR2X1 G5355 (.A1(W14868), .A2(W14780), .ZN(W16983));
  NOR2X1 G5356 (.A1(W10716), .A2(W6961), .ZN(W16982));
  NOR2X1 G5357 (.A1(W1448), .A2(W14279), .ZN(O6962));
  NOR2X1 G5358 (.A1(W16273), .A2(W15933), .ZN(W16990));
  NOR2X1 G5359 (.A1(W13695), .A2(W7210), .ZN(O6963));
  NOR2X1 G5360 (.A1(I919), .A2(W16807), .ZN(O1291));
  NOR2X1 G5361 (.A1(W13099), .A2(W5556), .ZN(W16977));
  NOR2X1 G5362 (.A1(I1784), .A2(W16158), .ZN(W16976));
  NOR2X1 G5363 (.A1(W10819), .A2(I21), .ZN(W16975));
  NOR2X1 G5364 (.A1(W3643), .A2(W22082), .ZN(O5650));
  NOR2X1 G5365 (.A1(W12744), .A2(I428), .ZN(W16973));
  NOR2X1 G5366 (.A1(W11872), .A2(W4155), .ZN(W16972));
  NOR2X1 G5367 (.A1(W379), .A2(W2514), .ZN(W16998));
  NOR2X1 G5368 (.A1(I140), .A2(W23064), .ZN(W31139));
  NOR2X1 G5369 (.A1(W14782), .A2(I1542), .ZN(O5655));
  NOR2X1 G5370 (.A1(W32893), .A2(W7066), .ZN(W33908));
  NOR2X1 G5371 (.A1(W25230), .A2(W16312), .ZN(O6949));
  NOR2X1 G5372 (.A1(I44), .A2(W8492), .ZN(W19702));
  NOR2X1 G5373 (.A1(W3342), .A2(W10049), .ZN(W17001));
  NOR2X1 G5374 (.A1(W28957), .A2(W9281), .ZN(O6953));
  NOR2X1 G5375 (.A1(W6953), .A2(W409), .ZN(W16999));
  NOR2X1 G5376 (.A1(W17999), .A2(W16787), .ZN(W19684));
  NOR2X1 G5377 (.A1(W1316), .A2(W16528), .ZN(W16997));
  NOR2X1 G5378 (.A1(W6369), .A2(W14784), .ZN(W31130));
  NOR2X1 G5379 (.A1(W26038), .A2(W25554), .ZN(O6954));
  NOR2X1 G5380 (.A1(W22106), .A2(W4551), .ZN(O6955));
  NOR2X1 G5381 (.A1(I1872), .A2(W1449), .ZN(W19705));
  NOR2X1 G5382 (.A1(W8303), .A2(W6588), .ZN(W16992));
  NOR2X1 G5383 (.A1(W29039), .A2(W3338), .ZN(O6958));
  NOR2X1 G5384 (.A1(W13070), .A2(W3206), .ZN(W17098));
  NOR2X1 G5385 (.A1(W3097), .A2(W5829), .ZN(W19662));
  NOR2X1 G5386 (.A1(W12644), .A2(W7790), .ZN(W17108));
  NOR2X1 G5387 (.A1(W17341), .A2(W10336), .ZN(W19663));
  NOR2X1 G5388 (.A1(W12822), .A2(W14867), .ZN(O6889));
  NOR2X1 G5389 (.A1(W10975), .A2(W12826), .ZN(O1318));
  NOR2X1 G5390 (.A1(W1734), .A2(W8645), .ZN(W17103));
  NOR2X1 G5391 (.A1(W10246), .A2(W1315), .ZN(O6891));
  NOR2X1 G5392 (.A1(W21709), .A2(W22511), .ZN(O6892));
  NOR2X1 G5393 (.A1(W10633), .A2(W1895), .ZN(W19660));
  NOR2X1 G5394 (.A1(W13734), .A2(I1436), .ZN(W17096));
  NOR2X1 G5395 (.A1(W14047), .A2(W24326), .ZN(W33810));
  NOR2X1 G5396 (.A1(W8913), .A2(W1217), .ZN(O1818));
  NOR2X1 G5397 (.A1(W16768), .A2(W13490), .ZN(O6897));
  NOR2X1 G5398 (.A1(I596), .A2(I276), .ZN(O6898));
  NOR2X1 G5399 (.A1(W13674), .A2(W4845), .ZN(O1819));
  NOR2X1 G5400 (.A1(W23528), .A2(W17871), .ZN(O5671));
  NOR2X1 G5401 (.A1(W1039), .A2(W13986), .ZN(O1820));
  NOR2X1 G5402 (.A1(W27578), .A2(W16977), .ZN(O6877));
  NOR2X1 G5403 (.A1(W13273), .A2(W32182), .ZN(W33775));
  NOR2X1 G5404 (.A1(W16584), .A2(W4819), .ZN(W17128));
  NOR2X1 G5405 (.A1(W13487), .A2(W14495), .ZN(O6874));
  NOR2X1 G5406 (.A1(W17039), .A2(W7687), .ZN(W17126));
  NOR2X1 G5407 (.A1(W3244), .A2(I809), .ZN(O6875));
  NOR2X1 G5408 (.A1(W4904), .A2(W11749), .ZN(O1325));
  NOR2X1 G5409 (.A1(W17995), .A2(W20062), .ZN(W31181));
  NOR2X1 G5410 (.A1(W347), .A2(W1214), .ZN(W33780));
  NOR2X1 G5411 (.A1(W12973), .A2(W4372), .ZN(O1315));
  NOR2X1 G5412 (.A1(W2405), .A2(W4990), .ZN(W33785));
  NOR2X1 G5413 (.A1(I1440), .A2(W3670), .ZN(O6879));
  NOR2X1 G5414 (.A1(W31392), .A2(W26302), .ZN(W33787));
  NOR2X1 G5415 (.A1(I1143), .A2(W12466), .ZN(W33788));
  NOR2X1 G5416 (.A1(I1267), .A2(W31059), .ZN(W33790));
  NOR2X1 G5417 (.A1(W6926), .A2(W17017), .ZN(W17114));
  NOR2X1 G5418 (.A1(W210), .A2(W14871), .ZN(O6881));
  NOR2X1 G5419 (.A1(W16196), .A2(W12360), .ZN(O1306));
  NOR2X1 G5420 (.A1(W2031), .A2(W15554), .ZN(W31160));
  NOR2X1 G5421 (.A1(W5373), .A2(W1879), .ZN(W17066));
  NOR2X1 G5422 (.A1(W30937), .A2(W1016), .ZN(W33846));
  NOR2X1 G5423 (.A1(W877), .A2(W10209), .ZN(W17063));
  NOR2X1 G5424 (.A1(W21593), .A2(I1650), .ZN(W33848));
  NOR2X1 G5425 (.A1(W33254), .A2(W223), .ZN(O6917));
  NOR2X1 G5426 (.A1(W16058), .A2(W14763), .ZN(W17060));
  NOR2X1 G5427 (.A1(I1722), .A2(W17048), .ZN(O6920));
  NOR2X1 G5428 (.A1(W8247), .A2(W7356), .ZN(W17068));
  NOR2X1 G5429 (.A1(W25557), .A2(W9038), .ZN(O6921));
  NOR2X1 G5430 (.A1(I244), .A2(W9857), .ZN(O5666));
  NOR2X1 G5431 (.A1(W11594), .A2(W31884), .ZN(W33856));
  NOR2X1 G5432 (.A1(W8563), .A2(I1302), .ZN(W33857));
  NOR2X1 G5433 (.A1(W145), .A2(W6225), .ZN(W17052));
  NOR2X1 G5434 (.A1(W10095), .A2(W16317), .ZN(W33859));
  NOR2X1 G5435 (.A1(W8852), .A2(W1465), .ZN(W17049));
  NOR2X1 G5436 (.A1(W6836), .A2(W5156), .ZN(W33862));
  NOR2X1 G5437 (.A1(W19650), .A2(W18809), .ZN(O6913));
  NOR2X1 G5438 (.A1(W3541), .A2(W10031), .ZN(W19673));
  NOR2X1 G5439 (.A1(W26312), .A2(W6807), .ZN(O6908));
  NOR2X1 G5440 (.A1(W27540), .A2(W32887), .ZN(W33832));
  NOR2X1 G5441 (.A1(W32661), .A2(W20566), .ZN(O6912));
  NOR2X1 G5442 (.A1(W4986), .A2(W10900), .ZN(O1312));
  NOR2X1 G5443 (.A1(W1439), .A2(W27968), .ZN(W33835));
  NOR2X1 G5444 (.A1(W25890), .A2(W31055), .ZN(W33836));
  NOR2X1 G5445 (.A1(W2886), .A2(W11357), .ZN(W19675));
  NOR2X1 G5446 (.A1(W9273), .A2(W30201), .ZN(O6965));
  NOR2X1 G5447 (.A1(W14029), .A2(W2599), .ZN(W17076));
  NOR2X1 G5448 (.A1(W5063), .A2(W9936), .ZN(W33841));
  NOR2X1 G5449 (.A1(W2016), .A2(W6345), .ZN(O1311));
  NOR2X1 G5450 (.A1(I32), .A2(W10316), .ZN(W17072));
  NOR2X1 G5451 (.A1(W14615), .A2(W8189), .ZN(W17071));
  NOR2X1 G5452 (.A1(W14233), .A2(W16834), .ZN(O5668));
  NOR2X1 G5453 (.A1(W9262), .A2(W5033), .ZN(O1309));
  NOR2X1 G5454 (.A1(W6652), .A2(W7095), .ZN(W16863));
  NOR2X1 G5455 (.A1(W9087), .A2(I1972), .ZN(W19743));
  NOR2X1 G5456 (.A1(W9352), .A2(W5806), .ZN(W16871));
  NOR2X1 G5457 (.A1(I1614), .A2(W14646), .ZN(O5638));
  NOR2X1 G5458 (.A1(W22384), .A2(W6729), .ZN(W31086));
  NOR2X1 G5459 (.A1(W7716), .A2(I968), .ZN(W16868));
  NOR2X1 G5460 (.A1(W14267), .A2(W15430), .ZN(W34033));
  NOR2X1 G5461 (.A1(I313), .A2(W7935), .ZN(O1841));
  NOR2X1 G5462 (.A1(W6613), .A2(W16706), .ZN(O1842));
  NOR2X1 G5463 (.A1(W15265), .A2(W21353), .ZN(O7025));
  NOR2X1 G5464 (.A1(W5144), .A2(W3478), .ZN(W16862));
  NOR2X1 G5465 (.A1(W11259), .A2(W9141), .ZN(W19749));
  NOR2X1 G5466 (.A1(W7357), .A2(W6178), .ZN(W19750));
  NOR2X1 G5467 (.A1(W32740), .A2(W28509), .ZN(W34041));
  NOR2X1 G5468 (.A1(W9105), .A2(W11660), .ZN(O5637));
  NOR2X1 G5469 (.A1(W6444), .A2(W13930), .ZN(W16857));
  NOR2X1 G5470 (.A1(W27316), .A2(W14012), .ZN(O7033));
  NOR2X1 G5471 (.A1(W11900), .A2(W13875), .ZN(O1844));
  NOR2X1 G5472 (.A1(I1333), .A2(W5541), .ZN(W16882));
  NOR2X1 G5473 (.A1(W1367), .A2(W10050), .ZN(W16890));
  NOR2X1 G5474 (.A1(W14556), .A2(W10404), .ZN(O5642));
  NOR2X1 G5475 (.A1(W9702), .A2(W10957), .ZN(W16888));
  NOR2X1 G5476 (.A1(W12230), .A2(W30453), .ZN(W31093));
  NOR2X1 G5477 (.A1(W9619), .A2(W19146), .ZN(W34013));
  NOR2X1 G5478 (.A1(W7366), .A2(W11123), .ZN(W16885));
  NOR2X1 G5479 (.A1(W4121), .A2(W5997), .ZN(W16884));
  NOR2X1 G5480 (.A1(W25158), .A2(W2699), .ZN(O5640));
  NOR2X1 G5481 (.A1(W3204), .A2(W8975), .ZN(W16854));
  NOR2X1 G5482 (.A1(W21806), .A2(W14575), .ZN(O7013));
  NOR2X1 G5483 (.A1(W15746), .A2(W21321), .ZN(W31090));
  NOR2X1 G5484 (.A1(W7894), .A2(I772), .ZN(W16879));
  NOR2X1 G5485 (.A1(W6076), .A2(W11196), .ZN(W16878));
  NOR2X1 G5486 (.A1(W11150), .A2(W3380), .ZN(W16877));
  NOR2X1 G5487 (.A1(W13531), .A2(W21620), .ZN(O5639));
  NOR2X1 G5488 (.A1(W32396), .A2(W12813), .ZN(O7022));
  NOR2X1 G5489 (.A1(W124), .A2(W9796), .ZN(O7051));
  NOR2X1 G5490 (.A1(W4277), .A2(W9402), .ZN(O1272));
  NOR2X1 G5491 (.A1(W28612), .A2(I1927), .ZN(O7044));
  NOR2X1 G5492 (.A1(W32635), .A2(W3011), .ZN(O7045));
  NOR2X1 G5493 (.A1(W32055), .A2(W1391), .ZN(O7046));
  NOR2X1 G5494 (.A1(W4279), .A2(W5046), .ZN(W16831));
  NOR2X1 G5495 (.A1(I1467), .A2(W5202), .ZN(W16830));
  NOR2X1 G5496 (.A1(W18903), .A2(W18931), .ZN(W19760));
  NOR2X1 G5497 (.A1(W9141), .A2(W14794), .ZN(W31072));
  NOR2X1 G5498 (.A1(W4678), .A2(W15875), .ZN(W16837));
  NOR2X1 G5499 (.A1(W19771), .A2(W9157), .ZN(O7052));
  NOR2X1 G5500 (.A1(W1430), .A2(W6497), .ZN(W16824));
  NOR2X1 G5501 (.A1(W9273), .A2(W18840), .ZN(W19763));
  NOR2X1 G5502 (.A1(I1415), .A2(W24530), .ZN(O7054));
  NOR2X1 G5503 (.A1(W14926), .A2(W17817), .ZN(O5632));
  NOR2X1 G5504 (.A1(W14160), .A2(W911), .ZN(W16819));
  NOR2X1 G5505 (.A1(W19645), .A2(W22009), .ZN(W34079));
  NOR2X1 G5506 (.A1(W22269), .A2(W31096), .ZN(O7057));
  NOR2X1 G5507 (.A1(W4585), .A2(W29314), .ZN(O7036));
  NOR2X1 G5508 (.A1(W13550), .A2(W9781), .ZN(W16853));
  NOR2X1 G5509 (.A1(W14695), .A2(W5934), .ZN(O7035));
  NOR2X1 G5510 (.A1(W8294), .A2(W1034), .ZN(O5636));
  NOR2X1 G5511 (.A1(W79), .A2(W12643), .ZN(O1845));
  NOR2X1 G5512 (.A1(W9309), .A2(W31797), .ZN(W34050));
  NOR2X1 G5513 (.A1(W13866), .A2(W2183), .ZN(W16848));
  NOR2X1 G5514 (.A1(W13608), .A2(W2648), .ZN(W16847));
  NOR2X1 G5515 (.A1(W5353), .A2(W6195), .ZN(W16846));
  NOR2X1 G5516 (.A1(W4607), .A2(I1626), .ZN(O1275));
  NOR2X1 G5517 (.A1(W2657), .A2(I793), .ZN(W16844));
  NOR2X1 G5518 (.A1(W15336), .A2(W4734), .ZN(W16843));
  NOR2X1 G5519 (.A1(W7216), .A2(W14947), .ZN(W16842));
  NOR2X1 G5520 (.A1(W22282), .A2(W21122), .ZN(W31081));
  NOR2X1 G5521 (.A1(W2826), .A2(W18918), .ZN(W19756));
  NOR2X1 G5522 (.A1(W14085), .A2(W1054), .ZN(W31080));
  NOR2X1 G5523 (.A1(W20132), .A2(W8196), .ZN(O5634));
  NOR2X1 G5524 (.A1(W4153), .A2(W3268), .ZN(W19718));
  NOR2X1 G5525 (.A1(W4863), .A2(W2116), .ZN(O1287));
  NOR2X1 G5526 (.A1(W170), .A2(W28101), .ZN(O6977));
  NOR2X1 G5527 (.A1(W19208), .A2(W9093), .ZN(O6978));
  NOR2X1 G5528 (.A1(W792), .A2(W1361), .ZN(W16947));
  NOR2X1 G5529 (.A1(W4319), .A2(W4679), .ZN(W16946));
  NOR2X1 G5530 (.A1(W3774), .A2(W19162), .ZN(W19717));
  NOR2X1 G5531 (.A1(W11251), .A2(W6824), .ZN(W16944));
  NOR2X1 G5532 (.A1(W17411), .A2(W12573), .ZN(W33959));
  NOR2X1 G5533 (.A1(W5503), .A2(W15212), .ZN(O6976));
  NOR2X1 G5534 (.A1(W5489), .A2(W14083), .ZN(W16941));
  NOR2X1 G5535 (.A1(W26267), .A2(W18286), .ZN(W31112));
  NOR2X1 G5536 (.A1(W22626), .A2(W2518), .ZN(O6981));
  NOR2X1 G5537 (.A1(W9136), .A2(W15291), .ZN(W16938));
  NOR2X1 G5538 (.A1(W14320), .A2(W4954), .ZN(W16937));
  NOR2X1 G5539 (.A1(W18657), .A2(I1553), .ZN(W19720));
  NOR2X1 G5540 (.A1(I338), .A2(W8016), .ZN(W16934));
  NOR2X1 G5541 (.A1(W13355), .A2(W8374), .ZN(O6985));
  NOR2X1 G5542 (.A1(W18252), .A2(W16352), .ZN(W31116));
  NOR2X1 G5543 (.A1(W6044), .A2(W4659), .ZN(W16969));
  NOR2X1 G5544 (.A1(W3083), .A2(W11272), .ZN(O1290));
  NOR2X1 G5545 (.A1(W20439), .A2(W7588), .ZN(W31125));
  NOR2X1 G5546 (.A1(W23510), .A2(W15744), .ZN(W31124));
  NOR2X1 G5547 (.A1(W17408), .A2(W19068), .ZN(O6966));
  NOR2X1 G5548 (.A1(W3868), .A2(W11088), .ZN(O6969));
  NOR2X1 G5549 (.A1(W13752), .A2(W5842), .ZN(W16961));
  NOR2X1 G5550 (.A1(W12623), .A2(W11933), .ZN(W33945));
  NOR2X1 G5551 (.A1(W182), .A2(W2504), .ZN(W19722));
  NOR2X1 G5552 (.A1(W4748), .A2(W7670), .ZN(W16958));
  NOR2X1 G5553 (.A1(W12866), .A2(W14538), .ZN(W19715));
  NOR2X1 G5554 (.A1(W10810), .A2(I1941), .ZN(O6972));
  NOR2X1 G5555 (.A1(W8800), .A2(W13625), .ZN(W16955));
  NOR2X1 G5556 (.A1(W23754), .A2(I164), .ZN(W31114));
  NOR2X1 G5557 (.A1(W26080), .A2(W2685), .ZN(W33952));
  NOR2X1 G5558 (.A1(W435), .A2(W419), .ZN(O6975));
  NOR2X1 G5559 (.A1(W9706), .A2(W12437), .ZN(W19733));
  NOR2X1 G5560 (.A1(W11604), .A2(W2595), .ZN(W31105));
  NOR2X1 G5561 (.A1(I1505), .A2(W30556), .ZN(W33988));
  NOR2X1 G5562 (.A1(W20132), .A2(W29445), .ZN(O7001));
  NOR2X1 G5563 (.A1(W4803), .A2(I1388), .ZN(W16909));
  NOR2X1 G5564 (.A1(W4328), .A2(W4263), .ZN(W16908));
  NOR2X1 G5565 (.A1(W18499), .A2(W14025), .ZN(O1836));
  NOR2X1 G5566 (.A1(W3510), .A2(W11958), .ZN(W33997));
  NOR2X1 G5567 (.A1(W13566), .A2(W6568), .ZN(O1279));
  NOR2X1 G5568 (.A1(W16886), .A2(W26559), .ZN(O6997));
  NOR2X1 G5569 (.A1(W16446), .A2(W574), .ZN(O1277));
  NOR2X1 G5570 (.A1(W12478), .A2(W16677), .ZN(W16899));
  NOR2X1 G5571 (.A1(W13290), .A2(I1149), .ZN(O7007));
  NOR2X1 G5572 (.A1(W5093), .A2(W9383), .ZN(W16897));
  NOR2X1 G5573 (.A1(W4855), .A2(I1755), .ZN(W16895));
  NOR2X1 G5574 (.A1(W2928), .A2(W11754), .ZN(O1839));
  NOR2X1 G5575 (.A1(W10125), .A2(W30935), .ZN(W34008));
  NOR2X1 G5576 (.A1(W8660), .A2(I334), .ZN(O6995));
  NOR2X1 G5577 (.A1(W4987), .A2(W12376), .ZN(W16931));
  NOR2X1 G5578 (.A1(W27770), .A2(I1672), .ZN(O6988));
  NOR2X1 G5579 (.A1(W22139), .A2(W21031), .ZN(O6989));
  NOR2X1 G5580 (.A1(W16668), .A2(W1628), .ZN(W16927));
  NOR2X1 G5581 (.A1(W6524), .A2(W4207), .ZN(W19724));
  NOR2X1 G5582 (.A1(W30688), .A2(W28611), .ZN(O6994));
  NOR2X1 G5583 (.A1(W16323), .A2(W9441), .ZN(O1284));
  NOR2X1 G5584 (.A1(W12608), .A2(W907), .ZN(W16923));
  NOR2X1 G5585 (.A1(W26982), .A2(W11286), .ZN(W31395));
  NOR2X1 G5586 (.A1(W13938), .A2(I192), .ZN(O1283));
  NOR2X1 G5587 (.A1(W1631), .A2(W5392), .ZN(O1282));
  NOR2X1 G5588 (.A1(W14809), .A2(W1859), .ZN(W16919));
  NOR2X1 G5589 (.A1(W12403), .A2(W11115), .ZN(W16918));
  NOR2X1 G5590 (.A1(W10264), .A2(W21453), .ZN(O5647));
  NOR2X1 G5591 (.A1(W5405), .A2(W9387), .ZN(O1281));
  NOR2X1 G5592 (.A1(W3895), .A2(W17459), .ZN(W19726));
  NOR2X1 G5593 (.A1(W5811), .A2(W15893), .ZN(W18598));
  NOR2X1 G5594 (.A1(W13311), .A2(W13867), .ZN(W18609));
  NOR2X1 G5595 (.A1(W26499), .A2(W27857), .ZN(W32228));
  NOR2X1 G5596 (.A1(I319), .A2(W20904), .ZN(O6153));
  NOR2X1 G5597 (.A1(W13194), .A2(W97), .ZN(W19130));
  NOR2X1 G5598 (.A1(W2150), .A2(W13600), .ZN(W32234));
  NOR2X1 G5599 (.A1(W4684), .A2(W31371), .ZN(O5902));
  NOR2X1 G5600 (.A1(W3661), .A2(W17763), .ZN(W32238));
  NOR2X1 G5601 (.A1(I1332), .A2(W18899), .ZN(W32240));
  NOR2X1 G5602 (.A1(W10327), .A2(I1184), .ZN(W18610));
  NOR2X1 G5603 (.A1(W13888), .A2(W10024), .ZN(O6158));
  NOR2X1 G5604 (.A1(W3340), .A2(W1255), .ZN(W19135));
  NOR2X1 G5605 (.A1(W14173), .A2(W29945), .ZN(O6160));
  NOR2X1 G5606 (.A1(W3679), .A2(W16682), .ZN(O1597));
  NOR2X1 G5607 (.A1(W1764), .A2(W3533), .ZN(W19136));
  NOR2X1 G5608 (.A1(W16252), .A2(W17737), .ZN(W19137));
  NOR2X1 G5609 (.A1(W19165), .A2(W1729), .ZN(O5901));
  NOR2X1 G5610 (.A1(W11145), .A2(W21316), .ZN(O6163));
  NOR2X1 G5611 (.A1(W9083), .A2(I1642), .ZN(O1604));
  NOR2X1 G5612 (.A1(W7742), .A2(W26875), .ZN(W32214));
  NOR2X1 G5613 (.A1(W711), .A2(W7661), .ZN(O1606));
  NOR2X1 G5614 (.A1(W17884), .A2(W16829), .ZN(O1605));
  NOR2X1 G5615 (.A1(W29659), .A2(W6958), .ZN(W32215));
  NOR2X1 G5616 (.A1(W8095), .A2(W5085), .ZN(O1710));
  NOR2X1 G5617 (.A1(W13212), .A2(W13607), .ZN(W18622));
  NOR2X1 G5618 (.A1(W31019), .A2(W9298), .ZN(O6147));
  NOR2X1 G5619 (.A1(W18621), .A2(W9078), .ZN(O6148));
  NOR2X1 G5620 (.A1(W9887), .A2(W6873), .ZN(W18587));
  NOR2X1 G5621 (.A1(W3323), .A2(W781), .ZN(W18618));
  NOR2X1 G5622 (.A1(W7771), .A2(W4195), .ZN(W32224));
  NOR2X1 G5623 (.A1(W1115), .A2(W6556), .ZN(W18615));
  NOR2X1 G5624 (.A1(W17418), .A2(W5362), .ZN(W18614));
  NOR2X1 G5625 (.A1(W6569), .A2(W21920), .ZN(W31710));
  NOR2X1 G5626 (.A1(W1828), .A2(W7009), .ZN(W18612));
  NOR2X1 G5627 (.A1(W660), .A2(W31056), .ZN(W32227));
  NOR2X1 G5628 (.A1(W17389), .A2(W17297), .ZN(O5899));
  NOR2X1 G5629 (.A1(W17486), .A2(I184), .ZN(W18568));
  NOR2X1 G5630 (.A1(W19742), .A2(W2254), .ZN(O6168));
  NOR2X1 G5631 (.A1(W13427), .A2(W15296), .ZN(W18566));
  NOR2X1 G5632 (.A1(W18345), .A2(W19834), .ZN(W32268));
  NOR2X1 G5633 (.A1(W9711), .A2(W16422), .ZN(W19145));
  NOR2X1 G5634 (.A1(W1602), .A2(W16324), .ZN(W18563));
  NOR2X1 G5635 (.A1(W2918), .A2(W9062), .ZN(W18562));
  NOR2X1 G5636 (.A1(W4177), .A2(W2175), .ZN(W18561));
  NOR2X1 G5637 (.A1(W7628), .A2(W9622), .ZN(W18569));
  NOR2X1 G5638 (.A1(W16524), .A2(W14646), .ZN(O1587));
  NOR2X1 G5639 (.A1(W10512), .A2(I1896), .ZN(O1715));
  NOR2X1 G5640 (.A1(W3905), .A2(W16516), .ZN(W19148));
  NOR2X1 G5641 (.A1(W19928), .A2(W15543), .ZN(W32276));
  NOR2X1 G5642 (.A1(W5087), .A2(I560), .ZN(W32278));
  NOR2X1 G5643 (.A1(W27352), .A2(W20553), .ZN(W32279));
  NOR2X1 G5644 (.A1(W6832), .A2(W14541), .ZN(W19149));
  NOR2X1 G5645 (.A1(W2128), .A2(W15048), .ZN(W18552));
  NOR2X1 G5646 (.A1(W14870), .A2(W1035), .ZN(W19140));
  NOR2X1 G5647 (.A1(W1603), .A2(W3170), .ZN(W18586));
  NOR2X1 G5648 (.A1(W32066), .A2(I1853), .ZN(W32253));
  NOR2X1 G5649 (.A1(W10551), .A2(W869), .ZN(O1593));
  NOR2X1 G5650 (.A1(W7359), .A2(W12979), .ZN(W18583));
  NOR2X1 G5651 (.A1(W8411), .A2(W14021), .ZN(O1592));
  NOR2X1 G5652 (.A1(W7399), .A2(W9914), .ZN(W19139));
  NOR2X1 G5653 (.A1(W3879), .A2(W1568), .ZN(W18580));
  NOR2X1 G5654 (.A1(W2745), .A2(W10230), .ZN(W18579));
  NOR2X1 G5655 (.A1(W2064), .A2(W29416), .ZN(O5905));
  NOR2X1 G5656 (.A1(W7121), .A2(W1277), .ZN(O1714));
  NOR2X1 G5657 (.A1(W24677), .A2(W20259), .ZN(W32259));
  NOR2X1 G5658 (.A1(W2610), .A2(W10806), .ZN(O1590));
  NOR2X1 G5659 (.A1(W28697), .A2(W26856), .ZN(W32260));
  NOR2X1 G5660 (.A1(W12241), .A2(W6737), .ZN(W31698));
  NOR2X1 G5661 (.A1(W17373), .A2(W13279), .ZN(O6167));
  NOR2X1 G5662 (.A1(W31431), .A2(W29303), .ZN(W31695));
  NOR2X1 G5663 (.A1(W24328), .A2(W31675), .ZN(W32162));
  NOR2X1 G5664 (.A1(W14378), .A2(W5957), .ZN(O1621));
  NOR2X1 G5665 (.A1(W6129), .A2(W12635), .ZN(W18683));
  NOR2X1 G5666 (.A1(W5047), .A2(W16206), .ZN(W18682));
  NOR2X1 G5667 (.A1(W11447), .A2(W21084), .ZN(O6123));
  NOR2X1 G5668 (.A1(W12472), .A2(W1735), .ZN(W18679));
  NOR2X1 G5669 (.A1(W12233), .A2(W14929), .ZN(W32160));
  NOR2X1 G5670 (.A1(W5590), .A2(W3219), .ZN(O1619));
  NOR2X1 G5671 (.A1(W29464), .A2(W12582), .ZN(W31728));
  NOR2X1 G5672 (.A1(W5022), .A2(W10018), .ZN(W18685));
  NOR2X1 G5673 (.A1(W198), .A2(W11770), .ZN(O6125));
  NOR2X1 G5674 (.A1(W11649), .A2(W28626), .ZN(W31727));
  NOR2X1 G5675 (.A1(W28746), .A2(W14072), .ZN(W32165));
  NOR2X1 G5676 (.A1(W2751), .A2(W17418), .ZN(W32168));
  NOR2X1 G5677 (.A1(W8761), .A2(W13518), .ZN(W18670));
  NOR2X1 G5678 (.A1(W21135), .A2(W27324), .ZN(O5913));
  NOR2X1 G5679 (.A1(W16222), .A2(I782), .ZN(W18668));
  NOR2X1 G5680 (.A1(W5713), .A2(W7142), .ZN(O6128));
  NOR2X1 G5681 (.A1(W23657), .A2(W3459), .ZN(O6114));
  NOR2X1 G5682 (.A1(W8848), .A2(W30165), .ZN(O6107));
  NOR2X1 G5683 (.A1(W4360), .A2(W7842), .ZN(W18701));
  NOR2X1 G5684 (.A1(W30983), .A2(W3657), .ZN(O6108));
  NOR2X1 G5685 (.A1(W22364), .A2(W25750), .ZN(O6109));
  NOR2X1 G5686 (.A1(W24307), .A2(W23529), .ZN(O6110));
  NOR2X1 G5687 (.A1(W21648), .A2(W7406), .ZN(O6111));
  NOR2X1 G5688 (.A1(W5080), .A2(W15267), .ZN(O6112));
  NOR2X1 G5689 (.A1(W2358), .A2(W11297), .ZN(O5915));
  NOR2X1 G5690 (.A1(W2732), .A2(W5988), .ZN(W18666));
  NOR2X1 G5691 (.A1(I1041), .A2(W15949), .ZN(W18693));
  NOR2X1 G5692 (.A1(W16929), .A2(W8343), .ZN(W18692));
  NOR2X1 G5693 (.A1(W29196), .A2(W27857), .ZN(O6116));
  NOR2X1 G5694 (.A1(W10707), .A2(W18259), .ZN(W18690));
  NOR2X1 G5695 (.A1(W17263), .A2(W2761), .ZN(W18688));
  NOR2X1 G5696 (.A1(W1000), .A2(W19743), .ZN(W32151));
  NOR2X1 G5697 (.A1(W19170), .A2(W18141), .ZN(O6120));
  NOR2X1 G5698 (.A1(W19678), .A2(W3977), .ZN(W32201));
  NOR2X1 G5699 (.A1(W4990), .A2(W9686), .ZN(O1614));
  NOR2X1 G5700 (.A1(W3559), .A2(W15585), .ZN(O6138));
  NOR2X1 G5701 (.A1(W292), .A2(W6135), .ZN(O6139));
  NOR2X1 G5702 (.A1(W8568), .A2(W8741), .ZN(W32194));
  NOR2X1 G5703 (.A1(W5853), .A2(W21331), .ZN(O5909));
  NOR2X1 G5704 (.A1(W17839), .A2(W15096), .ZN(O5908));
  NOR2X1 G5705 (.A1(W31152), .A2(W21354), .ZN(W32199));
  NOR2X1 G5706 (.A1(W20759), .A2(W8838), .ZN(O6144));
  NOR2X1 G5707 (.A1(W15769), .A2(W18395), .ZN(W19116));
  NOR2X1 G5708 (.A1(W17145), .A2(W8259), .ZN(W18636));
  NOR2X1 G5709 (.A1(W16121), .A2(W13264), .ZN(O6145));
  NOR2X1 G5710 (.A1(W13927), .A2(W1383), .ZN(W32204));
  NOR2X1 G5711 (.A1(W11543), .A2(I1930), .ZN(W31715));
  NOR2X1 G5712 (.A1(W8937), .A2(W6226), .ZN(W32206));
  NOR2X1 G5713 (.A1(W6081), .A2(W25690), .ZN(W32210));
  NOR2X1 G5714 (.A1(W5104), .A2(W7364), .ZN(W18630));
  NOR2X1 G5715 (.A1(W3388), .A2(W2407), .ZN(O5907));
  NOR2X1 G5716 (.A1(W9952), .A2(W25406), .ZN(W32180));
  NOR2X1 G5717 (.A1(W11911), .A2(W10774), .ZN(W18665));
  NOR2X1 G5718 (.A1(W9570), .A2(W2417), .ZN(O1708));
  NOR2X1 G5719 (.A1(I1957), .A2(W1001), .ZN(W18663));
  NOR2X1 G5720 (.A1(W10848), .A2(W28675), .ZN(W31725));
  NOR2X1 G5721 (.A1(W856), .A2(W13076), .ZN(W19114));
  NOR2X1 G5722 (.A1(W4040), .A2(I358), .ZN(W18660));
  NOR2X1 G5723 (.A1(W5202), .A2(W7883), .ZN(W18659));
  NOR2X1 G5724 (.A1(W15669), .A2(W25741), .ZN(W32179));
  NOR2X1 G5725 (.A1(W6562), .A2(W9171), .ZN(W18551));
  NOR2X1 G5726 (.A1(W28997), .A2(W5921), .ZN(O6133));
  NOR2X1 G5727 (.A1(W17215), .A2(W6704), .ZN(W32182));
  NOR2X1 G5728 (.A1(W14780), .A2(W16035), .ZN(W18654));
  NOR2X1 G5729 (.A1(W12915), .A2(W17431), .ZN(W18653));
  NOR2X1 G5730 (.A1(W4467), .A2(W19979), .ZN(W32183));
  NOR2X1 G5731 (.A1(W14687), .A2(W5853), .ZN(W19115));
  NOR2X1 G5732 (.A1(W19724), .A2(W13619), .ZN(W32186));
  NOR2X1 G5733 (.A1(W15712), .A2(I230), .ZN(O6225));
  NOR2X1 G5734 (.A1(W17416), .A2(W27702), .ZN(W32396));
  NOR2X1 G5735 (.A1(W14610), .A2(W13096), .ZN(O5875));
  NOR2X1 G5736 (.A1(W1932), .A2(W3690), .ZN(O1569));
  NOR2X1 G5737 (.A1(W14042), .A2(W17842), .ZN(W19194));
  NOR2X1 G5738 (.A1(W15273), .A2(W4500), .ZN(W18446));
  NOR2X1 G5739 (.A1(W23928), .A2(W3698), .ZN(W31643));
  NOR2X1 G5740 (.A1(W7357), .A2(I423), .ZN(W18444));
  NOR2X1 G5741 (.A1(W214), .A2(W9605), .ZN(W18443));
  NOR2X1 G5742 (.A1(W18670), .A2(W25223), .ZN(W32395));
  NOR2X1 G5743 (.A1(W2010), .A2(W11348), .ZN(W18441));
  NOR2X1 G5744 (.A1(I1959), .A2(W11962), .ZN(O5871));
  NOR2X1 G5745 (.A1(W16432), .A2(W16357), .ZN(W19197));
  NOR2X1 G5746 (.A1(W7043), .A2(W6136), .ZN(W19199));
  NOR2X1 G5747 (.A1(W19311), .A2(W18246), .ZN(O6231));
  NOR2X1 G5748 (.A1(W23167), .A2(W738), .ZN(O5867));
  NOR2X1 G5749 (.A1(W6532), .A2(W23066), .ZN(W32419));
  NOR2X1 G5750 (.A1(W3026), .A2(W12747), .ZN(O1567));
  NOR2X1 G5751 (.A1(W18899), .A2(W29502), .ZN(O5878));
  NOR2X1 G5752 (.A1(I522), .A2(W5882), .ZN(O1572));
  NOR2X1 G5753 (.A1(W13759), .A2(W14810), .ZN(W18470));
  NOR2X1 G5754 (.A1(W16051), .A2(W26396), .ZN(W32369));
  NOR2X1 G5755 (.A1(W18493), .A2(I346), .ZN(O5879));
  NOR2X1 G5756 (.A1(W3827), .A2(W9203), .ZN(W18466));
  NOR2X1 G5757 (.A1(I169), .A2(I110), .ZN(W32377));
  NOR2X1 G5758 (.A1(W14416), .A2(W1904), .ZN(W19185));
  NOR2X1 G5759 (.A1(W24354), .A2(W7177), .ZN(W31656));
  NOR2X1 G5760 (.A1(W16337), .A2(W4475), .ZN(O1566));
  NOR2X1 G5761 (.A1(W14949), .A2(W23658), .ZN(W32382));
  NOR2X1 G5762 (.A1(W4637), .A2(W16554), .ZN(W18459));
  NOR2X1 G5763 (.A1(W31173), .A2(W8430), .ZN(O6217));
  NOR2X1 G5764 (.A1(W8988), .A2(W11966), .ZN(W19189));
  NOR2X1 G5765 (.A1(W4676), .A2(W17168), .ZN(O6219));
  NOR2X1 G5766 (.A1(W16052), .A2(W30497), .ZN(O5876));
  NOR2X1 G5767 (.A1(W12796), .A2(W390), .ZN(W18454));
  NOR2X1 G5768 (.A1(W4009), .A2(W16181), .ZN(W31622));
  NOR2X1 G5769 (.A1(W703), .A2(W10374), .ZN(W18407));
  NOR2X1 G5770 (.A1(I100), .A2(W1769), .ZN(W18406));
  NOR2X1 G5771 (.A1(W23194), .A2(W9834), .ZN(W31624));
  NOR2X1 G5772 (.A1(W13320), .A2(W26902), .ZN(W32450));
  NOR2X1 G5773 (.A1(W10411), .A2(W10014), .ZN(W18403));
  NOR2X1 G5774 (.A1(W2075), .A2(W170), .ZN(W18402));
  NOR2X1 G5775 (.A1(W3114), .A2(I66), .ZN(W18401));
  NOR2X1 G5776 (.A1(W17588), .A2(W13543), .ZN(W18400));
  NOR2X1 G5777 (.A1(W11387), .A2(W3858), .ZN(O6241));
  NOR2X1 G5778 (.A1(W14474), .A2(W24518), .ZN(W32454));
  NOR2X1 G5779 (.A1(W2640), .A2(W6969), .ZN(W19216));
  NOR2X1 G5780 (.A1(W4906), .A2(I352), .ZN(W18396));
  NOR2X1 G5781 (.A1(W14637), .A2(W3784), .ZN(W32459));
  NOR2X1 G5782 (.A1(W2217), .A2(W16869), .ZN(W19219));
  NOR2X1 G5783 (.A1(W1282), .A2(W13874), .ZN(O5861));
  NOR2X1 G5784 (.A1(W26599), .A2(W11199), .ZN(W32464));
  NOR2X1 G5785 (.A1(W8155), .A2(W6389), .ZN(W18389));
  NOR2X1 G5786 (.A1(W10235), .A2(W1942), .ZN(W32429));
  NOR2X1 G5787 (.A1(W5724), .A2(W28600), .ZN(W32421));
  NOR2X1 G5788 (.A1(W16461), .A2(W3722), .ZN(W31634));
  NOR2X1 G5789 (.A1(W12668), .A2(W11988), .ZN(W19204));
  NOR2X1 G5790 (.A1(W903), .A2(I606), .ZN(W18424));
  NOR2X1 G5791 (.A1(W8212), .A2(W9108), .ZN(W18423));
  NOR2X1 G5792 (.A1(W12526), .A2(W12810), .ZN(W18422));
  NOR2X1 G5793 (.A1(W15756), .A2(W4881), .ZN(O1564));
  NOR2X1 G5794 (.A1(W11179), .A2(W8998), .ZN(W32428));
  NOR2X1 G5795 (.A1(W3398), .A2(W9500), .ZN(W32366));
  NOR2X1 G5796 (.A1(W26399), .A2(W17657), .ZN(W32430));
  NOR2X1 G5797 (.A1(W6861), .A2(W12789), .ZN(W31628));
  NOR2X1 G5798 (.A1(W4012), .A2(W836), .ZN(W19210));
  NOR2X1 G5799 (.A1(W14694), .A2(W7496), .ZN(O1726));
  NOR2X1 G5800 (.A1(W167), .A2(W7136), .ZN(W19212));
  NOR2X1 G5801 (.A1(W30277), .A2(W17930), .ZN(W32444));
  NOR2X1 G5802 (.A1(W15487), .A2(W23763), .ZN(W32445));
  NOR2X1 G5803 (.A1(W14053), .A2(W17782), .ZN(W31682));
  NOR2X1 G5804 (.A1(W1755), .A2(I132), .ZN(W18532));
  NOR2X1 G5805 (.A1(W18096), .A2(W3894), .ZN(O1583));
  NOR2X1 G5806 (.A1(W13764), .A2(W10778), .ZN(W31687));
  NOR2X1 G5807 (.A1(W30276), .A2(W3195), .ZN(W31686));
  NOR2X1 G5808 (.A1(W24957), .A2(W30663), .ZN(O5893));
  NOR2X1 G5809 (.A1(I9), .A2(W9448), .ZN(W32303));
  NOR2X1 G5810 (.A1(W15078), .A2(W9228), .ZN(W18526));
  NOR2X1 G5811 (.A1(W16867), .A2(I442), .ZN(W31683));
  NOR2X1 G5812 (.A1(W25427), .A2(W17590), .ZN(O6177));
  NOR2X1 G5813 (.A1(W15370), .A2(W403), .ZN(O1578));
  NOR2X1 G5814 (.A1(W21041), .A2(W1435), .ZN(O5892));
  NOR2X1 G5815 (.A1(W3024), .A2(W14601), .ZN(W18521));
  NOR2X1 G5816 (.A1(W7095), .A2(W4782), .ZN(O1577));
  NOR2X1 G5817 (.A1(W16276), .A2(W30588), .ZN(W32309));
  NOR2X1 G5818 (.A1(W19030), .A2(W3005), .ZN(O6185));
  NOR2X1 G5819 (.A1(W6316), .A2(W9020), .ZN(W19163));
  NOR2X1 G5820 (.A1(W8408), .A2(W16776), .ZN(W18516));
  NOR2X1 G5821 (.A1(W6035), .A2(W7244), .ZN(O1584));
  NOR2X1 G5822 (.A1(W22630), .A2(I1144), .ZN(O6174));
  NOR2X1 G5823 (.A1(W19863), .A2(W19763), .ZN(O5898));
  NOR2X1 G5824 (.A1(W5009), .A2(W11369), .ZN(O1716));
  NOR2X1 G5825 (.A1(W5447), .A2(W9863), .ZN(W18547));
  NOR2X1 G5826 (.A1(W25160), .A2(W27333), .ZN(O6176));
  NOR2X1 G5827 (.A1(W14947), .A2(W12755), .ZN(W32288));
  NOR2X1 G5828 (.A1(W19077), .A2(W1027), .ZN(O5897));
  NOR2X1 G5829 (.A1(I294), .A2(W2158), .ZN(O1717));
  NOR2X1 G5830 (.A1(W21343), .A2(W168), .ZN(O6187));
  NOR2X1 G5831 (.A1(W15943), .A2(W13047), .ZN(W18540));
  NOR2X1 G5832 (.A1(W12869), .A2(W14304), .ZN(W31689));
  NOR2X1 G5833 (.A1(W13872), .A2(W13353), .ZN(W18538));
  NOR2X1 G5834 (.A1(W16291), .A2(W754), .ZN(W18537));
  NOR2X1 G5835 (.A1(W1787), .A2(W27062), .ZN(O5894));
  NOR2X1 G5836 (.A1(W22811), .A2(W12260), .ZN(W32295));
  NOR2X1 G5837 (.A1(W3438), .A2(W2856), .ZN(W18534));
  NOR2X1 G5838 (.A1(W462), .A2(W18627), .ZN(O5886));
  NOR2X1 G5839 (.A1(W3285), .A2(I1910), .ZN(W18493));
  NOR2X1 G5840 (.A1(W12587), .A2(W25777), .ZN(W32338));
  NOR2X1 G5841 (.A1(W14867), .A2(W32206), .ZN(O6199));
  NOR2X1 G5842 (.A1(W4924), .A2(W24391), .ZN(W32340));
  NOR2X1 G5843 (.A1(W10410), .A2(W1420), .ZN(O5887));
  NOR2X1 G5844 (.A1(W31948), .A2(W29340), .ZN(O6201));
  NOR2X1 G5845 (.A1(W1837), .A2(W12374), .ZN(O1723));
  NOR2X1 G5846 (.A1(W27627), .A2(W29677), .ZN(W32345));
  NOR2X1 G5847 (.A1(W19127), .A2(W14555), .ZN(O1722));
  NOR2X1 G5848 (.A1(W22324), .A2(W19207), .ZN(W32348));
  NOR2X1 G5849 (.A1(W28103), .A2(I1982), .ZN(O6203));
  NOR2X1 G5850 (.A1(W5622), .A2(W9866), .ZN(W18481));
  NOR2X1 G5851 (.A1(W18940), .A2(I1296), .ZN(O1724));
  NOR2X1 G5852 (.A1(W1364), .A2(W3888), .ZN(W18478));
  NOR2X1 G5853 (.A1(W1805), .A2(W10064), .ZN(W19179));
  NOR2X1 G5854 (.A1(W10582), .A2(W25049), .ZN(O6210));
  NOR2X1 G5855 (.A1(W6216), .A2(W2429), .ZN(W19181));
  NOR2X1 G5856 (.A1(W12906), .A2(I483), .ZN(O6189));
  NOR2X1 G5857 (.A1(W5028), .A2(W12256), .ZN(O1576));
  NOR2X1 G5858 (.A1(W13148), .A2(W28980), .ZN(W32313));
  NOR2X1 G5859 (.A1(W30626), .A2(W14187), .ZN(W32315));
  NOR2X1 G5860 (.A1(W10490), .A2(W1970), .ZN(W32316));
  NOR2X1 G5861 (.A1(W5986), .A2(W28607), .ZN(W32317));
  NOR2X1 G5862 (.A1(W15836), .A2(W14997), .ZN(W19164));
  NOR2X1 G5863 (.A1(W8972), .A2(W3029), .ZN(W19165));
  NOR2X1 G5864 (.A1(W18216), .A2(W31881), .ZN(W32321));
  NOR2X1 G5865 (.A1(W19012), .A2(W9240), .ZN(O5916));
  NOR2X1 G5866 (.A1(W2775), .A2(W6838), .ZN(W18505));
  NOR2X1 G5867 (.A1(W27694), .A2(W13424), .ZN(W31680));
  NOR2X1 G5868 (.A1(W20769), .A2(I512), .ZN(O6190));
  NOR2X1 G5869 (.A1(W9429), .A2(W11166), .ZN(O6193));
  NOR2X1 G5870 (.A1(I162), .A2(W17881), .ZN(W18500));
  NOR2X1 G5871 (.A1(W6332), .A2(W8093), .ZN(W31676));
  NOR2X1 G5872 (.A1(W15008), .A2(W14562), .ZN(W32333));
  NOR2X1 G5873 (.A1(I988), .A2(W14801), .ZN(W18913));
  NOR2X1 G5874 (.A1(W17239), .A2(W1318), .ZN(W31923));
  NOR2X1 G5875 (.A1(W10868), .A2(W11890), .ZN(W18922));
  NOR2X1 G5876 (.A1(W11284), .A2(W4750), .ZN(W18921));
  NOR2X1 G5877 (.A1(W18989), .A2(W27599), .ZN(O6013));
  NOR2X1 G5878 (.A1(W3631), .A2(W3078), .ZN(W18919));
  NOR2X1 G5879 (.A1(W18115), .A2(I633), .ZN(W18917));
  NOR2X1 G5880 (.A1(W2961), .A2(W30338), .ZN(W31929));
  NOR2X1 G5881 (.A1(W24751), .A2(W9190), .ZN(W31932));
  NOR2X1 G5882 (.A1(W30862), .A2(W11767), .ZN(O6011));
  NOR2X1 G5883 (.A1(W16851), .A2(W7431), .ZN(O1676));
  NOR2X1 G5884 (.A1(W10983), .A2(W14964), .ZN(W19044));
  NOR2X1 G5885 (.A1(W901), .A2(W9639), .ZN(O6017));
  NOR2X1 G5886 (.A1(W17909), .A2(W5825), .ZN(W18908));
  NOR2X1 G5887 (.A1(W12125), .A2(W20234), .ZN(O5950));
  NOR2X1 G5888 (.A1(W16332), .A2(W8910), .ZN(W31939));
  NOR2X1 G5889 (.A1(W13496), .A2(W6349), .ZN(W18905));
  NOR2X1 G5890 (.A1(W17295), .A2(W27890), .ZN(W31941));
  NOR2X1 G5891 (.A1(W8456), .A2(W3096), .ZN(W18933));
  NOR2X1 G5892 (.A1(W6668), .A2(W18094), .ZN(W31906));
  NOR2X1 G5893 (.A1(I1920), .A2(I1194), .ZN(W31908));
  NOR2X1 G5894 (.A1(W16225), .A2(W2177), .ZN(W18940));
  NOR2X1 G5895 (.A1(W2342), .A2(I144), .ZN(W18938));
  NOR2X1 G5896 (.A1(W20563), .A2(W9106), .ZN(O5957));
  NOR2X1 G5897 (.A1(W16471), .A2(W7252), .ZN(O1694));
  NOR2X1 G5898 (.A1(W14654), .A2(W10529), .ZN(W18935));
  NOR2X1 G5899 (.A1(W8048), .A2(W6600), .ZN(W18934));
  NOR2X1 G5900 (.A1(W33), .A2(W18555), .ZN(W18903));
  NOR2X1 G5901 (.A1(W22339), .A2(W8393), .ZN(W31913));
  NOR2X1 G5902 (.A1(W1120), .A2(W10071), .ZN(W19038));
  NOR2X1 G5903 (.A1(W18837), .A2(W19713), .ZN(W31915));
  NOR2X1 G5904 (.A1(W29442), .A2(I1020), .ZN(O5956));
  NOR2X1 G5905 (.A1(W469), .A2(W18537), .ZN(O6009));
  NOR2X1 G5906 (.A1(W20858), .A2(W8428), .ZN(O6010));
  NOR2X1 G5907 (.A1(W17400), .A2(W17493), .ZN(W18926));
  NOR2X1 G5908 (.A1(W14325), .A2(W4610), .ZN(W19052));
  NOR2X1 G5909 (.A1(W21641), .A2(W11852), .ZN(W31965));
  NOR2X1 G5910 (.A1(W17232), .A2(W9323), .ZN(W19050));
  NOR2X1 G5911 (.A1(W25871), .A2(W13581), .ZN(O6029));
  NOR2X1 G5912 (.A1(W22005), .A2(W29077), .ZN(W31972));
  NOR2X1 G5913 (.A1(W15693), .A2(W14420), .ZN(O1666));
  NOR2X1 G5914 (.A1(W11268), .A2(W17286), .ZN(W18878));
  NOR2X1 G5915 (.A1(W1753), .A2(W29926), .ZN(O6030));
  NOR2X1 G5916 (.A1(W30108), .A2(W30953), .ZN(O6032));
  NOR2X1 G5917 (.A1(I946), .A2(W532), .ZN(W31964));
  NOR2X1 G5918 (.A1(W13568), .A2(W17728), .ZN(W18873));
  NOR2X1 G5919 (.A1(W19976), .A2(W12157), .ZN(O6033));
  NOR2X1 G5920 (.A1(W27623), .A2(W29925), .ZN(O5947));
  NOR2X1 G5921 (.A1(I1364), .A2(W12106), .ZN(O6034));
  NOR2X1 G5922 (.A1(W4091), .A2(W15650), .ZN(O1663));
  NOR2X1 G5923 (.A1(I563), .A2(W829), .ZN(W18867));
  NOR2X1 G5924 (.A1(W14679), .A2(W1542), .ZN(W18866));
  NOR2X1 G5925 (.A1(W20386), .A2(W31910), .ZN(W31985));
  NOR2X1 G5926 (.A1(W25024), .A2(W14237), .ZN(W31953));
  NOR2X1 G5927 (.A1(W28520), .A2(W9058), .ZN(O6020));
  NOR2X1 G5928 (.A1(W12914), .A2(W11120), .ZN(W18901));
  NOR2X1 G5929 (.A1(W25421), .A2(W9344), .ZN(W31797));
  NOR2X1 G5930 (.A1(W13464), .A2(W1467), .ZN(W31948));
  NOR2X1 G5931 (.A1(W9931), .A2(W16297), .ZN(W18897));
  NOR2X1 G5932 (.A1(W19371), .A2(W11037), .ZN(W31951));
  NOR2X1 G5933 (.A1(W11526), .A2(W1113), .ZN(O1673));
  NOR2X1 G5934 (.A1(W15542), .A2(W7028), .ZN(O1672));
  NOR2X1 G5935 (.A1(W1068), .A2(I506), .ZN(W19034));
  NOR2X1 G5936 (.A1(I1421), .A2(W12140), .ZN(W18892));
  NOR2X1 G5937 (.A1(W18237), .A2(W17768), .ZN(W18891));
  NOR2X1 G5938 (.A1(W17391), .A2(W28735), .ZN(O5949));
  NOR2X1 G5939 (.A1(W4713), .A2(W542), .ZN(W18889));
  NOR2X1 G5940 (.A1(W18355), .A2(I483), .ZN(O6027));
  NOR2X1 G5941 (.A1(W327), .A2(W7865), .ZN(W18887));
  NOR2X1 G5942 (.A1(W12601), .A2(W4921), .ZN(W31962));
  NOR2X1 G5943 (.A1(W6792), .A2(W5743), .ZN(W18991));
  NOR2X1 G5944 (.A1(W17916), .A2(W18821), .ZN(O1689));
  NOR2X1 G5945 (.A1(W15913), .A2(W8319), .ZN(O1688));
  NOR2X1 G5946 (.A1(W713), .A2(W12608), .ZN(W18997));
  NOR2X1 G5947 (.A1(I387), .A2(W24542), .ZN(W31843));
  NOR2X1 G5948 (.A1(W6479), .A2(W9566), .ZN(W18995));
  NOR2X1 G5949 (.A1(W21210), .A2(W3679), .ZN(O5973));
  NOR2X1 G5950 (.A1(W12855), .A2(W10750), .ZN(W31847));
  NOR2X1 G5951 (.A1(W15624), .A2(W16436), .ZN(W18992));
  NOR2X1 G5952 (.A1(W14860), .A2(W5856), .ZN(W19000));
  NOR2X1 G5953 (.A1(W10989), .A2(W3017), .ZN(W18990));
  NOR2X1 G5954 (.A1(W19453), .A2(W30484), .ZN(W31848));
  NOR2X1 G5955 (.A1(W8180), .A2(W22835), .ZN(O5974));
  NOR2X1 G5956 (.A1(W15022), .A2(W4124), .ZN(O1687));
  NOR2X1 G5957 (.A1(W24292), .A2(W1303), .ZN(O5962));
  NOR2X1 G5958 (.A1(W5388), .A2(W12925), .ZN(W18985));
  NOR2X1 G5959 (.A1(W8036), .A2(W546), .ZN(W19023));
  NOR2X1 G5960 (.A1(W9431), .A2(W2387), .ZN(W19025));
  NOR2X1 G5961 (.A1(W6013), .A2(W17697), .ZN(O1691));
  NOR2X1 G5962 (.A1(W21277), .A2(W20148), .ZN(W31824));
  NOR2X1 G5963 (.A1(W6214), .A2(I284), .ZN(W19016));
  NOR2X1 G5964 (.A1(W13725), .A2(W10845), .ZN(W19018));
  NOR2X1 G5965 (.A1(W4995), .A2(W7037), .ZN(W19014));
  NOR2X1 G5966 (.A1(W15930), .A2(W23168), .ZN(O5966));
  NOR2X1 G5967 (.A1(W18000), .A2(W1109), .ZN(W31830));
  NOR2X1 G5968 (.A1(W24345), .A2(W14588), .ZN(W31831));
  NOR2X1 G5969 (.A1(W11836), .A2(W7063), .ZN(W19010));
  NOR2X1 G5970 (.A1(I1065), .A2(I494), .ZN(W18981));
  NOR2X1 G5971 (.A1(W29050), .A2(W15307), .ZN(O5963));
  NOR2X1 G5972 (.A1(W14265), .A2(W27492), .ZN(W31835));
  NOR2X1 G5973 (.A1(W90), .A2(W18736), .ZN(W19006));
  NOR2X1 G5974 (.A1(W22122), .A2(W23147), .ZN(W31836));
  NOR2X1 G5975 (.A1(W24154), .A2(W26065), .ZN(O5969));
  NOR2X1 G5976 (.A1(W1365), .A2(W14660), .ZN(W19020));
  NOR2X1 G5977 (.A1(W13316), .A2(W16048), .ZN(O1690));
  NOR2X1 G5978 (.A1(I614), .A2(W14690), .ZN(W18953));
  NOR2X1 G5979 (.A1(W3731), .A2(W16388), .ZN(W18961));
  NOR2X1 G5980 (.A1(W13836), .A2(W11165), .ZN(W18960));
  NOR2X1 G5981 (.A1(W15278), .A2(W28440), .ZN(O5996));
  NOR2X1 G5982 (.A1(W8770), .A2(W7634), .ZN(O1680));
  NOR2X1 G5983 (.A1(W10107), .A2(W3317), .ZN(W31884));
  NOR2X1 G5984 (.A1(W13394), .A2(W21807), .ZN(O5998));
  NOR2X1 G5985 (.A1(W14198), .A2(W11356), .ZN(W18955));
  NOR2X1 G5986 (.A1(W19323), .A2(W27595), .ZN(O5999));
  NOR2X1 G5987 (.A1(W1539), .A2(W27627), .ZN(O5995));
  NOR2X1 G5988 (.A1(W24709), .A2(W18688), .ZN(W31892));
  NOR2X1 G5989 (.A1(W25309), .A2(W17673), .ZN(W31896));
  NOR2X1 G5990 (.A1(W14839), .A2(W11145), .ZN(W19030));
  NOR2X1 G5991 (.A1(W1157), .A2(W13529), .ZN(W18948));
  NOR2X1 G5992 (.A1(W432), .A2(W1545), .ZN(W19032));
  NOR2X1 G5993 (.A1(W31120), .A2(W27361), .ZN(O5959));
  NOR2X1 G5994 (.A1(W30164), .A2(W14913), .ZN(O6004));
  NOR2X1 G5995 (.A1(W1468), .A2(W22558), .ZN(O6005));
  NOR2X1 G5996 (.A1(W18652), .A2(I1901), .ZN(W18971));
  NOR2X1 G5997 (.A1(W17513), .A2(W28633), .ZN(O5983));
  NOR2X1 G5998 (.A1(W1766), .A2(W8890), .ZN(O1684));
  NOR2X1 G5999 (.A1(W8107), .A2(W13572), .ZN(W18977));
  NOR2X1 G6000 (.A1(W11051), .A2(W4276), .ZN(W31863));
  NOR2X1 G6001 (.A1(W5934), .A2(W30248), .ZN(W31864));
  NOR2X1 G6002 (.A1(W18423), .A2(W6776), .ZN(W18974));
  NOR2X1 G6003 (.A1(W5166), .A2(I479), .ZN(W18973));
  NOR2X1 G6004 (.A1(W31687), .A2(W20888), .ZN(O5989));
  NOR2X1 G6005 (.A1(W1145), .A2(W23589), .ZN(O6035));
  NOR2X1 G6006 (.A1(W29302), .A2(W3834), .ZN(W31873));
  NOR2X1 G6007 (.A1(W27706), .A2(W26642), .ZN(W31874));
  NOR2X1 G6008 (.A1(W29116), .A2(W4909), .ZN(O5991));
  NOR2X1 G6009 (.A1(W6134), .A2(W18368), .ZN(W18966));
  NOR2X1 G6010 (.A1(W29481), .A2(I1992), .ZN(W31813));
  NOR2X1 G6011 (.A1(W4392), .A2(W1371), .ZN(W31877));
  NOR2X1 G6012 (.A1(W30616), .A2(W10039), .ZN(W31812));
  NOR2X1 G6013 (.A1(W18445), .A2(I1550), .ZN(W18751));
  NOR2X1 G6014 (.A1(W12680), .A2(W13735), .ZN(W18761));
  NOR2X1 G6015 (.A1(W14391), .A2(W21416), .ZN(W32089));
  NOR2X1 G6016 (.A1(W6902), .A2(W3902), .ZN(W18758));
  NOR2X1 G6017 (.A1(W32060), .A2(W14269), .ZN(W32090));
  NOR2X1 G6018 (.A1(W9880), .A2(W13744), .ZN(O1637));
  NOR2X1 G6019 (.A1(W182), .A2(W667), .ZN(O1636));
  NOR2X1 G6020 (.A1(W25112), .A2(W7154), .ZN(W32094));
  NOR2X1 G6021 (.A1(W18860), .A2(W7330), .ZN(W32095));
  NOR2X1 G6022 (.A1(W2893), .A2(W7192), .ZN(W18762));
  NOR2X1 G6023 (.A1(W3226), .A2(W5816), .ZN(W18750));
  NOR2X1 G6024 (.A1(W19699), .A2(W26283), .ZN(O5925));
  NOR2X1 G6025 (.A1(W26137), .A2(I1352), .ZN(O5924));
  NOR2X1 G6026 (.A1(W5036), .A2(W1570), .ZN(W18747));
  NOR2X1 G6027 (.A1(W1785), .A2(W12341), .ZN(W19092));
  NOR2X1 G6028 (.A1(I480), .A2(W17375), .ZN(W19093));
  NOR2X1 G6029 (.A1(W6377), .A2(W3288), .ZN(W18743));
  NOR2X1 G6030 (.A1(W4276), .A2(W13433), .ZN(W18742));
  NOR2X1 G6031 (.A1(W2340), .A2(W4285), .ZN(W18771));
  NOR2X1 G6032 (.A1(W16794), .A2(W8), .ZN(W18781));
  NOR2X1 G6033 (.A1(W2320), .A2(W12315), .ZN(W18779));
  NOR2X1 G6034 (.A1(W15646), .A2(W12299), .ZN(W19081));
  NOR2X1 G6035 (.A1(W22823), .A2(W1887), .ZN(O6079));
  NOR2X1 G6036 (.A1(W12470), .A2(W14558), .ZN(O6080));
  NOR2X1 G6037 (.A1(W16003), .A2(W24093), .ZN(W32074));
  NOR2X1 G6038 (.A1(W13815), .A2(W12484), .ZN(W19082));
  NOR2X1 G6039 (.A1(W5238), .A2(W20767), .ZN(O6081));
  NOR2X1 G6040 (.A1(W20892), .A2(W31510), .ZN(W31746));
  NOR2X1 G6041 (.A1(W12155), .A2(W585), .ZN(W19083));
  NOR2X1 G6042 (.A1(W21221), .A2(W7797), .ZN(W32078));
  NOR2X1 G6043 (.A1(W13378), .A2(W16192), .ZN(O1702));
  NOR2X1 G6044 (.A1(W18877), .A2(W2635), .ZN(W32081));
  NOR2X1 G6045 (.A1(W14905), .A2(I1353), .ZN(W32083));
  NOR2X1 G6046 (.A1(W25131), .A2(W27429), .ZN(W31753));
  NOR2X1 G6047 (.A1(W16578), .A2(W7333), .ZN(W32085));
  NOR2X1 G6048 (.A1(W9453), .A2(W7253), .ZN(W19101));
  NOR2X1 G6049 (.A1(W11091), .A2(W14019), .ZN(W32120));
  NOR2X1 G6050 (.A1(W6444), .A2(W8192), .ZN(O1629));
  NOR2X1 G6051 (.A1(W8908), .A2(W4963), .ZN(W18719));
  NOR2X1 G6052 (.A1(W10572), .A2(W18544), .ZN(W18718));
  NOR2X1 G6053 (.A1(W3185), .A2(W2925), .ZN(W19100));
  NOR2X1 G6054 (.A1(W22006), .A2(W170), .ZN(W32122));
  NOR2X1 G6055 (.A1(W5421), .A2(W5727), .ZN(W18715));
  NOR2X1 G6056 (.A1(W3214), .A2(W13301), .ZN(W32123));
  NOR2X1 G6057 (.A1(W5887), .A2(I291), .ZN(W18722));
  NOR2X1 G6058 (.A1(W11087), .A2(W11069), .ZN(W32125));
  NOR2X1 G6059 (.A1(W10367), .A2(W9276), .ZN(O6101));
  NOR2X1 G6060 (.A1(W7590), .A2(W20712), .ZN(W32129));
  NOR2X1 G6061 (.A1(W16013), .A2(W13029), .ZN(W19103));
  NOR2X1 G6062 (.A1(W28050), .A2(W15368), .ZN(W32132));
  NOR2X1 G6063 (.A1(W1560), .A2(W15800), .ZN(W18706));
  NOR2X1 G6064 (.A1(I1887), .A2(W24599), .ZN(O6104));
  NOR2X1 G6065 (.A1(W16640), .A2(W14057), .ZN(W19104));
  NOR2X1 G6066 (.A1(W16232), .A2(W5495), .ZN(W18730));
  NOR2X1 G6067 (.A1(W295), .A2(W12073), .ZN(W18739));
  NOR2X1 G6068 (.A1(W23440), .A2(W3720), .ZN(W31743));
  NOR2X1 G6069 (.A1(W28810), .A2(W15313), .ZN(W31735));
  NOR2X1 G6070 (.A1(W16679), .A2(W6143), .ZN(W18735));
  NOR2X1 G6071 (.A1(W20607), .A2(W11423), .ZN(W32111));
  NOR2X1 G6072 (.A1(W13828), .A2(W9430), .ZN(W18733));
  NOR2X1 G6073 (.A1(W2044), .A2(W26265), .ZN(W32112));
  NOR2X1 G6074 (.A1(W23941), .A2(W17763), .ZN(O6096));
  NOR2X1 G6075 (.A1(W14237), .A2(W22255), .ZN(O6076));
  NOR2X1 G6076 (.A1(W6791), .A2(W4969), .ZN(W19099));
  NOR2X1 G6077 (.A1(W18095), .A2(I983), .ZN(W18728));
  NOR2X1 G6078 (.A1(W2372), .A2(W12996), .ZN(W32115));
  NOR2X1 G6079 (.A1(W7978), .A2(W15210), .ZN(W18726));
  NOR2X1 G6080 (.A1(W6132), .A2(W2644), .ZN(W32116));
  NOR2X1 G6081 (.A1(W7996), .A2(W27435), .ZN(W32118));
  NOR2X1 G6082 (.A1(W16203), .A2(W9335), .ZN(W18723));
  NOR2X1 G6083 (.A1(W11708), .A2(I1274), .ZN(W19065));
  NOR2X1 G6084 (.A1(W15820), .A2(W17178), .ZN(O5941));
  NOR2X1 G6085 (.A1(W22341), .A2(W3787), .ZN(O6050));
  NOR2X1 G6086 (.A1(W4243), .A2(W10146), .ZN(W32011));
  NOR2X1 G6087 (.A1(W11303), .A2(W23364), .ZN(O6052));
  NOR2X1 G6088 (.A1(W8830), .A2(W16943), .ZN(O1659));
  NOR2X1 G6089 (.A1(W4434), .A2(I793), .ZN(W32013));
  NOR2X1 G6090 (.A1(W2927), .A2(W16894), .ZN(O1657));
  NOR2X1 G6091 (.A1(W2956), .A2(W19984), .ZN(O6054));
  NOR2X1 G6092 (.A1(W7324), .A2(W10816), .ZN(W18843));
  NOR2X1 G6093 (.A1(W8629), .A2(W2880), .ZN(O6058));
  NOR2X1 G6094 (.A1(I1425), .A2(W8807), .ZN(W18828));
  NOR2X1 G6095 (.A1(W5255), .A2(W10780), .ZN(W18826));
  NOR2X1 G6096 (.A1(W6670), .A2(W24529), .ZN(W31771));
  NOR2X1 G6097 (.A1(W5916), .A2(W8740), .ZN(O5935));
  NOR2X1 G6098 (.A1(W909), .A2(W18939), .ZN(O6064));
  NOR2X1 G6099 (.A1(W29405), .A2(W18818), .ZN(W32032));
  NOR2X1 G6100 (.A1(W6659), .A2(W3935), .ZN(W32033));
  NOR2X1 G6101 (.A1(W11322), .A2(W18084), .ZN(W18853));
  NOR2X1 G6102 (.A1(W3356), .A2(W19584), .ZN(O5944));
  NOR2X1 G6103 (.A1(W16118), .A2(W3559), .ZN(W18861));
  NOR2X1 G6104 (.A1(I480), .A2(W4043), .ZN(W18860));
  NOR2X1 G6105 (.A1(W31850), .A2(W31182), .ZN(W31989));
  NOR2X1 G6106 (.A1(W18205), .A2(W11750), .ZN(W18858));
  NOR2X1 G6107 (.A1(W16757), .A2(W16045), .ZN(W18857));
  NOR2X1 G6108 (.A1(W14114), .A2(W11680), .ZN(O6038));
  NOR2X1 G6109 (.A1(W16662), .A2(I728), .ZN(O1661));
  NOR2X1 G6110 (.A1(W6667), .A2(W28971), .ZN(W32034));
  NOR2X1 G6111 (.A1(W2236), .A2(W315), .ZN(W31783));
  NOR2X1 G6112 (.A1(W11818), .A2(W18457), .ZN(O6042));
  NOR2X1 G6113 (.A1(I1825), .A2(I182), .ZN(W31998));
  NOR2X1 G6114 (.A1(W1484), .A2(W3246), .ZN(W18848));
  NOR2X1 G6115 (.A1(W28386), .A2(W14624), .ZN(O6046));
  NOR2X1 G6116 (.A1(W17931), .A2(W15995), .ZN(W18845));
  NOR2X1 G6117 (.A1(W11614), .A2(W13446), .ZN(W19061));
  NOR2X1 G6118 (.A1(I501), .A2(I1015), .ZN(W18790));
  NOR2X1 G6119 (.A1(W14937), .A2(W5187), .ZN(W18799));
  NOR2X1 G6120 (.A1(W26273), .A2(W11051), .ZN(O5932));
  NOR2X1 G6121 (.A1(W274), .A2(W3445), .ZN(W18797));
  NOR2X1 G6122 (.A1(W12337), .A2(W15331), .ZN(W18796));
  NOR2X1 G6123 (.A1(W28366), .A2(W351), .ZN(W32055));
  NOR2X1 G6124 (.A1(W9515), .A2(W8639), .ZN(W19077));
  NOR2X1 G6125 (.A1(W10134), .A2(W608), .ZN(W18792));
  NOR2X1 G6126 (.A1(W17071), .A2(W13897), .ZN(W18791));
  NOR2X1 G6127 (.A1(W18546), .A2(W321), .ZN(W32051));
  NOR2X1 G6128 (.A1(W14207), .A2(W11399), .ZN(W18789));
  NOR2X1 G6129 (.A1(W14433), .A2(I315), .ZN(W18788));
  NOR2X1 G6130 (.A1(W12180), .A2(W22939), .ZN(O6073));
  NOR2X1 G6131 (.A1(W25323), .A2(W17984), .ZN(O6075));
  NOR2X1 G6132 (.A1(W13347), .A2(W4094), .ZN(W32064));
  NOR2X1 G6133 (.A1(W5231), .A2(W2345), .ZN(W19078));
  NOR2X1 G6134 (.A1(W12233), .A2(W16509), .ZN(W18783));
  NOR2X1 G6135 (.A1(W14548), .A2(W10157), .ZN(W18810));
  NOR2X1 G6136 (.A1(W379), .A2(W2970), .ZN(W18818));
  NOR2X1 G6137 (.A1(W5914), .A2(W2438), .ZN(O6065));
  NOR2X1 G6138 (.A1(I226), .A2(W24716), .ZN(O6066));
  NOR2X1 G6139 (.A1(W13076), .A2(W30912), .ZN(O6067));
  NOR2X1 G6140 (.A1(I1802), .A2(W1731), .ZN(O5933));
  NOR2X1 G6141 (.A1(W16106), .A2(W4004), .ZN(W18813));
  NOR2X1 G6142 (.A1(I1977), .A2(W15194), .ZN(O1652));
  NOR2X1 G6143 (.A1(W30533), .A2(W31980), .ZN(W32041));
  NOR2X1 G6144 (.A1(W21324), .A2(W29442), .ZN(O6244));
  NOR2X1 G6145 (.A1(W28641), .A2(W15892), .ZN(W32043));
  NOR2X1 G6146 (.A1(W4009), .A2(W7338), .ZN(W18808));
  NOR2X1 G6147 (.A1(W9286), .A2(W7387), .ZN(W18807));
  NOR2X1 G6148 (.A1(W6090), .A2(W17771), .ZN(W18806));
  NOR2X1 G6149 (.A1(W4743), .A2(W14730), .ZN(W18805));
  NOR2X1 G6150 (.A1(W26039), .A2(W13385), .ZN(O6069));
  NOR2X1 G6151 (.A1(W19969), .A2(W2177), .ZN(W32047));
  NOR2X1 G6152 (.A1(W8365), .A2(W9498), .ZN(W32892));
  NOR2X1 G6153 (.A1(I697), .A2(W16993), .ZN(W17983));
  NOR2X1 G6154 (.A1(W5650), .A2(W2745), .ZN(W17981));
  NOR2X1 G6155 (.A1(W1036), .A2(W8553), .ZN(W17979));
  NOR2X1 G6156 (.A1(W14101), .A2(W9216), .ZN(W17978));
  NOR2X1 G6157 (.A1(W12667), .A2(W2361), .ZN(W17977));
  NOR2X1 G6158 (.A1(I240), .A2(W16158), .ZN(O1753));
  NOR2X1 G6159 (.A1(W6513), .A2(W16114), .ZN(W17975));
  NOR2X1 G6160 (.A1(W18442), .A2(W11510), .ZN(W19360));
  NOR2X1 G6161 (.A1(W5718), .A2(I995), .ZN(O5801));
  NOR2X1 G6162 (.A1(W24411), .A2(W28061), .ZN(W32893));
  NOR2X1 G6163 (.A1(W3342), .A2(W1108), .ZN(W19361));
  NOR2X1 G6164 (.A1(W13777), .A2(W15696), .ZN(W17970));
  NOR2X1 G6165 (.A1(W6700), .A2(W6321), .ZN(O6450));
  NOR2X1 G6166 (.A1(W7068), .A2(W13187), .ZN(W17968));
  NOR2X1 G6167 (.A1(W1135), .A2(W658), .ZN(W31463));
  NOR2X1 G6168 (.A1(W6526), .A2(W7029), .ZN(W17966));
  NOR2X1 G6169 (.A1(W30129), .A2(W3570), .ZN(W31461));
  NOR2X1 G6170 (.A1(W8109), .A2(W11719), .ZN(W17993));
  NOR2X1 G6171 (.A1(W7965), .A2(W4628), .ZN(W18003));
  NOR2X1 G6172 (.A1(W15805), .A2(W15580), .ZN(W19348));
  NOR2X1 G6173 (.A1(W10836), .A2(W11518), .ZN(W19349));
  NOR2X1 G6174 (.A1(W5430), .A2(I532), .ZN(W17999));
  NOR2X1 G6175 (.A1(W11424), .A2(I905), .ZN(O1480));
  NOR2X1 G6176 (.A1(W9936), .A2(W12061), .ZN(W31472));
  NOR2X1 G6177 (.A1(W3686), .A2(W23438), .ZN(O6441));
  NOR2X1 G6178 (.A1(W1771), .A2(W6898), .ZN(W17994));
  NOR2X1 G6179 (.A1(W10973), .A2(W1944), .ZN(W17963));
  NOR2X1 G6180 (.A1(W15996), .A2(W5076), .ZN(W17991));
  NOR2X1 G6181 (.A1(W4683), .A2(W5755), .ZN(W17990));
  NOR2X1 G6182 (.A1(W5848), .A2(W21089), .ZN(O5803));
  NOR2X1 G6183 (.A1(W3126), .A2(W13807), .ZN(W32879));
  NOR2X1 G6184 (.A1(W13435), .A2(W27391), .ZN(O6444));
  NOR2X1 G6185 (.A1(W7537), .A2(W9548), .ZN(W19355));
  NOR2X1 G6186 (.A1(W24035), .A2(W20000), .ZN(O6445));
  NOR2X1 G6187 (.A1(W9202), .A2(W20577), .ZN(W32929));
  NOR2X1 G6188 (.A1(W2069), .A2(W11511), .ZN(W17942));
  NOR2X1 G6189 (.A1(W16306), .A2(W16379), .ZN(O1472));
  NOR2X1 G6190 (.A1(W17833), .A2(W326), .ZN(W17940));
  NOR2X1 G6191 (.A1(W824), .A2(W24080), .ZN(W32922));
  NOR2X1 G6192 (.A1(W8369), .A2(W28680), .ZN(O6457));
  NOR2X1 G6193 (.A1(W6221), .A2(I550), .ZN(O1471));
  NOR2X1 G6194 (.A1(W21539), .A2(W17343), .ZN(O6458));
  NOR2X1 G6195 (.A1(W11417), .A2(W15216), .ZN(W32927));
  NOR2X1 G6196 (.A1(W19274), .A2(W3206), .ZN(W32915));
  NOR2X1 G6197 (.A1(W6119), .A2(W1950), .ZN(O6460));
  NOR2X1 G6198 (.A1(I1562), .A2(W19230), .ZN(O1758));
  NOR2X1 G6199 (.A1(W2805), .A2(W6441), .ZN(W19373));
  NOR2X1 G6200 (.A1(W12236), .A2(W9037), .ZN(W17929));
  NOR2X1 G6201 (.A1(I166), .A2(W14858), .ZN(W32939));
  NOR2X1 G6202 (.A1(W8743), .A2(W2462), .ZN(W17925));
  NOR2X1 G6203 (.A1(W6341), .A2(W411), .ZN(W17924));
  NOR2X1 G6204 (.A1(W12849), .A2(W4036), .ZN(O6465));
  NOR2X1 G6205 (.A1(W18941), .A2(W16735), .ZN(O1756));
  NOR2X1 G6206 (.A1(W5942), .A2(W6551), .ZN(W17962));
  NOR2X1 G6207 (.A1(W13858), .A2(W1624), .ZN(W17961));
  NOR2X1 G6208 (.A1(W16895), .A2(W28990), .ZN(W32901));
  NOR2X1 G6209 (.A1(W22955), .A2(W28250), .ZN(O5799));
  NOR2X1 G6210 (.A1(W13244), .A2(W13845), .ZN(W17958));
  NOR2X1 G6211 (.A1(W2125), .A2(W9462), .ZN(W17957));
  NOR2X1 G6212 (.A1(W10148), .A2(W3275), .ZN(W17956));
  NOR2X1 G6213 (.A1(W4602), .A2(I1822), .ZN(W19368));
  NOR2X1 G6214 (.A1(W18407), .A2(W12490), .ZN(W32867));
  NOR2X1 G6215 (.A1(W17211), .A2(W15723), .ZN(W17951));
  NOR2X1 G6216 (.A1(W11719), .A2(W21395), .ZN(O6453));
  NOR2X1 G6217 (.A1(W16502), .A2(W13926), .ZN(O1475));
  NOR2X1 G6218 (.A1(W8755), .A2(I1126), .ZN(W17947));
  NOR2X1 G6219 (.A1(W8494), .A2(W2096), .ZN(W32910));
  NOR2X1 G6220 (.A1(W2052), .A2(W21829), .ZN(W32911));
  NOR2X1 G6221 (.A1(W10400), .A2(W4863), .ZN(W17944));
  NOR2X1 G6222 (.A1(W29485), .A2(W13081), .ZN(O6411));
  NOR2X1 G6223 (.A1(W2999), .A2(W18735), .ZN(O5812));
  NOR2X1 G6224 (.A1(W1678), .A2(W14079), .ZN(W18060));
  NOR2X1 G6225 (.A1(W14380), .A2(W1903), .ZN(O1493));
  NOR2X1 G6226 (.A1(W17183), .A2(W17950), .ZN(O1492));
  NOR2X1 G6227 (.A1(W12960), .A2(W13364), .ZN(O1491));
  NOR2X1 G6228 (.A1(W2067), .A2(I1964), .ZN(W18054));
  NOR2X1 G6229 (.A1(W26351), .A2(W342), .ZN(O5808));
  NOR2X1 G6230 (.A1(W29504), .A2(W17762), .ZN(W32817));
  NOR2X1 G6231 (.A1(W17261), .A2(W31036), .ZN(O5814));
  NOR2X1 G6232 (.A1(W8000), .A2(W30014), .ZN(O5807));
  NOR2X1 G6233 (.A1(W13282), .A2(W5710), .ZN(O5806));
  NOR2X1 G6234 (.A1(W9204), .A2(W8115), .ZN(W19335));
  NOR2X1 G6235 (.A1(W6948), .A2(W25540), .ZN(W32830));
  NOR2X1 G6236 (.A1(W13589), .A2(W9181), .ZN(W18045));
  NOR2X1 G6237 (.A1(W7155), .A2(W14073), .ZN(O6420));
  NOR2X1 G6238 (.A1(W1677), .A2(I450), .ZN(O6421));
  NOR2X1 G6239 (.A1(W7472), .A2(W17183), .ZN(W18041));
  NOR2X1 G6240 (.A1(W4409), .A2(W2421), .ZN(W18071));
  NOR2X1 G6241 (.A1(W18810), .A2(W2974), .ZN(O6394));
  NOR2X1 G6242 (.A1(W785), .A2(W3313), .ZN(W18078));
  NOR2X1 G6243 (.A1(W1019), .A2(W6917), .ZN(O5815));
  NOR2X1 G6244 (.A1(W4827), .A2(W7220), .ZN(W32790));
  NOR2X1 G6245 (.A1(W2875), .A2(W30733), .ZN(W32791));
  NOR2X1 G6246 (.A1(W24067), .A2(W9883), .ZN(O6396));
  NOR2X1 G6247 (.A1(W4849), .A2(W8811), .ZN(W19324));
  NOR2X1 G6248 (.A1(W823), .A2(W14542), .ZN(O6398));
  NOR2X1 G6249 (.A1(W16501), .A2(I1280), .ZN(W18040));
  NOR2X1 G6250 (.A1(W24711), .A2(W24276), .ZN(O6399));
  NOR2X1 G6251 (.A1(W22163), .A2(W11883), .ZN(W31500));
  NOR2X1 G6252 (.A1(W6640), .A2(I917), .ZN(W18068));
  NOR2X1 G6253 (.A1(W449), .A2(W14573), .ZN(O1495));
  NOR2X1 G6254 (.A1(W15130), .A2(W14861), .ZN(O1494));
  NOR2X1 G6255 (.A1(W114), .A2(W20780), .ZN(O6404));
  NOR2X1 G6256 (.A1(W4427), .A2(W4870), .ZN(O6405));
  NOR2X1 G6257 (.A1(W22586), .A2(W21803), .ZN(W32860));
  NOR2X1 G6258 (.A1(W18327), .A2(W23678), .ZN(O6429));
  NOR2X1 G6259 (.A1(W22327), .A2(W14767), .ZN(W31475));
  NOR2X1 G6260 (.A1(W30580), .A2(W7566), .ZN(O6431));
  NOR2X1 G6261 (.A1(W5126), .A2(W5449), .ZN(W18019));
  NOR2X1 G6262 (.A1(W18806), .A2(W7327), .ZN(W19342));
  NOR2X1 G6263 (.A1(W7715), .A2(W13827), .ZN(W18017));
  NOR2X1 G6264 (.A1(W19587), .A2(W23036), .ZN(O6435));
  NOR2X1 G6265 (.A1(W19951), .A2(W15085), .ZN(W32858));
  NOR2X1 G6266 (.A1(W11038), .A2(W14127), .ZN(W18023));
  NOR2X1 G6267 (.A1(W9023), .A2(W254), .ZN(O1485));
  NOR2X1 G6268 (.A1(W8472), .A2(W13021), .ZN(W19344));
  NOR2X1 G6269 (.A1(W8156), .A2(W6601), .ZN(W19345));
  NOR2X1 G6270 (.A1(W12268), .A2(W9220), .ZN(W19346));
  NOR2X1 G6271 (.A1(W5532), .A2(W8851), .ZN(W19347));
  NOR2X1 G6272 (.A1(W24225), .A2(W18747), .ZN(O6436));
  NOR2X1 G6273 (.A1(W14135), .A2(W232), .ZN(O1482));
  NOR2X1 G6274 (.A1(W27044), .A2(W17410), .ZN(W32866));
  NOR2X1 G6275 (.A1(W24729), .A2(W30930), .ZN(W31479));
  NOR2X1 G6276 (.A1(W4465), .A2(W2540), .ZN(O6422));
  NOR2X1 G6277 (.A1(W10277), .A2(I906), .ZN(W18038));
  NOR2X1 G6278 (.A1(W32749), .A2(W12530), .ZN(O6423));
  NOR2X1 G6279 (.A1(W8644), .A2(W2522), .ZN(W18036));
  NOR2X1 G6280 (.A1(W24538), .A2(W8348), .ZN(W31480));
  NOR2X1 G6281 (.A1(I227), .A2(W975), .ZN(O6424));
  NOR2X1 G6282 (.A1(W8929), .A2(W28683), .ZN(W32839));
  NOR2X1 G6283 (.A1(W15621), .A2(I1926), .ZN(W18032));
  NOR2X1 G6284 (.A1(W19133), .A2(W12856), .ZN(W19378));
  NOR2X1 G6285 (.A1(W15104), .A2(W1603), .ZN(W18030));
  NOR2X1 G6286 (.A1(W13942), .A2(I1667), .ZN(O6426));
  NOR2X1 G6287 (.A1(W10099), .A2(W3964), .ZN(W31478));
  NOR2X1 G6288 (.A1(W16716), .A2(W16056), .ZN(W18027));
  NOR2X1 G6289 (.A1(W4359), .A2(W11478), .ZN(W32846));
  NOR2X1 G6290 (.A1(W13420), .A2(W7393), .ZN(W19340));
  NOR2X1 G6291 (.A1(I1084), .A2(W909), .ZN(W18024));
  NOR2X1 G6292 (.A1(W6668), .A2(W13044), .ZN(W17809));
  NOR2X1 G6293 (.A1(W14964), .A2(W7796), .ZN(W17820));
  NOR2X1 G6294 (.A1(W21389), .A2(W1796), .ZN(O6523));
  NOR2X1 G6295 (.A1(W2261), .A2(W7577), .ZN(W17816));
  NOR2X1 G6296 (.A1(W8642), .A2(W431), .ZN(O1450));
  NOR2X1 G6297 (.A1(W11827), .A2(W30725), .ZN(W33061));
  NOR2X1 G6298 (.A1(W10140), .A2(W14439), .ZN(W17812));
  NOR2X1 G6299 (.A1(W11662), .A2(W12484), .ZN(W17811));
  NOR2X1 G6300 (.A1(I640), .A2(W16281), .ZN(W33066));
  NOR2X1 G6301 (.A1(W9300), .A2(W2386), .ZN(W17822));
  NOR2X1 G6302 (.A1(W8327), .A2(W1858), .ZN(W17808));
  NOR2X1 G6303 (.A1(W27025), .A2(W3976), .ZN(W33068));
  NOR2X1 G6304 (.A1(W29947), .A2(W14430), .ZN(W33069));
  NOR2X1 G6305 (.A1(W10707), .A2(W14946), .ZN(O1448));
  NOR2X1 G6306 (.A1(W15707), .A2(W30851), .ZN(O5773));
  NOR2X1 G6307 (.A1(W9679), .A2(W1190), .ZN(O5772));
  NOR2X1 G6308 (.A1(W6871), .A2(W6641), .ZN(W17802));
  NOR2X1 G6309 (.A1(W18249), .A2(W26628), .ZN(O5771));
  NOR2X1 G6310 (.A1(W1139), .A2(W3689), .ZN(W33042));
  NOR2X1 G6311 (.A1(I1490), .A2(W10416), .ZN(W17842));
  NOR2X1 G6312 (.A1(W23469), .A2(W29861), .ZN(W31424));
  NOR2X1 G6313 (.A1(W12283), .A2(W14846), .ZN(W19409));
  NOR2X1 G6314 (.A1(W5660), .A2(W14918), .ZN(W17839));
  NOR2X1 G6315 (.A1(W8707), .A2(W12434), .ZN(W17838));
  NOR2X1 G6316 (.A1(W32032), .A2(W11641), .ZN(W33039));
  NOR2X1 G6317 (.A1(W9091), .A2(W15437), .ZN(W19411));
  NOR2X1 G6318 (.A1(W27425), .A2(W10119), .ZN(W33041));
  NOR2X1 G6319 (.A1(W1052), .A2(W8440), .ZN(W17800));
  NOR2X1 G6320 (.A1(W25663), .A2(W12483), .ZN(O6516));
  NOR2X1 G6321 (.A1(W4615), .A2(W4213), .ZN(W33048));
  NOR2X1 G6322 (.A1(W15467), .A2(I170), .ZN(W17828));
  NOR2X1 G6323 (.A1(W9032), .A2(W8663), .ZN(W17827));
  NOR2X1 G6324 (.A1(W31885), .A2(W21176), .ZN(W33051));
  NOR2X1 G6325 (.A1(W17239), .A2(I410), .ZN(W17825));
  NOR2X1 G6326 (.A1(W7214), .A2(W4951), .ZN(O1452));
  NOR2X1 G6327 (.A1(W13398), .A2(W1031), .ZN(W17772));
  NOR2X1 G6328 (.A1(W7021), .A2(W9164), .ZN(O6537));
  NOR2X1 G6329 (.A1(W5463), .A2(I266), .ZN(O6538));
  NOR2X1 G6330 (.A1(W2569), .A2(I1235), .ZN(W17779));
  NOR2X1 G6331 (.A1(W1479), .A2(W8205), .ZN(W17778));
  NOR2X1 G6332 (.A1(W6235), .A2(W17547), .ZN(W19426));
  NOR2X1 G6333 (.A1(W23996), .A2(W590), .ZN(O6539));
  NOR2X1 G6334 (.A1(W10325), .A2(W4251), .ZN(W19427));
  NOR2X1 G6335 (.A1(W11432), .A2(W3327), .ZN(W33097));
  NOR2X1 G6336 (.A1(W22715), .A2(W2644), .ZN(W33087));
  NOR2X1 G6337 (.A1(W8490), .A2(W6110), .ZN(W17771));
  NOR2X1 G6338 (.A1(W4433), .A2(W2494), .ZN(O1773));
  NOR2X1 G6339 (.A1(W6198), .A2(W900), .ZN(W33104));
  NOR2X1 G6340 (.A1(W6404), .A2(W10746), .ZN(W17767));
  NOR2X1 G6341 (.A1(W12082), .A2(W4367), .ZN(O6543));
  NOR2X1 G6342 (.A1(W15446), .A2(W5180), .ZN(W19431));
  NOR2X1 G6343 (.A1(W11925), .A2(W21907), .ZN(W33110));
  NOR2X1 G6344 (.A1(I700), .A2(I1540), .ZN(W17762));
  NOR2X1 G6345 (.A1(W11604), .A2(I1609), .ZN(W17790));
  NOR2X1 G6346 (.A1(W2863), .A2(W31481), .ZN(W33073));
  NOR2X1 G6347 (.A1(W1157), .A2(W3415), .ZN(O6530));
  NOR2X1 G6348 (.A1(I686), .A2(W4438), .ZN(W17797));
  NOR2X1 G6349 (.A1(W14880), .A2(W16049), .ZN(O1446));
  NOR2X1 G6350 (.A1(W8439), .A2(W7766), .ZN(W17795));
  NOR2X1 G6351 (.A1(W7078), .A2(W7076), .ZN(W31404));
  NOR2X1 G6352 (.A1(W2512), .A2(W13962), .ZN(O6531));
  NOR2X1 G6353 (.A1(W4913), .A2(W30131), .ZN(O6532));
  NOR2X1 G6354 (.A1(W4290), .A2(W29540), .ZN(W33029));
  NOR2X1 G6355 (.A1(W363), .A2(W15072), .ZN(W17789));
  NOR2X1 G6356 (.A1(W9613), .A2(W7361), .ZN(W17788));
  NOR2X1 G6357 (.A1(W19433), .A2(W4438), .ZN(W33083));
  NOR2X1 G6358 (.A1(W3265), .A2(W15063), .ZN(W31401));
  NOR2X1 G6359 (.A1(W5000), .A2(W1652), .ZN(W17785));
  NOR2X1 G6360 (.A1(W16909), .A2(W8066), .ZN(W31400));
  NOR2X1 G6361 (.A1(W5542), .A2(I85), .ZN(W17783));
  NOR2X1 G6362 (.A1(W9846), .A2(W9519), .ZN(W17893));
  NOR2X1 G6363 (.A1(W11284), .A2(W2487), .ZN(W17902));
  NOR2X1 G6364 (.A1(W10986), .A2(I679), .ZN(W19384));
  NOR2X1 G6365 (.A1(I724), .A2(W9024), .ZN(W17899));
  NOR2X1 G6366 (.A1(W1820), .A2(W3894), .ZN(W17898));
  NOR2X1 G6367 (.A1(I544), .A2(W14246), .ZN(O5791));
  NOR2X1 G6368 (.A1(W2774), .A2(W2373), .ZN(W17896));
  NOR2X1 G6369 (.A1(W2079), .A2(W25110), .ZN(W31444));
  NOR2X1 G6370 (.A1(W10677), .A2(I488), .ZN(W17894));
  NOR2X1 G6371 (.A1(I386), .A2(W14857), .ZN(W32967));
  NOR2X1 G6372 (.A1(W7135), .A2(W7609), .ZN(W19387));
  NOR2X1 G6373 (.A1(W5131), .A2(W2386), .ZN(O1761));
  NOR2X1 G6374 (.A1(W22614), .A2(W14262), .ZN(W31443));
  NOR2X1 G6375 (.A1(W19810), .A2(I1252), .ZN(W32980));
  NOR2X1 G6376 (.A1(W11958), .A2(W1267), .ZN(O1464));
  NOR2X1 G6377 (.A1(W15372), .A2(W7807), .ZN(O1463));
  NOR2X1 G6378 (.A1(W5278), .A2(I1473), .ZN(W19390));
  NOR2X1 G6379 (.A1(W792), .A2(W12342), .ZN(W17885));
  NOR2X1 G6380 (.A1(W7905), .A2(W3109), .ZN(W19381));
  NOR2X1 G6381 (.A1(W30309), .A2(W15341), .ZN(W31449));
  NOR2X1 G6382 (.A1(W17259), .A2(W9680), .ZN(W17918));
  NOR2X1 G6383 (.A1(W29732), .A2(W32808), .ZN(W32948));
  NOR2X1 G6384 (.A1(W15809), .A2(W14738), .ZN(W19380));
  NOR2X1 G6385 (.A1(W12140), .A2(I1675), .ZN(O6469));
  NOR2X1 G6386 (.A1(W17637), .A2(W23531), .ZN(O6471));
  NOR2X1 G6387 (.A1(W4699), .A2(W10837), .ZN(W32955));
  NOR2X1 G6388 (.A1(W19955), .A2(W15085), .ZN(O6473));
  NOR2X1 G6389 (.A1(W15731), .A2(W9535), .ZN(O1462));
  NOR2X1 G6390 (.A1(W12692), .A2(W15838), .ZN(W17910));
  NOR2X1 G6391 (.A1(W11764), .A2(W29200), .ZN(W32960));
  NOR2X1 G6392 (.A1(W13273), .A2(W4710), .ZN(O1759));
  NOR2X1 G6393 (.A1(W109), .A2(W3835), .ZN(W17907));
  NOR2X1 G6394 (.A1(W17142), .A2(W1117), .ZN(W17906));
  NOR2X1 G6395 (.A1(I854), .A2(W22123), .ZN(W32962));
  NOR2X1 G6396 (.A1(W2811), .A2(W7603), .ZN(O6476));
  NOR2X1 G6397 (.A1(W16624), .A2(W11112), .ZN(W19402));
  NOR2X1 G6398 (.A1(W5571), .A2(W8757), .ZN(W17864));
  NOR2X1 G6399 (.A1(W6835), .A2(W856), .ZN(O1456));
  NOR2X1 G6400 (.A1(W3346), .A2(W1822), .ZN(W17860));
  NOR2X1 G6401 (.A1(W5635), .A2(W21872), .ZN(W33006));
  NOR2X1 G6402 (.A1(W16407), .A2(W5466), .ZN(W17858));
  NOR2X1 G6403 (.A1(I1758), .A2(W5971), .ZN(W31431));
  NOR2X1 G6404 (.A1(W30273), .A2(I1310), .ZN(O6503));
  NOR2X1 G6405 (.A1(W17554), .A2(W13475), .ZN(O6505));
  NOR2X1 G6406 (.A1(W11270), .A2(W22186), .ZN(O6498));
  NOR2X1 G6407 (.A1(W11542), .A2(W19013), .ZN(O5785));
  NOR2X1 G6408 (.A1(W12696), .A2(I1314), .ZN(W17851));
  NOR2X1 G6409 (.A1(W19260), .A2(W23740), .ZN(O5784));
  NOR2X1 G6410 (.A1(W8474), .A2(W7420), .ZN(O6508));
  NOR2X1 G6411 (.A1(W30684), .A2(W1969), .ZN(W33022));
  NOR2X1 G6412 (.A1(W12770), .A2(W6292), .ZN(W19405));
  NOR2X1 G6413 (.A1(W27185), .A2(W7693), .ZN(W33026));
  NOR2X1 G6414 (.A1(W3048), .A2(W9788), .ZN(W31426));
  NOR2X1 G6415 (.A1(W11311), .A2(W10392), .ZN(W17874));
  NOR2X1 G6416 (.A1(W17405), .A2(W18028), .ZN(O6488));
  NOR2X1 G6417 (.A1(W30083), .A2(W16529), .ZN(W31440));
  NOR2X1 G6418 (.A1(W15357), .A2(W2599), .ZN(W17880));
  NOR2X1 G6419 (.A1(W24259), .A2(W1987), .ZN(O6490));
  NOR2X1 G6420 (.A1(W25376), .A2(W26976), .ZN(O6491));
  NOR2X1 G6421 (.A1(W23595), .A2(I1850), .ZN(W31439));
  NOR2X1 G6422 (.A1(I268), .A2(W14640), .ZN(W17876));
  NOR2X1 G6423 (.A1(W7782), .A2(W11389), .ZN(W17875));
  NOR2X1 G6424 (.A1(W259), .A2(I1659), .ZN(O6392));
  NOR2X1 G6425 (.A1(W502), .A2(W622), .ZN(W19394));
  NOR2X1 G6426 (.A1(W6557), .A2(W15637), .ZN(W32993));
  NOR2X1 G6427 (.A1(W27882), .A2(W20301), .ZN(O5789));
  NOR2X1 G6428 (.A1(I1253), .A2(W531), .ZN(W19396));
  NOR2X1 G6429 (.A1(W18031), .A2(W18228), .ZN(O6495));
  NOR2X1 G6430 (.A1(W14244), .A2(W6264), .ZN(O1457));
  NOR2X1 G6431 (.A1(W25179), .A2(W10481), .ZN(O6497));
  NOR2X1 G6432 (.A1(W710), .A2(I885), .ZN(W18281));
  NOR2X1 G6433 (.A1(W28827), .A2(W11764), .ZN(W32562));
  NOR2X1 G6434 (.A1(W14819), .A2(W13665), .ZN(O1734));
  NOR2X1 G6435 (.A1(W18709), .A2(W14451), .ZN(W19253));
  NOR2X1 G6436 (.A1(W2350), .A2(W9745), .ZN(O1735));
  NOR2X1 G6437 (.A1(W17696), .A2(W7585), .ZN(O6294));
  NOR2X1 G6438 (.A1(W40), .A2(W7954), .ZN(W31568));
  NOR2X1 G6439 (.A1(I1943), .A2(W10715), .ZN(W18283));
  NOR2X1 G6440 (.A1(I1059), .A2(W2514), .ZN(O6295));
  NOR2X1 G6441 (.A1(W3036), .A2(W10921), .ZN(W18292));
  NOR2X1 G6442 (.A1(W21749), .A2(W30216), .ZN(W32572));
  NOR2X1 G6443 (.A1(W18050), .A2(W6032), .ZN(W32573));
  NOR2X1 G6444 (.A1(W8145), .A2(W4084), .ZN(W19258));
  NOR2X1 G6445 (.A1(W5243), .A2(W3117), .ZN(W19259));
  NOR2X1 G6446 (.A1(W28884), .A2(W11475), .ZN(W32578));
  NOR2X1 G6447 (.A1(W15707), .A2(I81), .ZN(W32580));
  NOR2X1 G6448 (.A1(W2910), .A2(W29641), .ZN(W32581));
  NOR2X1 G6449 (.A1(W5428), .A2(W9250), .ZN(W18273));
  NOR2X1 G6450 (.A1(W2868), .A2(W3300), .ZN(O6285));
  NOR2X1 G6451 (.A1(W25231), .A2(W24553), .ZN(O5847));
  NOR2X1 G6452 (.A1(W29809), .A2(W26575), .ZN(W32543));
  NOR2X1 G6453 (.A1(W14052), .A2(W9914), .ZN(W18306));
  NOR2X1 G6454 (.A1(W16079), .A2(W6129), .ZN(O6279));
  NOR2X1 G6455 (.A1(W22518), .A2(W27012), .ZN(W32546));
  NOR2X1 G6456 (.A1(W727), .A2(W4372), .ZN(W31581));
  NOR2X1 G6457 (.A1(W2202), .A2(W2757), .ZN(W18302));
  NOR2X1 G6458 (.A1(W6157), .A2(W4803), .ZN(W31580));
  NOR2X1 G6459 (.A1(W9712), .A2(W9086), .ZN(W18272));
  NOR2X1 G6460 (.A1(W13333), .A2(W3245), .ZN(W19250));
  NOR2X1 G6461 (.A1(W8353), .A2(W19697), .ZN(O6287));
  NOR2X1 G6462 (.A1(W4178), .A2(W3578), .ZN(O5846));
  NOR2X1 G6463 (.A1(W10650), .A2(W7310), .ZN(W18296));
  NOR2X1 G6464 (.A1(W420), .A2(W2614), .ZN(W18295));
  NOR2X1 G6465 (.A1(W3615), .A2(W23551), .ZN(O6289));
  NOR2X1 G6466 (.A1(W29074), .A2(W32149), .ZN(W32560));
  NOR2X1 G6467 (.A1(I1955), .A2(W4366), .ZN(O1525));
  NOR2X1 G6468 (.A1(I337), .A2(W3314), .ZN(O1527));
  NOR2X1 G6469 (.A1(W19775), .A2(W18508), .ZN(O5839));
  NOR2X1 G6470 (.A1(W18020), .A2(W18295), .ZN(O6309));
  NOR2X1 G6471 (.A1(W3768), .A2(W8284), .ZN(W18247));
  NOR2X1 G6472 (.A1(W1189), .A2(W3814), .ZN(W18246));
  NOR2X1 G6473 (.A1(W5314), .A2(W17987), .ZN(W18245));
  NOR2X1 G6474 (.A1(W29066), .A2(I235), .ZN(W31554));
  NOR2X1 G6475 (.A1(W4045), .A2(W1754), .ZN(W19266));
  NOR2X1 G6476 (.A1(W288), .A2(W16461), .ZN(W18252));
  NOR2X1 G6477 (.A1(W20697), .A2(I219), .ZN(W32615));
  NOR2X1 G6478 (.A1(W11318), .A2(W10045), .ZN(O1524));
  NOR2X1 G6479 (.A1(W1791), .A2(W9725), .ZN(O5836));
  NOR2X1 G6480 (.A1(W1339), .A2(W13122), .ZN(W18237));
  NOR2X1 G6481 (.A1(W8119), .A2(W18042), .ZN(W18236));
  NOR2X1 G6482 (.A1(W22857), .A2(W28148), .ZN(W31550));
  NOR2X1 G6483 (.A1(W17392), .A2(W5987), .ZN(W32619));
  NOR2X1 G6484 (.A1(W5053), .A2(W19116), .ZN(O6317));
  NOR2X1 G6485 (.A1(W14059), .A2(W18465), .ZN(O6304));
  NOR2X1 G6486 (.A1(W19973), .A2(W29562), .ZN(W32582));
  NOR2X1 G6487 (.A1(W10445), .A2(W12607), .ZN(W32583));
  NOR2X1 G6488 (.A1(W7597), .A2(W1988), .ZN(O1533));
  NOR2X1 G6489 (.A1(W9867), .A2(I1931), .ZN(O6303));
  NOR2X1 G6490 (.A1(W17754), .A2(W3781), .ZN(W32593));
  NOR2X1 G6491 (.A1(W2894), .A2(W9494), .ZN(O1530));
  NOR2X1 G6492 (.A1(W14620), .A2(W13383), .ZN(W18264));
  NOR2X1 G6493 (.A1(W10533), .A2(W15060), .ZN(W18263));
  NOR2X1 G6494 (.A1(W15102), .A2(W8436), .ZN(W19244));
  NOR2X1 G6495 (.A1(W963), .A2(W29694), .ZN(O6305));
  NOR2X1 G6496 (.A1(I42), .A2(W25228), .ZN(W32597));
  NOR2X1 G6497 (.A1(W2071), .A2(W12591), .ZN(W32598));
  NOR2X1 G6498 (.A1(W7302), .A2(W7640), .ZN(W18256));
  NOR2X1 G6499 (.A1(W32498), .A2(W1168), .ZN(O6306));
  NOR2X1 G6500 (.A1(W2751), .A2(W28522), .ZN(O6307));
  NOR2X1 G6501 (.A1(W10707), .A2(W7436), .ZN(O6308));
  NOR2X1 G6502 (.A1(W3001), .A2(W26988), .ZN(W32493));
  NOR2X1 G6503 (.A1(W10346), .A2(I1724), .ZN(W32483));
  NOR2X1 G6504 (.A1(W13887), .A2(W13450), .ZN(W18368));
  NOR2X1 G6505 (.A1(W26306), .A2(W30775), .ZN(O6251));
  NOR2X1 G6506 (.A1(W27642), .A2(W22134), .ZN(W31608));
  NOR2X1 G6507 (.A1(W20115), .A2(W15198), .ZN(O5859));
  NOR2X1 G6508 (.A1(W12), .A2(W587), .ZN(W18364));
  NOR2X1 G6509 (.A1(W12809), .A2(W16695), .ZN(O1557));
  NOR2X1 G6510 (.A1(W633), .A2(W24009), .ZN(O6255));
  NOR2X1 G6511 (.A1(W30166), .A2(W15), .ZN(O5860));
  NOR2X1 G6512 (.A1(W16135), .A2(W1175), .ZN(W18359));
  NOR2X1 G6513 (.A1(W10229), .A2(W1227), .ZN(W18358));
  NOR2X1 G6514 (.A1(W30078), .A2(W5929), .ZN(O6256));
  NOR2X1 G6515 (.A1(W7081), .A2(I1337), .ZN(W18356));
  NOR2X1 G6516 (.A1(W11795), .A2(W25631), .ZN(W32497));
  NOR2X1 G6517 (.A1(W5469), .A2(W18929), .ZN(W19229));
  NOR2X1 G6518 (.A1(W4645), .A2(W10147), .ZN(W18353));
  NOR2X1 G6519 (.A1(W29397), .A2(W29125), .ZN(W32500));
  NOR2X1 G6520 (.A1(W10202), .A2(W21257), .ZN(O6247));
  NOR2X1 G6521 (.A1(W1818), .A2(W25457), .ZN(O6245));
  NOR2X1 G6522 (.A1(I915), .A2(W3008), .ZN(W18386));
  NOR2X1 G6523 (.A1(W4322), .A2(I1107), .ZN(W32467));
  NOR2X1 G6524 (.A1(W5706), .A2(W11665), .ZN(W32469));
  NOR2X1 G6525 (.A1(W2644), .A2(W1051), .ZN(W32470));
  NOR2X1 G6526 (.A1(W2667), .A2(W14414), .ZN(W18382));
  NOR2X1 G6527 (.A1(W3506), .A2(W1081), .ZN(O6246));
  NOR2X1 G6528 (.A1(W11456), .A2(W22022), .ZN(W31614));
  NOR2X1 G6529 (.A1(W20031), .A2(W26115), .ZN(W32501));
  NOR2X1 G6530 (.A1(W13495), .A2(W11487), .ZN(W18378));
  NOR2X1 G6531 (.A1(W13247), .A2(W24126), .ZN(W31612));
  NOR2X1 G6532 (.A1(W2503), .A2(W9359), .ZN(W18375));
  NOR2X1 G6533 (.A1(W1616), .A2(W3259), .ZN(W18374));
  NOR2X1 G6534 (.A1(W14984), .A2(W3337), .ZN(W18373));
  NOR2X1 G6535 (.A1(W2375), .A2(W17771), .ZN(W19224));
  NOR2X1 G6536 (.A1(W29847), .A2(W19500), .ZN(W32481));
  NOR2X1 G6537 (.A1(W4451), .A2(W14184), .ZN(W18322));
  NOR2X1 G6538 (.A1(W17827), .A2(I1113), .ZN(W18330));
  NOR2X1 G6539 (.A1(W4760), .A2(W18727), .ZN(W31599));
  NOR2X1 G6540 (.A1(W13988), .A2(W13387), .ZN(W18328));
  NOR2X1 G6541 (.A1(W2635), .A2(W24345), .ZN(O6271));
  NOR2X1 G6542 (.A1(W13917), .A2(W6422), .ZN(W32525));
  NOR2X1 G6543 (.A1(W11546), .A2(W14979), .ZN(W18325));
  NOR2X1 G6544 (.A1(W14593), .A2(W11583), .ZN(O1546));
  NOR2X1 G6545 (.A1(W1992), .A2(W29928), .ZN(W32526));
  NOR2X1 G6546 (.A1(W16854), .A2(W4667), .ZN(O1547));
  NOR2X1 G6547 (.A1(W784), .A2(W3969), .ZN(W32527));
  NOR2X1 G6548 (.A1(W8552), .A2(W4089), .ZN(W32528));
  NOR2X1 G6549 (.A1(W5825), .A2(W15935), .ZN(O1731));
  NOR2X1 G6550 (.A1(W12904), .A2(W1556), .ZN(W31597));
  NOR2X1 G6551 (.A1(W2946), .A2(W14523), .ZN(W18316));
  NOR2X1 G6552 (.A1(W6700), .A2(W18258), .ZN(W18315));
  NOR2X1 G6553 (.A1(W11668), .A2(W19596), .ZN(O5852));
  NOR2X1 G6554 (.A1(W16278), .A2(W4307), .ZN(W32537));
  NOR2X1 G6555 (.A1(W24406), .A2(W27161), .ZN(O5856));
  NOR2X1 G6556 (.A1(W19148), .A2(W1345), .ZN(W32504));
  NOR2X1 G6557 (.A1(W1911), .A2(W3470), .ZN(W18348));
  NOR2X1 G6558 (.A1(W7455), .A2(W9480), .ZN(W32505));
  NOR2X1 G6559 (.A1(W2106), .A2(W14208), .ZN(W19231));
  NOR2X1 G6560 (.A1(W24447), .A2(W3608), .ZN(W32507));
  NOR2X1 G6561 (.A1(W10378), .A2(W31335), .ZN(O6260));
  NOR2X1 G6562 (.A1(W14723), .A2(W1802), .ZN(W19232));
  NOR2X1 G6563 (.A1(W22603), .A2(W24132), .ZN(W32511));
  NOR2X1 G6564 (.A1(W27907), .A2(W5943), .ZN(O5834));
  NOR2X1 G6565 (.A1(I902), .A2(W9049), .ZN(W19234));
  NOR2X1 G6566 (.A1(W2277), .A2(W9810), .ZN(W18339));
  NOR2X1 G6567 (.A1(W13334), .A2(W9685), .ZN(W19236));
  NOR2X1 G6568 (.A1(W1182), .A2(W17415), .ZN(W18335));
  NOR2X1 G6569 (.A1(W14707), .A2(W11194), .ZN(W18334));
  NOR2X1 G6570 (.A1(W13028), .A2(W27046), .ZN(O6268));
  NOR2X1 G6571 (.A1(W23361), .A2(W18796), .ZN(O6269));
  NOR2X1 G6572 (.A1(I109), .A2(W7286), .ZN(W19304));
  NOR2X1 G6573 (.A1(W3292), .A2(W11470), .ZN(W31517));
  NOR2X1 G6574 (.A1(W18304), .A2(I1428), .ZN(W19302));
  NOR2X1 G6575 (.A1(W24635), .A2(W32635), .ZN(O6367));
  NOR2X1 G6576 (.A1(W7961), .A2(W12968), .ZN(O5821));
  NOR2X1 G6577 (.A1(W5787), .A2(W14882), .ZN(O1509));
  NOR2X1 G6578 (.A1(W1189), .A2(W1598), .ZN(W32723));
  NOR2X1 G6579 (.A1(W598), .A2(W5956), .ZN(W18129));
  NOR2X1 G6580 (.A1(W3930), .A2(W26505), .ZN(W32724));
  NOR2X1 G6581 (.A1(W7892), .A2(W9818), .ZN(O6366));
  NOR2X1 G6582 (.A1(W3389), .A2(W14809), .ZN(O1507));
  NOR2X1 G6583 (.A1(W16270), .A2(W95), .ZN(O6368));
  NOR2X1 G6584 (.A1(W1325), .A2(W5853), .ZN(O1743));
  NOR2X1 G6585 (.A1(W7067), .A2(W17680), .ZN(W18123));
  NOR2X1 G6586 (.A1(W27130), .A2(W10409), .ZN(W32728));
  NOR2X1 G6587 (.A1(W27704), .A2(W23010), .ZN(O5820));
  NOR2X1 G6588 (.A1(W14722), .A2(W15915), .ZN(O1744));
  NOR2X1 G6589 (.A1(W9577), .A2(W14522), .ZN(W18119));
  NOR2X1 G6590 (.A1(W2662), .A2(W15232), .ZN(W18144));
  NOR2X1 G6591 (.A1(W1718), .A2(W5994), .ZN(W18152));
  NOR2X1 G6592 (.A1(I621), .A2(W12734), .ZN(O6358));
  NOR2X1 G6593 (.A1(W8609), .A2(W10128), .ZN(W18150));
  NOR2X1 G6594 (.A1(W2320), .A2(W8626), .ZN(W18149));
  NOR2X1 G6595 (.A1(W27177), .A2(W7115), .ZN(W32705));
  NOR2X1 G6596 (.A1(W9970), .A2(W16825), .ZN(W19297));
  NOR2X1 G6597 (.A1(W10263), .A2(W16650), .ZN(O1512));
  NOR2X1 G6598 (.A1(W22200), .A2(W10354), .ZN(O6362));
  NOR2X1 G6599 (.A1(W3427), .A2(W4578), .ZN(O6372));
  NOR2X1 G6600 (.A1(W16039), .A2(W13071), .ZN(W18143));
  NOR2X1 G6601 (.A1(W15834), .A2(W1890), .ZN(O1511));
  NOR2X1 G6602 (.A1(W651), .A2(W9154), .ZN(W18141));
  NOR2X1 G6603 (.A1(W10625), .A2(W14079), .ZN(W19298));
  NOR2X1 G6604 (.A1(W11617), .A2(W1028), .ZN(O1510));
  NOR2X1 G6605 (.A1(W8580), .A2(W16394), .ZN(W19299));
  NOR2X1 G6606 (.A1(W10509), .A2(W23129), .ZN(W31518));
  NOR2X1 G6607 (.A1(W16749), .A2(W8748), .ZN(O1745));
  NOR2X1 G6608 (.A1(W16102), .A2(W17241), .ZN(W19312));
  NOR2X1 G6609 (.A1(I501), .A2(W9668), .ZN(W18098));
  NOR2X1 G6610 (.A1(W12629), .A2(W4820), .ZN(W18097));
  NOR2X1 G6611 (.A1(W11859), .A2(W14173), .ZN(O5818));
  NOR2X1 G6612 (.A1(W16826), .A2(W13150), .ZN(O6389));
  NOR2X1 G6613 (.A1(W4995), .A2(W7439), .ZN(W19314));
  NOR2X1 G6614 (.A1(W9481), .A2(W18493), .ZN(W19316));
  NOR2X1 G6615 (.A1(W1269), .A2(W21248), .ZN(W32775));
  NOR2X1 G6616 (.A1(W8480), .A2(W18305), .ZN(W19311));
  NOR2X1 G6617 (.A1(W25345), .A2(W30758), .ZN(W32778));
  NOR2X1 G6618 (.A1(W1196), .A2(W3279), .ZN(W18088));
  NOR2X1 G6619 (.A1(W6597), .A2(W13714), .ZN(W19318));
  NOR2X1 G6620 (.A1(W7977), .A2(W8260), .ZN(O1746));
  NOR2X1 G6621 (.A1(W13091), .A2(W7288), .ZN(W31505));
  NOR2X1 G6622 (.A1(W27538), .A2(W4833), .ZN(W32782));
  NOR2X1 G6623 (.A1(W5675), .A2(W2538), .ZN(O1499));
  NOR2X1 G6624 (.A1(W28785), .A2(W29855), .ZN(O5816));
  NOR2X1 G6625 (.A1(W3746), .A2(W4040), .ZN(W18109));
  NOR2X1 G6626 (.A1(W12265), .A2(I578), .ZN(W32733));
  NOR2X1 G6627 (.A1(W14360), .A2(W13239), .ZN(W31512));
  NOR2X1 G6628 (.A1(W19161), .A2(I668), .ZN(O6379));
  NOR2X1 G6629 (.A1(W15369), .A2(W16010), .ZN(W32745));
  NOR2X1 G6630 (.A1(W16612), .A2(W32006), .ZN(O6381));
  NOR2X1 G6631 (.A1(W13998), .A2(W4121), .ZN(W32751));
  NOR2X1 G6632 (.A1(W2616), .A2(I1507), .ZN(W18111));
  NOR2X1 G6633 (.A1(W8888), .A2(W23205), .ZN(O5819));
  NOR2X1 G6634 (.A1(W18758), .A2(W4731), .ZN(O1742));
  NOR2X1 G6635 (.A1(W19975), .A2(W12356), .ZN(O6383));
  NOR2X1 G6636 (.A1(W8731), .A2(W14221), .ZN(O6384));
  NOR2X1 G6637 (.A1(W17091), .A2(W27171), .ZN(W32760));
  NOR2X1 G6638 (.A1(W26623), .A2(W13552), .ZN(W32763));
  NOR2X1 G6639 (.A1(W12911), .A2(I145), .ZN(W18103));
  NOR2X1 G6640 (.A1(W11561), .A2(W11960), .ZN(W18102));
  NOR2X1 G6641 (.A1(W15823), .A2(W17227), .ZN(W32766));
  NOR2X1 G6642 (.A1(W14465), .A2(I1271), .ZN(W19284));
  NOR2X1 G6643 (.A1(W15962), .A2(W8984), .ZN(O1520));
  NOR2X1 G6644 (.A1(W10877), .A2(W29654), .ZN(O6327));
  NOR2X1 G6645 (.A1(W15890), .A2(I304), .ZN(W18209));
  NOR2X1 G6646 (.A1(W11131), .A2(W8592), .ZN(W18206));
  NOR2X1 G6647 (.A1(W2805), .A2(W8159), .ZN(W31533));
  NOR2X1 G6648 (.A1(I1478), .A2(W18361), .ZN(W19282));
  NOR2X1 G6649 (.A1(W20796), .A2(W11616), .ZN(O5828));
  NOR2X1 G6650 (.A1(W29440), .A2(W16103), .ZN(O6333));
  NOR2X1 G6651 (.A1(W25204), .A2(W31219), .ZN(W32642));
  NOR2X1 G6652 (.A1(W5086), .A2(W736), .ZN(W18200));
  NOR2X1 G6653 (.A1(W10788), .A2(W21664), .ZN(O6334));
  NOR2X1 G6654 (.A1(W19298), .A2(W12645), .ZN(W32658));
  NOR2X1 G6655 (.A1(W31724), .A2(W2658), .ZN(W32659));
  NOR2X1 G6656 (.A1(W2150), .A2(W16559), .ZN(W31531));
  NOR2X1 G6657 (.A1(W12998), .A2(W12715), .ZN(W32661));
  NOR2X1 G6658 (.A1(W21498), .A2(W6127), .ZN(W32662));
  NOR2X1 G6659 (.A1(W23809), .A2(W0), .ZN(O5827));
  NOR2X1 G6660 (.A1(W29841), .A2(W5351), .ZN(O6323));
  NOR2X1 G6661 (.A1(W19329), .A2(W7412), .ZN(W32624));
  NOR2X1 G6662 (.A1(W6221), .A2(W10465), .ZN(W32625));
  NOR2X1 G6663 (.A1(I565), .A2(W9648), .ZN(W18228));
  NOR2X1 G6664 (.A1(W16438), .A2(I1062), .ZN(W18227));
  NOR2X1 G6665 (.A1(W19657), .A2(W29926), .ZN(O6319));
  NOR2X1 G6666 (.A1(W17092), .A2(I1393), .ZN(W18225));
  NOR2X1 G6667 (.A1(W6614), .A2(W16326), .ZN(W19272));
  NOR2X1 G6668 (.A1(W17860), .A2(W16558), .ZN(W32629));
  NOR2X1 G6669 (.A1(W31434), .A2(W32295), .ZN(W32664));
  NOR2X1 G6670 (.A1(W201), .A2(W10031), .ZN(W19274));
  NOR2X1 G6671 (.A1(W4638), .A2(W7447), .ZN(W18219));
  NOR2X1 G6672 (.A1(W9079), .A2(W5616), .ZN(W18218));
  NOR2X1 G6673 (.A1(W10028), .A2(W8772), .ZN(W19275));
  NOR2X1 G6674 (.A1(W38), .A2(W13326), .ZN(W32636));
  NOR2X1 G6675 (.A1(W6239), .A2(W1979), .ZN(W19276));
  NOR2X1 G6676 (.A1(I1748), .A2(W28747), .ZN(O5831));
  NOR2X1 G6677 (.A1(W2898), .A2(W3768), .ZN(W18163));
  NOR2X1 G6678 (.A1(W17587), .A2(W8283), .ZN(W18171));
  NOR2X1 G6679 (.A1(W9441), .A2(W12085), .ZN(W18170));
  NOR2X1 G6680 (.A1(W26634), .A2(W22959), .ZN(O5824));
  NOR2X1 G6681 (.A1(W3097), .A2(W13933), .ZN(W18168));
  NOR2X1 G6682 (.A1(W21961), .A2(W2387), .ZN(W31522));
  NOR2X1 G6683 (.A1(W13056), .A2(W14173), .ZN(W18166));
  NOR2X1 G6684 (.A1(W7924), .A2(I1416), .ZN(W18165));
  NOR2X1 G6685 (.A1(W26063), .A2(W5672), .ZN(O6349));
  NOR2X1 G6686 (.A1(W29289), .A2(W16292), .ZN(W32686));
  NOR2X1 G6687 (.A1(I322), .A2(W2413), .ZN(O1513));
  NOR2X1 G6688 (.A1(W10106), .A2(W12492), .ZN(W18159));
  NOR2X1 G6689 (.A1(W25829), .A2(W31843), .ZN(W32698));
  NOR2X1 G6690 (.A1(W9996), .A2(W13192), .ZN(W18157));
  NOR2X1 G6691 (.A1(W14142), .A2(I1064), .ZN(W19295));
  NOR2X1 G6692 (.A1(W3220), .A2(W13705), .ZN(W18155));
  NOR2X1 G6693 (.A1(W31542), .A2(W4840), .ZN(O6355));
  NOR2X1 G6694 (.A1(W28483), .A2(W529), .ZN(O6340));
  NOR2X1 G6695 (.A1(W3425), .A2(W19069), .ZN(W19287));
  NOR2X1 G6696 (.A1(I14), .A2(W5782), .ZN(O1517));
  NOR2X1 G6697 (.A1(W17430), .A2(W17480), .ZN(W18189));
  NOR2X1 G6698 (.A1(W3623), .A2(W2793), .ZN(W18188));
  NOR2X1 G6699 (.A1(W17774), .A2(W18130), .ZN(W18186));
  NOR2X1 G6700 (.A1(W18118), .A2(W285), .ZN(W32670));
  NOR2X1 G6701 (.A1(W29258), .A2(W26520), .ZN(W32673));
  NOR2X1 G6702 (.A1(W11927), .A2(W30225), .ZN(W32674));
  NOR2X1 G6703 (.A1(W4589), .A2(W14072), .ZN(W16494));
  NOR2X1 G6704 (.A1(W12663), .A2(W266), .ZN(W18180));
  NOR2X1 G6705 (.A1(W31594), .A2(I228), .ZN(O6344));
  NOR2X1 G6706 (.A1(W1697), .A2(I1558), .ZN(O6346));
  NOR2X1 G6707 (.A1(W6621), .A2(W16756), .ZN(W18176));
  NOR2X1 G6708 (.A1(I872), .A2(W12360), .ZN(W18175));
  NOR2X1 G6709 (.A1(W16610), .A2(W31769), .ZN(O6347));
  NOR2X1 G6710 (.A1(I102), .A2(W12643), .ZN(W32685));
  NOR2X1 G6711 (.A1(W14800), .A2(W6936), .ZN(W20437));
  NOR2X1 G6712 (.A1(W10579), .A2(W16280), .ZN(W20434));
  NOR2X1 G6713 (.A1(W790), .A2(W6810), .ZN(W14814));
  NOR2X1 G6714 (.A1(W4843), .A2(I1516), .ZN(W14813));
  NOR2X1 G6715 (.A1(W9940), .A2(W12335), .ZN(O919));
  NOR2X1 G6716 (.A1(W643), .A2(W28540), .ZN(W35995));
  NOR2X1 G6717 (.A1(W5041), .A2(I116), .ZN(W20435));
  NOR2X1 G6718 (.A1(W7110), .A2(W5862), .ZN(W35999));
  NOR2X1 G6719 (.A1(W19253), .A2(I172), .ZN(W20436));
  NOR2X1 G6720 (.A1(W4423), .A2(W12791), .ZN(O921));
  NOR2X1 G6721 (.A1(W18248), .A2(W35827), .ZN(O8136));
  NOR2X1 G6722 (.A1(W2766), .A2(W23654), .ZN(W30355));
  NOR2X1 G6723 (.A1(W8836), .A2(W5653), .ZN(W14804));
  NOR2X1 G6724 (.A1(W391), .A2(W11052), .ZN(W14803));
  NOR2X1 G6725 (.A1(W1686), .A2(W35374), .ZN(O8138));
  NOR2X1 G6726 (.A1(W18221), .A2(W29871), .ZN(O8139));
  NOR2X1 G6727 (.A1(W27852), .A2(W30267), .ZN(O8141));
  NOR2X1 G6728 (.A1(W5891), .A2(W14111), .ZN(O8142));
  NOR2X1 G6729 (.A1(W3137), .A2(W5182), .ZN(O924));
  NOR2X1 G6730 (.A1(W7465), .A2(W855), .ZN(O8119));
  NOR2X1 G6731 (.A1(W1190), .A2(W22), .ZN(W14831));
  NOR2X1 G6732 (.A1(W26025), .A2(W5896), .ZN(W30360));
  NOR2X1 G6733 (.A1(W1985), .A2(W6031), .ZN(W14829));
  NOR2X1 G6734 (.A1(W19044), .A2(W3159), .ZN(W20430));
  NOR2X1 G6735 (.A1(W33790), .A2(W12253), .ZN(O8121));
  NOR2X1 G6736 (.A1(W12744), .A2(W6426), .ZN(W14826));
  NOR2X1 G6737 (.A1(W2681), .A2(W6067), .ZN(W14825));
  NOR2X1 G6738 (.A1(W28278), .A2(W8069), .ZN(O5296));
  NOR2X1 G6739 (.A1(W27027), .A2(W12092), .ZN(O5297));
  NOR2X1 G6740 (.A1(W16882), .A2(W29220), .ZN(O8123));
  NOR2X1 G6741 (.A1(I628), .A2(W2965), .ZN(O8124));
  NOR2X1 G6742 (.A1(W5534), .A2(W741), .ZN(W35981));
  NOR2X1 G6743 (.A1(W8581), .A2(W6392), .ZN(W30358));
  NOR2X1 G6744 (.A1(W9156), .A2(W20146), .ZN(W35989));
  NOR2X1 G6745 (.A1(W17582), .A2(W19164), .ZN(W30356));
  NOR2X1 G6746 (.A1(W13337), .A2(I827), .ZN(W14771));
  NOR2X1 G6747 (.A1(W6273), .A2(W10663), .ZN(W14779));
  NOR2X1 G6748 (.A1(W13831), .A2(W35978), .ZN(O8158));
  NOR2X1 G6749 (.A1(W4160), .A2(W11687), .ZN(W14777));
  NOR2X1 G6750 (.A1(W3359), .A2(W8170), .ZN(W20447));
  NOR2X1 G6751 (.A1(W29567), .A2(W20859), .ZN(O8160));
  NOR2X1 G6752 (.A1(W9225), .A2(W6937), .ZN(W20448));
  NOR2X1 G6753 (.A1(W326), .A2(W917), .ZN(W14773));
  NOR2X1 G6754 (.A1(W10392), .A2(W9182), .ZN(O914));
  NOR2X1 G6755 (.A1(W25788), .A2(W25482), .ZN(O8157));
  NOR2X1 G6756 (.A1(W6699), .A2(W15793), .ZN(O8161));
  NOR2X1 G6757 (.A1(W14960), .A2(W18365), .ZN(O8162));
  NOR2X1 G6758 (.A1(W429), .A2(W10823), .ZN(W20449));
  NOR2X1 G6759 (.A1(I1915), .A2(W3564), .ZN(W20450));
  NOR2X1 G6760 (.A1(W13406), .A2(W11429), .ZN(O2012));
  NOR2X1 G6761 (.A1(I1045), .A2(W2572), .ZN(W14763));
  NOR2X1 G6762 (.A1(W6032), .A2(W18877), .ZN(W20454));
  NOR2X1 G6763 (.A1(W13702), .A2(I1334), .ZN(O5292));
  NOR2X1 G6764 (.A1(W16012), .A2(I1740), .ZN(W36022));
  NOR2X1 G6765 (.A1(W418), .A2(W11184), .ZN(W14797));
  NOR2X1 G6766 (.A1(W5755), .A2(W19101), .ZN(W20440));
  NOR2X1 G6767 (.A1(W3185), .A2(W7002), .ZN(O917));
  NOR2X1 G6768 (.A1(W9330), .A2(W4608), .ZN(W20441));
  NOR2X1 G6769 (.A1(W20685), .A2(W8379), .ZN(O8147));
  NOR2X1 G6770 (.A1(W9912), .A2(W19778), .ZN(W30353));
  NOR2X1 G6771 (.A1(W6495), .A2(W4038), .ZN(W14791));
  NOR2X1 G6772 (.A1(W29012), .A2(W15429), .ZN(W36021));
  NOR2X1 G6773 (.A1(W4514), .A2(I661), .ZN(W14833));
  NOR2X1 G6774 (.A1(W8516), .A2(W8662), .ZN(O5295));
  NOR2X1 G6775 (.A1(W34828), .A2(W6453), .ZN(O8149));
  NOR2X1 G6776 (.A1(W23520), .A2(W25497), .ZN(W30350));
  NOR2X1 G6777 (.A1(W11583), .A2(I603), .ZN(W14785));
  NOR2X1 G6778 (.A1(W940), .A2(W22538), .ZN(W30349));
  NOR2X1 G6779 (.A1(W18186), .A2(W4133), .ZN(O8153));
  NOR2X1 G6780 (.A1(W11148), .A2(W14455), .ZN(W14781));
  NOR2X1 G6781 (.A1(W6727), .A2(W11602), .ZN(W30384));
  NOR2X1 G6782 (.A1(W35703), .A2(W33837), .ZN(O8073));
  NOR2X1 G6783 (.A1(W25699), .A2(W11084), .ZN(O5310));
  NOR2X1 G6784 (.A1(W34719), .A2(W18218), .ZN(O8075));
  NOR2X1 G6785 (.A1(W20374), .A2(W29269), .ZN(W30388));
  NOR2X1 G6786 (.A1(W4682), .A2(I934), .ZN(O5308));
  NOR2X1 G6787 (.A1(I1663), .A2(W12840), .ZN(W14890));
  NOR2X1 G6788 (.A1(W23735), .A2(W9838), .ZN(W35908));
  NOR2X1 G6789 (.A1(I216), .A2(W9118), .ZN(W35909));
  NOR2X1 G6790 (.A1(I711), .A2(W198), .ZN(O8072));
  NOR2X1 G6791 (.A1(W259), .A2(W10686), .ZN(W14884));
  NOR2X1 G6792 (.A1(W15036), .A2(W4148), .ZN(O2002));
  NOR2X1 G6793 (.A1(W11507), .A2(W11162), .ZN(O8082));
  NOR2X1 G6794 (.A1(W1508), .A2(W14382), .ZN(W14881));
  NOR2X1 G6795 (.A1(W13735), .A2(W5602), .ZN(W14880));
  NOR2X1 G6796 (.A1(W8908), .A2(W29362), .ZN(O8085));
  NOR2X1 G6797 (.A1(W20078), .A2(W3685), .ZN(W30382));
  NOR2X1 G6798 (.A1(W2223), .A2(I950), .ZN(W14877));
  NOR2X1 G6799 (.A1(W7687), .A2(W23556), .ZN(O8062));
  NOR2X1 G6800 (.A1(W7190), .A2(W12129), .ZN(W14912));
  NOR2X1 G6801 (.A1(W9108), .A2(W9350), .ZN(W14911));
  NOR2X1 G6802 (.A1(W1492), .A2(W13084), .ZN(W14910));
  NOR2X1 G6803 (.A1(W142), .A2(W29045), .ZN(W35879));
  NOR2X1 G6804 (.A1(W3596), .A2(W7442), .ZN(W14908));
  NOR2X1 G6805 (.A1(W15855), .A2(I20), .ZN(W35880));
  NOR2X1 G6806 (.A1(W595), .A2(W16393), .ZN(W35881));
  NOR2X1 G6807 (.A1(W16036), .A2(W7459), .ZN(W20397));
  NOR2X1 G6808 (.A1(W23417), .A2(W13466), .ZN(W35920));
  NOR2X1 G6809 (.A1(W22886), .A2(I137), .ZN(O8063));
  NOR2X1 G6810 (.A1(W23086), .A2(W13129), .ZN(O5312));
  NOR2X1 G6811 (.A1(W2686), .A2(W28783), .ZN(W35889));
  NOR2X1 G6812 (.A1(W23326), .A2(I1508), .ZN(O8066));
  NOR2X1 G6813 (.A1(W16594), .A2(W860), .ZN(W30392));
  NOR2X1 G6814 (.A1(W6558), .A2(W2528), .ZN(W20400));
  NOR2X1 G6815 (.A1(W5334), .A2(W9421), .ZN(W14897));
  NOR2X1 G6816 (.A1(W497), .A2(W8467), .ZN(W14844));
  NOR2X1 G6817 (.A1(W1271), .A2(W5478), .ZN(O928));
  NOR2X1 G6818 (.A1(W9174), .A2(W9262), .ZN(W14852));
  NOR2X1 G6819 (.A1(W21243), .A2(I447), .ZN(W35954));
  NOR2X1 G6820 (.A1(W6105), .A2(W8675), .ZN(O927));
  NOR2X1 G6821 (.A1(W9869), .A2(W5491), .ZN(O8109));
  NOR2X1 G6822 (.A1(W13159), .A2(W14790), .ZN(O926));
  NOR2X1 G6823 (.A1(I988), .A2(W11071), .ZN(W14846));
  NOR2X1 G6824 (.A1(W6751), .A2(W13598), .ZN(W14845));
  NOR2X1 G6825 (.A1(I12), .A2(W15354), .ZN(O2007));
  NOR2X1 G6826 (.A1(W2374), .A2(W4359), .ZN(W20423));
  NOR2X1 G6827 (.A1(W14840), .A2(W119), .ZN(O2009));
  NOR2X1 G6828 (.A1(W24042), .A2(W9725), .ZN(W30364));
  NOR2X1 G6829 (.A1(W24840), .A2(W18293), .ZN(W30363));
  NOR2X1 G6830 (.A1(W34417), .A2(W15664), .ZN(O8115));
  NOR2X1 G6831 (.A1(W19744), .A2(W11980), .ZN(O8116));
  NOR2X1 G6832 (.A1(W976), .A2(W12191), .ZN(W14836));
  NOR2X1 G6833 (.A1(W6538), .A2(W5985), .ZN(W14835));
  NOR2X1 G6834 (.A1(W13506), .A2(W4243), .ZN(O5305));
  NOR2X1 G6835 (.A1(W4275), .A2(W3981), .ZN(W30379));
  NOR2X1 G6836 (.A1(W2916), .A2(W1390), .ZN(W20410));
  NOR2X1 G6837 (.A1(W13343), .A2(W5001), .ZN(W14873));
  NOR2X1 G6838 (.A1(W5254), .A2(W10392), .ZN(W14872));
  NOR2X1 G6839 (.A1(W9744), .A2(W5691), .ZN(O2004));
  NOR2X1 G6840 (.A1(W9531), .A2(W942), .ZN(W20412));
  NOR2X1 G6841 (.A1(W5291), .A2(W4085), .ZN(W14869));
  NOR2X1 G6842 (.A1(W53), .A2(W11921), .ZN(O8090));
  NOR2X1 G6843 (.A1(I1177), .A2(W520), .ZN(W14760));
  NOR2X1 G6844 (.A1(W9465), .A2(W3389), .ZN(W14866));
  NOR2X1 G6845 (.A1(W14722), .A2(W18775), .ZN(W35932));
  NOR2X1 G6846 (.A1(I306), .A2(W16200), .ZN(W35934));
  NOR2X1 G6847 (.A1(W28157), .A2(W20297), .ZN(O8097));
  NOR2X1 G6848 (.A1(W27514), .A2(W25054), .ZN(W30373));
  NOR2X1 G6849 (.A1(W31042), .A2(W33306), .ZN(O8099));
  NOR2X1 G6850 (.A1(W19782), .A2(W15964), .ZN(W20418));
  NOR2X1 G6851 (.A1(W5290), .A2(W14523), .ZN(W14650));
  NOR2X1 G6852 (.A1(W7998), .A2(W8645), .ZN(W14658));
  NOR2X1 G6853 (.A1(I798), .A2(W6752), .ZN(W30297));
  NOR2X1 G6854 (.A1(W3250), .A2(W14906), .ZN(W36162));
  NOR2X1 G6855 (.A1(W3993), .A2(W11636), .ZN(W14655));
  NOR2X1 G6856 (.A1(W19501), .A2(W16572), .ZN(O8235));
  NOR2X1 G6857 (.A1(W5462), .A2(W6597), .ZN(W14653));
  NOR2X1 G6858 (.A1(W11879), .A2(W7697), .ZN(W30296));
  NOR2X1 G6859 (.A1(W18013), .A2(W8204), .ZN(W36165));
  NOR2X1 G6860 (.A1(W8029), .A2(W12885), .ZN(W14659));
  NOR2X1 G6861 (.A1(W13624), .A2(W13431), .ZN(W14649));
  NOR2X1 G6862 (.A1(W16930), .A2(W12866), .ZN(O5275));
  NOR2X1 G6863 (.A1(W2880), .A2(W20406), .ZN(W20500));
  NOR2X1 G6864 (.A1(W14280), .A2(W10598), .ZN(W14646));
  NOR2X1 G6865 (.A1(W11941), .A2(W7727), .ZN(O895));
  NOR2X1 G6866 (.A1(W29837), .A2(W347), .ZN(W36168));
  NOR2X1 G6867 (.A1(W34511), .A2(W6239), .ZN(O8238));
  NOR2X1 G6868 (.A1(W13624), .A2(W5896), .ZN(W20501));
  NOR2X1 G6869 (.A1(W11893), .A2(W15710), .ZN(O5276));
  NOR2X1 G6870 (.A1(I872), .A2(W3428), .ZN(O897));
  NOR2X1 G6871 (.A1(W7084), .A2(W32719), .ZN(W36147));
  NOR2X1 G6872 (.A1(W10316), .A2(W5898), .ZN(W14674));
  NOR2X1 G6873 (.A1(W10959), .A2(W7994), .ZN(O896));
  NOR2X1 G6874 (.A1(W17001), .A2(W15487), .ZN(O5277));
  NOR2X1 G6875 (.A1(W1576), .A2(W12706), .ZN(W14671));
  NOR2X1 G6876 (.A1(W31369), .A2(W12730), .ZN(O8227));
  NOR2X1 G6877 (.A1(W7198), .A2(W23821), .ZN(O8228));
  NOR2X1 G6878 (.A1(W30144), .A2(W19682), .ZN(W36171));
  NOR2X1 G6879 (.A1(W33860), .A2(W265), .ZN(O8231));
  NOR2X1 G6880 (.A1(W2003), .A2(W5464), .ZN(W14666));
  NOR2X1 G6881 (.A1(I1851), .A2(W1165), .ZN(W14665));
  NOR2X1 G6882 (.A1(W6133), .A2(W6704), .ZN(W14664));
  NOR2X1 G6883 (.A1(W973), .A2(W5445), .ZN(O8233));
  NOR2X1 G6884 (.A1(W797), .A2(W8430), .ZN(W20496));
  NOR2X1 G6885 (.A1(W8391), .A2(I104), .ZN(W14660));
  NOR2X1 G6886 (.A1(W4854), .A2(W221), .ZN(W14609));
  NOR2X1 G6887 (.A1(W29742), .A2(W2499), .ZN(W36202));
  NOR2X1 G6888 (.A1(W123), .A2(W2972), .ZN(O8256));
  NOR2X1 G6889 (.A1(W8544), .A2(W13130), .ZN(W14615));
  NOR2X1 G6890 (.A1(W1676), .A2(W9301), .ZN(W14614));
  NOR2X1 G6891 (.A1(W5251), .A2(W8745), .ZN(W36206));
  NOR2X1 G6892 (.A1(I635), .A2(I729), .ZN(W14612));
  NOR2X1 G6893 (.A1(W166), .A2(W3115), .ZN(W14611));
  NOR2X1 G6894 (.A1(I1819), .A2(I270), .ZN(O8258));
  NOR2X1 G6895 (.A1(W15672), .A2(W10345), .ZN(W30275));
  NOR2X1 G6896 (.A1(W7532), .A2(W9691), .ZN(W14608));
  NOR2X1 G6897 (.A1(W14936), .A2(W22939), .ZN(O8259));
  NOR2X1 G6898 (.A1(W5826), .A2(W25871), .ZN(W30274));
  NOR2X1 G6899 (.A1(W7197), .A2(W3900), .ZN(W14605));
  NOR2X1 G6900 (.A1(W14065), .A2(W21549), .ZN(W30271));
  NOR2X1 G6901 (.A1(W10270), .A2(W11750), .ZN(W20516));
  NOR2X1 G6902 (.A1(W13377), .A2(W21421), .ZN(O8261));
  NOR2X1 G6903 (.A1(W4022), .A2(W7624), .ZN(W14601));
  NOR2X1 G6904 (.A1(W33246), .A2(W18109), .ZN(O8250));
  NOR2X1 G6905 (.A1(W8548), .A2(W1514), .ZN(O8241));
  NOR2X1 G6906 (.A1(W27469), .A2(W33275), .ZN(O8243));
  NOR2X1 G6907 (.A1(W9778), .A2(W14419), .ZN(W36178));
  NOR2X1 G6908 (.A1(W25351), .A2(W12375), .ZN(O8244));
  NOR2X1 G6909 (.A1(W15659), .A2(W21704), .ZN(O5273));
  NOR2X1 G6910 (.A1(W7715), .A2(I621), .ZN(W14634));
  NOR2X1 G6911 (.A1(W18030), .A2(W8636), .ZN(O2019));
  NOR2X1 G6912 (.A1(W33859), .A2(W20071), .ZN(W36188));
  NOR2X1 G6913 (.A1(W1700), .A2(W6733), .ZN(W36146));
  NOR2X1 G6914 (.A1(W548), .A2(W25663), .ZN(W30282));
  NOR2X1 G6915 (.A1(W12016), .A2(I813), .ZN(O890));
  NOR2X1 G6916 (.A1(W9963), .A2(W25987), .ZN(W30281));
  NOR2X1 G6917 (.A1(W1583), .A2(W27203), .ZN(W30276));
  NOR2X1 G6918 (.A1(W13505), .A2(W9001), .ZN(W14621));
  NOR2X1 G6919 (.A1(W12289), .A2(W13338), .ZN(W36198));
  NOR2X1 G6920 (.A1(W10417), .A2(W850), .ZN(W36199));
  NOR2X1 G6921 (.A1(W4587), .A2(W17657), .ZN(W20473));
  NOR2X1 G6922 (.A1(I1395), .A2(W27039), .ZN(W30333));
  NOR2X1 G6923 (.A1(W1033), .A2(W30020), .ZN(W36071));
  NOR2X1 G6924 (.A1(W9268), .A2(W763), .ZN(O8184));
  NOR2X1 G6925 (.A1(W4794), .A2(W622), .ZN(W14732));
  NOR2X1 G6926 (.A1(W14800), .A2(W17679), .ZN(O5284));
  NOR2X1 G6927 (.A1(I1619), .A2(W5544), .ZN(W14727));
  NOR2X1 G6928 (.A1(W6875), .A2(W29244), .ZN(W36084));
  NOR2X1 G6929 (.A1(W10831), .A2(W1539), .ZN(W14725));
  NOR2X1 G6930 (.A1(W17622), .A2(W14929), .ZN(O5289));
  NOR2X1 G6931 (.A1(W5611), .A2(W22790), .ZN(W30321));
  NOR2X1 G6932 (.A1(W13405), .A2(W14703), .ZN(W36089));
  NOR2X1 G6933 (.A1(W5326), .A2(W9470), .ZN(O909));
  NOR2X1 G6934 (.A1(W5058), .A2(W17317), .ZN(W20475));
  NOR2X1 G6935 (.A1(W27622), .A2(W19292), .ZN(O8196));
  NOR2X1 G6936 (.A1(W12502), .A2(W1012), .ZN(W36095));
  NOR2X1 G6937 (.A1(W13695), .A2(W6981), .ZN(O906));
  NOR2X1 G6938 (.A1(W34408), .A2(W10291), .ZN(O8197));
  NOR2X1 G6939 (.A1(I648), .A2(W14430), .ZN(W14750));
  NOR2X1 G6940 (.A1(W1341), .A2(W9254), .ZN(W14759));
  NOR2X1 G6941 (.A1(W15405), .A2(W13542), .ZN(W20457));
  NOR2X1 G6942 (.A1(W1817), .A2(W29473), .ZN(O5291));
  NOR2X1 G6943 (.A1(I1259), .A2(W13648), .ZN(O913));
  NOR2X1 G6944 (.A1(W8028), .A2(I1665), .ZN(W14754));
  NOR2X1 G6945 (.A1(W3386), .A2(W805), .ZN(W14753));
  NOR2X1 G6946 (.A1(W135), .A2(I1216), .ZN(W30339));
  NOR2X1 G6947 (.A1(W6220), .A2(W23539), .ZN(O8173));
  NOR2X1 G6948 (.A1(W7), .A2(I1147), .ZN(W14715));
  NOR2X1 G6949 (.A1(W11820), .A2(W7896), .ZN(W14749));
  NOR2X1 G6950 (.A1(W4849), .A2(W24331), .ZN(O8174));
  NOR2X1 G6951 (.A1(W10300), .A2(W7344), .ZN(W14747));
  NOR2X1 G6952 (.A1(W6185), .A2(I1619), .ZN(W14746));
  NOR2X1 G6953 (.A1(W15785), .A2(W28672), .ZN(O8175));
  NOR2X1 G6954 (.A1(W16487), .A2(W11972), .ZN(W30335));
  NOR2X1 G6955 (.A1(W21208), .A2(W11448), .ZN(W36063));
  NOR2X1 G6956 (.A1(W11715), .A2(W12595), .ZN(W14687));
  NOR2X1 G6957 (.A1(W27068), .A2(W24252), .ZN(W30315));
  NOR2X1 G6958 (.A1(W34866), .A2(W32458), .ZN(O8213));
  NOR2X1 G6959 (.A1(W19212), .A2(W14585), .ZN(O5282));
  NOR2X1 G6960 (.A1(W22673), .A2(W9188), .ZN(W30307));
  NOR2X1 G6961 (.A1(W16316), .A2(W9015), .ZN(O8217));
  NOR2X1 G6962 (.A1(W13895), .A2(W9090), .ZN(W14690));
  NOR2X1 G6963 (.A1(W13413), .A2(W24919), .ZN(O8218));
  NOR2X1 G6964 (.A1(W1987), .A2(W26555), .ZN(W30306));
  NOR2X1 G6965 (.A1(W12835), .A2(W4947), .ZN(W14697));
  NOR2X1 G6966 (.A1(W12757), .A2(W9893), .ZN(W14686));
  NOR2X1 G6967 (.A1(W6740), .A2(W14898), .ZN(W36131));
  NOR2X1 G6968 (.A1(I943), .A2(W12043), .ZN(W20489));
  NOR2X1 G6969 (.A1(W20275), .A2(W8234), .ZN(O8223));
  NOR2X1 G6970 (.A1(W2597), .A2(W17706), .ZN(W30305));
  NOR2X1 G6971 (.A1(I1031), .A2(W2248), .ZN(O899));
  NOR2X1 G6972 (.A1(W2512), .A2(I1672), .ZN(O898));
  NOR2X1 G6973 (.A1(W6881), .A2(W2689), .ZN(O5279));
  NOR2X1 G6974 (.A1(W28355), .A2(W8472), .ZN(O5283));
  NOR2X1 G6975 (.A1(W12836), .A2(W12880), .ZN(W20476));
  NOR2X1 G6976 (.A1(W4950), .A2(W18946), .ZN(O2015));
  NOR2X1 G6977 (.A1(I934), .A2(I290), .ZN(W36103));
  NOR2X1 G6978 (.A1(W14283), .A2(W14916), .ZN(W20478));
  NOR2X1 G6979 (.A1(W15048), .A2(W10913), .ZN(W20479));
  NOR2X1 G6980 (.A1(W16781), .A2(W29151), .ZN(W30319));
  NOR2X1 G6981 (.A1(W2023), .A2(W12954), .ZN(O905));
  NOR2X1 G6982 (.A1(W1315), .A2(I684), .ZN(W14707));
  NOR2X1 G6983 (.A1(W9560), .A2(W9172), .ZN(W14913));
  NOR2X1 G6984 (.A1(W19318), .A2(W27457), .ZN(W30317));
  NOR2X1 G6985 (.A1(W4631), .A2(W13135), .ZN(W14704));
  NOR2X1 G6986 (.A1(W20542), .A2(W33446), .ZN(W36111));
  NOR2X1 G6987 (.A1(W32636), .A2(W25861), .ZN(O8207));
  NOR2X1 G6988 (.A1(W23411), .A2(W30759), .ZN(O8209));
  NOR2X1 G6989 (.A1(W14205), .A2(W29396), .ZN(O8210));
  NOR2X1 G6990 (.A1(W21562), .A2(W19487), .ZN(O8211));
  NOR2X1 G6991 (.A1(W16205), .A2(W18834), .ZN(W20316));
  NOR2X1 G6992 (.A1(W31342), .A2(W1718), .ZN(W35671));
  NOR2X1 G6993 (.A1(W11208), .A2(W15970), .ZN(O5352));
  NOR2X1 G6994 (.A1(W1023), .A2(W6165), .ZN(O5350));
  NOR2X1 G6995 (.A1(W2386), .A2(W10927), .ZN(W15133));
  NOR2X1 G6996 (.A1(W7297), .A2(W2843), .ZN(O7958));
  NOR2X1 G6997 (.A1(W2069), .A2(W5105), .ZN(W15130));
  NOR2X1 G6998 (.A1(W10292), .A2(W20532), .ZN(O7959));
  NOR2X1 G6999 (.A1(W10074), .A2(W3018), .ZN(W15128));
  NOR2X1 G7000 (.A1(W29900), .A2(W7661), .ZN(W30471));
  NOR2X1 G7001 (.A1(I1392), .A2(W5067), .ZN(W15126));
  NOR2X1 G7002 (.A1(W3175), .A2(W11265), .ZN(O965));
  NOR2X1 G7003 (.A1(W20749), .A2(W575), .ZN(O7962));
  NOR2X1 G7004 (.A1(W8448), .A2(W349), .ZN(W15122));
  NOR2X1 G7005 (.A1(W9669), .A2(I1412), .ZN(O963));
  NOR2X1 G7006 (.A1(W32946), .A2(W5314), .ZN(W35685));
  NOR2X1 G7007 (.A1(W13809), .A2(W24796), .ZN(O5348));
  NOR2X1 G7008 (.A1(W14959), .A2(W15384), .ZN(W20319));
  NOR2X1 G7009 (.A1(W12855), .A2(W13468), .ZN(W15146));
  NOR2X1 G7010 (.A1(W1999), .A2(W2629), .ZN(W15155));
  NOR2X1 G7011 (.A1(W23750), .A2(W10048), .ZN(W30477));
  NOR2X1 G7012 (.A1(W18105), .A2(W13822), .ZN(W20308));
  NOR2X1 G7013 (.A1(W22338), .A2(W30559), .ZN(O7945));
  NOR2X1 G7014 (.A1(W27615), .A2(W26685), .ZN(W35659));
  NOR2X1 G7015 (.A1(W2165), .A2(W19620), .ZN(O7947));
  NOR2X1 G7016 (.A1(W9039), .A2(W14867), .ZN(W15149));
  NOR2X1 G7017 (.A1(W31384), .A2(W4357), .ZN(W35662));
  NOR2X1 G7018 (.A1(W17058), .A2(W4008), .ZN(W20320));
  NOR2X1 G7019 (.A1(I917), .A2(W4884), .ZN(O968));
  NOR2X1 G7020 (.A1(W17147), .A2(W27818), .ZN(O5353));
  NOR2X1 G7021 (.A1(I922), .A2(I664), .ZN(W15143));
  NOR2X1 G7022 (.A1(W7227), .A2(W4365), .ZN(W15142));
  NOR2X1 G7023 (.A1(W2274), .A2(W14938), .ZN(W15141));
  NOR2X1 G7024 (.A1(W5977), .A2(W32945), .ZN(O7951));
  NOR2X1 G7025 (.A1(W23654), .A2(W9532), .ZN(O7952));
  NOR2X1 G7026 (.A1(W7395), .A2(W9329), .ZN(W15086));
  NOR2X1 G7027 (.A1(W11593), .A2(W6508), .ZN(W15095));
  NOR2X1 G7028 (.A1(W8320), .A2(W5066), .ZN(W15093));
  NOR2X1 G7029 (.A1(W1630), .A2(W10111), .ZN(W35707));
  NOR2X1 G7030 (.A1(W2049), .A2(W10269), .ZN(W15091));
  NOR2X1 G7031 (.A1(W29899), .A2(W2154), .ZN(O7970));
  NOR2X1 G7032 (.A1(W13271), .A2(W6287), .ZN(O7971));
  NOR2X1 G7033 (.A1(W6038), .A2(I60), .ZN(W15088));
  NOR2X1 G7034 (.A1(W13035), .A2(I1528), .ZN(W20329));
  NOR2X1 G7035 (.A1(W9350), .A2(I162), .ZN(W15097));
  NOR2X1 G7036 (.A1(I825), .A2(W5904), .ZN(W15085));
  NOR2X1 G7037 (.A1(W27942), .A2(W4717), .ZN(W35714));
  NOR2X1 G7038 (.A1(W10620), .A2(W6599), .ZN(W15082));
  NOR2X1 G7039 (.A1(W5718), .A2(W16566), .ZN(W20331));
  NOR2X1 G7040 (.A1(W24551), .A2(W8744), .ZN(O7976));
  NOR2X1 G7041 (.A1(W2227), .A2(W10824), .ZN(W15079));
  NOR2X1 G7042 (.A1(W10994), .A2(W6260), .ZN(W15078));
  NOR2X1 G7043 (.A1(W29870), .A2(W5540), .ZN(O7977));
  NOR2X1 G7044 (.A1(W6596), .A2(W5488), .ZN(W15106));
  NOR2X1 G7045 (.A1(W8032), .A2(W1349), .ZN(W35691));
  NOR2X1 G7046 (.A1(W4790), .A2(W9083), .ZN(W15115));
  NOR2X1 G7047 (.A1(W16088), .A2(W576), .ZN(O5347));
  NOR2X1 G7048 (.A1(W7809), .A2(W4816), .ZN(W15113));
  NOR2X1 G7049 (.A1(W23656), .A2(W7465), .ZN(O5343));
  NOR2X1 G7050 (.A1(W4532), .A2(W13131), .ZN(W15109));
  NOR2X1 G7051 (.A1(W30590), .A2(W30239), .ZN(W35697));
  NOR2X1 G7052 (.A1(W9537), .A2(I1154), .ZN(W15107));
  NOR2X1 G7053 (.A1(W30444), .A2(W12850), .ZN(O7941));
  NOR2X1 G7054 (.A1(W82), .A2(W13503), .ZN(W15105));
  NOR2X1 G7055 (.A1(W289), .A2(W9595), .ZN(W20325));
  NOR2X1 G7056 (.A1(W9582), .A2(W9214), .ZN(O960));
  NOR2X1 G7057 (.A1(W7255), .A2(W2074), .ZN(W15102));
  NOR2X1 G7058 (.A1(W8695), .A2(W7911), .ZN(W15101));
  NOR2X1 G7059 (.A1(W33215), .A2(I1738), .ZN(O7969));
  NOR2X1 G7060 (.A1(W9085), .A2(W12323), .ZN(W15098));
  NOR2X1 G7061 (.A1(W33299), .A2(W18060), .ZN(O7908));
  NOR2X1 G7062 (.A1(W30349), .A2(W25393), .ZN(W35591));
  NOR2X1 G7063 (.A1(W11183), .A2(W11999), .ZN(W15214));
  NOR2X1 G7064 (.A1(W27868), .A2(W26), .ZN(O7904));
  NOR2X1 G7065 (.A1(W10104), .A2(W17053), .ZN(O7905));
  NOR2X1 G7066 (.A1(W1502), .A2(W14236), .ZN(W15211));
  NOR2X1 G7067 (.A1(W18750), .A2(W14018), .ZN(W20290));
  NOR2X1 G7068 (.A1(W8483), .A2(W12779), .ZN(W15207));
  NOR2X1 G7069 (.A1(W33501), .A2(W168), .ZN(O7907));
  NOR2X1 G7070 (.A1(W5963), .A2(W1995), .ZN(W15216));
  NOR2X1 G7071 (.A1(I895), .A2(W5878), .ZN(W15204));
  NOR2X1 G7072 (.A1(W547), .A2(W3389), .ZN(W15202));
  NOR2X1 G7073 (.A1(W15426), .A2(W223), .ZN(O7911));
  NOR2X1 G7074 (.A1(W18315), .A2(W18357), .ZN(O7912));
  NOR2X1 G7075 (.A1(W1757), .A2(W3113), .ZN(W15199));
  NOR2X1 G7076 (.A1(W23801), .A2(W34303), .ZN(O7914));
  NOR2X1 G7077 (.A1(W13422), .A2(W7494), .ZN(O7915));
  NOR2X1 G7078 (.A1(W23997), .A2(W24988), .ZN(O5364));
  NOR2X1 G7079 (.A1(W6806), .A2(W8022), .ZN(W20283));
  NOR2X1 G7080 (.A1(W7868), .A2(W13216), .ZN(W15239));
  NOR2X1 G7081 (.A1(W17310), .A2(W7692), .ZN(W20277));
  NOR2X1 G7082 (.A1(W13809), .A2(W19213), .ZN(O5372));
  NOR2X1 G7083 (.A1(W14606), .A2(W9376), .ZN(O7888));
  NOR2X1 G7084 (.A1(W13324), .A2(W4421), .ZN(W35573));
  NOR2X1 G7085 (.A1(W14724), .A2(W231), .ZN(W15232));
  NOR2X1 G7086 (.A1(W7127), .A2(W5730), .ZN(W15231));
  NOR2X1 G7087 (.A1(W1304), .A2(W5299), .ZN(W15230));
  NOR2X1 G7088 (.A1(W4072), .A2(W33439), .ZN(O7918));
  NOR2X1 G7089 (.A1(W953), .A2(W12126), .ZN(W20285));
  NOR2X1 G7090 (.A1(W10226), .A2(W31627), .ZN(W35584));
  NOR2X1 G7091 (.A1(W14646), .A2(W2673), .ZN(W15221));
  NOR2X1 G7092 (.A1(W17641), .A2(W141), .ZN(W20287));
  NOR2X1 G7093 (.A1(W3440), .A2(W4445), .ZN(W15219));
  NOR2X1 G7094 (.A1(W27349), .A2(W1894), .ZN(W30502));
  NOR2X1 G7095 (.A1(W9807), .A2(W20925), .ZN(O7901));
  NOR2X1 G7096 (.A1(W30005), .A2(W28076), .ZN(W35640));
  NOR2X1 G7097 (.A1(W4868), .A2(W9956), .ZN(W15175));
  NOR2X1 G7098 (.A1(W13261), .A2(W7370), .ZN(W15174));
  NOR2X1 G7099 (.A1(W30704), .A2(W1943), .ZN(W35634));
  NOR2X1 G7100 (.A1(W12610), .A2(W31233), .ZN(W35636));
  NOR2X1 G7101 (.A1(W3937), .A2(W8518), .ZN(O5360));
  NOR2X1 G7102 (.A1(W12939), .A2(W1287), .ZN(W30484));
  NOR2X1 G7103 (.A1(W12377), .A2(W6991), .ZN(W15169));
  NOR2X1 G7104 (.A1(W3144), .A2(W9499), .ZN(W15168));
  NOR2X1 G7105 (.A1(W3777), .A2(W9411), .ZN(O7929));
  NOR2X1 G7106 (.A1(I944), .A2(W945), .ZN(W15165));
  NOR2X1 G7107 (.A1(W35229), .A2(W27891), .ZN(O7936));
  NOR2X1 G7108 (.A1(W5500), .A2(W5392), .ZN(W20304));
  NOR2X1 G7109 (.A1(I813), .A2(W5921), .ZN(W15162));
  NOR2X1 G7110 (.A1(W12809), .A2(W7087), .ZN(O5358));
  NOR2X1 G7111 (.A1(W11810), .A2(W4650), .ZN(W15160));
  NOR2X1 G7112 (.A1(W34707), .A2(W25969), .ZN(O7937));
  NOR2X1 G7113 (.A1(W3160), .A2(W14639), .ZN(O969));
  NOR2X1 G7114 (.A1(W11982), .A2(W8608), .ZN(W15185));
  NOR2X1 G7115 (.A1(W35421), .A2(W5110), .ZN(O7919));
  NOR2X1 G7116 (.A1(I253), .A2(W17049), .ZN(O7920));
  NOR2X1 G7117 (.A1(I1243), .A2(W8100), .ZN(O5363));
  NOR2X1 G7118 (.A1(I1455), .A2(W7088), .ZN(O7922));
  NOR2X1 G7119 (.A1(W9963), .A2(W5815), .ZN(W15189));
  NOR2X1 G7120 (.A1(W11462), .A2(W14061), .ZN(W15188));
  NOR2X1 G7121 (.A1(W2557), .A2(W9975), .ZN(W30491));
  NOR2X1 G7122 (.A1(W7262), .A2(W13093), .ZN(W15186));
  NOR2X1 G7123 (.A1(W25236), .A2(W31733), .ZN(O7978));
  NOR2X1 G7124 (.A1(W29164), .A2(W10), .ZN(W30490));
  NOR2X1 G7125 (.A1(W7687), .A2(W25272), .ZN(W30488));
  NOR2X1 G7126 (.A1(W6171), .A2(W3183), .ZN(W15182));
  NOR2X1 G7127 (.A1(W1462), .A2(W11923), .ZN(O1971));
  NOR2X1 G7128 (.A1(W2473), .A2(W11888), .ZN(W15180));
  NOR2X1 G7129 (.A1(W31522), .A2(W11871), .ZN(W35630));
  NOR2X1 G7130 (.A1(W5732), .A2(W33469), .ZN(O7928));
  NOR2X1 G7131 (.A1(W8121), .A2(W4957), .ZN(W20372));
  NOR2X1 G7132 (.A1(W1795), .A2(W1224), .ZN(O8024));
  NOR2X1 G7133 (.A1(W20105), .A2(W16151), .ZN(W20368));
  NOR2X1 G7134 (.A1(W34833), .A2(W22933), .ZN(W35813));
  NOR2X1 G7135 (.A1(I572), .A2(W1974), .ZN(W14970));
  NOR2X1 G7136 (.A1(W16662), .A2(W3949), .ZN(O8026));
  NOR2X1 G7137 (.A1(W1323), .A2(W13081), .ZN(O8027));
  NOR2X1 G7138 (.A1(W5387), .A2(W4051), .ZN(W14967));
  NOR2X1 G7139 (.A1(W15417), .A2(W750), .ZN(W30419));
  NOR2X1 G7140 (.A1(W26082), .A2(W11474), .ZN(O5328));
  NOR2X1 G7141 (.A1(W16524), .A2(W5934), .ZN(W20374));
  NOR2X1 G7142 (.A1(I1317), .A2(W8427), .ZN(W20375));
  NOR2X1 G7143 (.A1(W11067), .A2(I1712), .ZN(W20377));
  NOR2X1 G7144 (.A1(W11407), .A2(W10697), .ZN(O937));
  NOR2X1 G7145 (.A1(W7197), .A2(W12372), .ZN(W35829));
  NOR2X1 G7146 (.A1(W7434), .A2(W2656), .ZN(W14956));
  NOR2X1 G7147 (.A1(W6530), .A2(W11916), .ZN(O8033));
  NOR2X1 G7148 (.A1(W1207), .A2(W33511), .ZN(O8034));
  NOR2X1 G7149 (.A1(W3056), .A2(W1361), .ZN(W14986));
  NOR2X1 G7150 (.A1(W6174), .A2(I1012), .ZN(O8013));
  NOR2X1 G7151 (.A1(W25745), .A2(W881), .ZN(O8015));
  NOR2X1 G7152 (.A1(W7077), .A2(W13091), .ZN(O1988));
  NOR2X1 G7153 (.A1(W118), .A2(W31480), .ZN(O8019));
  NOR2X1 G7154 (.A1(W4595), .A2(W11675), .ZN(W14992));
  NOR2X1 G7155 (.A1(I1021), .A2(W18214), .ZN(W20361));
  NOR2X1 G7156 (.A1(W20623), .A2(W23931), .ZN(W35799));
  NOR2X1 G7157 (.A1(W3588), .A2(W35196), .ZN(W35800));
  NOR2X1 G7158 (.A1(W12220), .A2(W25958), .ZN(O8035));
  NOR2X1 G7159 (.A1(W5376), .A2(W5725), .ZN(W14985));
  NOR2X1 G7160 (.A1(W10113), .A2(W2663), .ZN(O1990));
  NOR2X1 G7161 (.A1(W21494), .A2(W26707), .ZN(W30426));
  NOR2X1 G7162 (.A1(W4116), .A2(W2811), .ZN(W14981));
  NOR2X1 G7163 (.A1(W8136), .A2(W11543), .ZN(W14980));
  NOR2X1 G7164 (.A1(W7161), .A2(W13691), .ZN(W14979));
  NOR2X1 G7165 (.A1(W759), .A2(W9831), .ZN(W35807));
  NOR2X1 G7166 (.A1(W19638), .A2(W10506), .ZN(O1996));
  NOR2X1 G7167 (.A1(W12930), .A2(W6450), .ZN(W20386));
  NOR2X1 G7168 (.A1(W35781), .A2(W26868), .ZN(W35854));
  NOR2X1 G7169 (.A1(W6127), .A2(W13747), .ZN(W14932));
  NOR2X1 G7170 (.A1(W9363), .A2(W20470), .ZN(O8048));
  NOR2X1 G7171 (.A1(W25529), .A2(W4178), .ZN(O8049));
  NOR2X1 G7172 (.A1(I1045), .A2(W6209), .ZN(W14929));
  NOR2X1 G7173 (.A1(W13947), .A2(W2050), .ZN(W14928));
  NOR2X1 G7174 (.A1(W320), .A2(W14488), .ZN(W14927));
  NOR2X1 G7175 (.A1(W3525), .A2(W2966), .ZN(W35850));
  NOR2X1 G7176 (.A1(W107), .A2(W6608), .ZN(W14925));
  NOR2X1 G7177 (.A1(W20755), .A2(W28202), .ZN(O5317));
  NOR2X1 G7178 (.A1(W29716), .A2(W15285), .ZN(O5316));
  NOR2X1 G7179 (.A1(W10581), .A2(W7535), .ZN(O1999));
  NOR2X1 G7180 (.A1(W14848), .A2(W22051), .ZN(W35871));
  NOR2X1 G7181 (.A1(W11998), .A2(W11798), .ZN(O932));
  NOR2X1 G7182 (.A1(W9409), .A2(W6132), .ZN(W14915));
  NOR2X1 G7183 (.A1(W16410), .A2(W191), .ZN(W20396));
  NOR2X1 G7184 (.A1(W1792), .A2(W16100), .ZN(O1995));
  NOR2X1 G7185 (.A1(W25272), .A2(W9287), .ZN(O8036));
  NOR2X1 G7186 (.A1(W2876), .A2(W10216), .ZN(O1994));
  NOR2X1 G7187 (.A1(W20459), .A2(W24404), .ZN(O8038));
  NOR2X1 G7188 (.A1(W23155), .A2(W28393), .ZN(O5322));
  NOR2X1 G7189 (.A1(W1359), .A2(I1145), .ZN(W20381));
  NOR2X1 G7190 (.A1(W18739), .A2(W12301), .ZN(O8039));
  NOR2X1 G7191 (.A1(W3978), .A2(W5263), .ZN(W14946));
  NOR2X1 G7192 (.A1(W12262), .A2(W11045), .ZN(W14945));
  NOR2X1 G7193 (.A1(W12620), .A2(W12807), .ZN(W14999));
  NOR2X1 G7194 (.A1(W11243), .A2(W10294), .ZN(W30409));
  NOR2X1 G7195 (.A1(W24204), .A2(W10626), .ZN(W30407));
  NOR2X1 G7196 (.A1(W8293), .A2(W3122), .ZN(O933));
  NOR2X1 G7197 (.A1(W31697), .A2(I178), .ZN(W35845));
  NOR2X1 G7198 (.A1(I1944), .A2(W11682), .ZN(W35846));
  NOR2X1 G7199 (.A1(W1738), .A2(W6588), .ZN(W14938));
  NOR2X1 G7200 (.A1(W3323), .A2(W24527), .ZN(W30406));
  NOR2X1 G7201 (.A1(W13348), .A2(W27628), .ZN(W30441));
  NOR2X1 G7202 (.A1(W18337), .A2(W963), .ZN(O7988));
  NOR2X1 G7203 (.A1(W12195), .A2(W31583), .ZN(W35741));
  NOR2X1 G7204 (.A1(W9739), .A2(I533), .ZN(W15053));
  NOR2X1 G7205 (.A1(I1616), .A2(W7270), .ZN(W15052));
  NOR2X1 G7206 (.A1(W14992), .A2(I375), .ZN(W15051));
  NOR2X1 G7207 (.A1(W358), .A2(W12868), .ZN(O953));
  NOR2X1 G7208 (.A1(W7877), .A2(W35435), .ZN(O7991));
  NOR2X1 G7209 (.A1(W1442), .A2(W1745), .ZN(W15048));
  NOR2X1 G7210 (.A1(W11773), .A2(W13085), .ZN(W15056));
  NOR2X1 G7211 (.A1(W7392), .A2(I602), .ZN(W20340));
  NOR2X1 G7212 (.A1(W4114), .A2(W846), .ZN(W15044));
  NOR2X1 G7213 (.A1(W34179), .A2(W22085), .ZN(O7994));
  NOR2X1 G7214 (.A1(W13689), .A2(W5086), .ZN(W20342));
  NOR2X1 G7215 (.A1(W4425), .A2(W1463), .ZN(W15041));
  NOR2X1 G7216 (.A1(W218), .A2(W23283), .ZN(W35749));
  NOR2X1 G7217 (.A1(W9055), .A2(W4607), .ZN(W20343));
  NOR2X1 G7218 (.A1(W152), .A2(W4920), .ZN(O7997));
  NOR2X1 G7219 (.A1(W7362), .A2(W27516), .ZN(W35731));
  NOR2X1 G7220 (.A1(W4188), .A2(W30922), .ZN(O7979));
  NOR2X1 G7221 (.A1(W10402), .A2(I455), .ZN(W20333));
  NOR2X1 G7222 (.A1(W4230), .A2(W3253), .ZN(W15072));
  NOR2X1 G7223 (.A1(W2422), .A2(W12241), .ZN(O5336));
  NOR2X1 G7224 (.A1(W13070), .A2(W2831), .ZN(W15070));
  NOR2X1 G7225 (.A1(W4222), .A2(W16069), .ZN(W35728));
  NOR2X1 G7226 (.A1(W6795), .A2(W6268), .ZN(W15068));
  NOR2X1 G7227 (.A1(W15770), .A2(W9956), .ZN(O1978));
  NOR2X1 G7228 (.A1(W13144), .A2(W14082), .ZN(W15037));
  NOR2X1 G7229 (.A1(W30985), .A2(W30058), .ZN(W35732));
  NOR2X1 G7230 (.A1(W4025), .A2(W6917), .ZN(W30444));
  NOR2X1 G7231 (.A1(W10071), .A2(W9699), .ZN(W15062));
  NOR2X1 G7232 (.A1(W13925), .A2(W3194), .ZN(O955));
  NOR2X1 G7233 (.A1(W8860), .A2(W3120), .ZN(W15060));
  NOR2X1 G7234 (.A1(W11382), .A2(W341), .ZN(O7986));
  NOR2X1 G7235 (.A1(I1574), .A2(W811), .ZN(W15057));
  NOR2X1 G7236 (.A1(W17771), .A2(W7722), .ZN(W20355));
  NOR2X1 G7237 (.A1(W5728), .A2(I904), .ZN(W15017));
  NOR2X1 G7238 (.A1(W13106), .A2(W21754), .ZN(O8005));
  NOR2X1 G7239 (.A1(W1517), .A2(W1602), .ZN(W15015));
  NOR2X1 G7240 (.A1(W10033), .A2(W10330), .ZN(W35773));
  NOR2X1 G7241 (.A1(W16391), .A2(W1352), .ZN(W35774));
  NOR2X1 G7242 (.A1(W2867), .A2(W27997), .ZN(O8007));
  NOR2X1 G7243 (.A1(W22967), .A2(W1896), .ZN(W35779));
  NOR2X1 G7244 (.A1(W8548), .A2(W28180), .ZN(O8008));
  NOR2X1 G7245 (.A1(W5279), .A2(W1546), .ZN(W15018));
  NOR2X1 G7246 (.A1(W4150), .A2(W15781), .ZN(W35782));
  NOR2X1 G7247 (.A1(W10899), .A2(W1769), .ZN(W15007));
  NOR2X1 G7248 (.A1(W1982), .A2(W3614), .ZN(W15006));
  NOR2X1 G7249 (.A1(I1458), .A2(W10095), .ZN(W15005));
  NOR2X1 G7250 (.A1(W6418), .A2(W6687), .ZN(W15003));
  NOR2X1 G7251 (.A1(W3834), .A2(W3064), .ZN(W15002));
  NOR2X1 G7252 (.A1(W6470), .A2(W1260), .ZN(W15001));
  NOR2X1 G7253 (.A1(W31717), .A2(W304), .ZN(O8011));
  NOR2X1 G7254 (.A1(W11791), .A2(W3999), .ZN(W15028));
  NOR2X1 G7255 (.A1(W13100), .A2(W12006), .ZN(W15036));
  NOR2X1 G7256 (.A1(W18173), .A2(W7554), .ZN(O7998));
  NOR2X1 G7257 (.A1(W10463), .A2(W15025), .ZN(O1979));
  NOR2X1 G7258 (.A1(W23809), .A2(W28869), .ZN(O5332));
  NOR2X1 G7259 (.A1(W14184), .A2(W16587), .ZN(W20346));
  NOR2X1 G7260 (.A1(W26547), .A2(W24311), .ZN(W30437));
  NOR2X1 G7261 (.A1(W128), .A2(W32291), .ZN(W35758));
  NOR2X1 G7262 (.A1(W4408), .A2(W10844), .ZN(O1981));
  NOR2X1 G7263 (.A1(W32386), .A2(W7636), .ZN(O8262));
  NOR2X1 G7264 (.A1(W22527), .A2(W10458), .ZN(W30436));
  NOR2X1 G7265 (.A1(W12497), .A2(W3925), .ZN(W20351));
  NOR2X1 G7266 (.A1(W8509), .A2(W7297), .ZN(O946));
  NOR2X1 G7267 (.A1(W12820), .A2(W7399), .ZN(W15023));
  NOR2X1 G7268 (.A1(W16815), .A2(W167), .ZN(W35768));
  NOR2X1 G7269 (.A1(I1173), .A2(W538), .ZN(O1984));
  NOR2X1 G7270 (.A1(W27165), .A2(W28139), .ZN(O5331));
  NOR2X1 G7271 (.A1(W3013), .A2(W9078), .ZN(W14172));
  NOR2X1 G7272 (.A1(W27635), .A2(W7211), .ZN(W30133));
  NOR2X1 G7273 (.A1(W3192), .A2(W32011), .ZN(O8519));
  NOR2X1 G7274 (.A1(W3648), .A2(W5354), .ZN(W14181));
  NOR2X1 G7275 (.A1(W16415), .A2(W24431), .ZN(W36642));
  NOR2X1 G7276 (.A1(W32808), .A2(W23744), .ZN(O8521));
  NOR2X1 G7277 (.A1(W5687), .A2(I10), .ZN(W36645));
  NOR2X1 G7278 (.A1(W10002), .A2(W29332), .ZN(W36647));
  NOR2X1 G7279 (.A1(I1259), .A2(W2789), .ZN(O834));
  NOR2X1 G7280 (.A1(W181), .A2(W8838), .ZN(W20649));
  NOR2X1 G7281 (.A1(W856), .A2(W8590), .ZN(W20654));
  NOR2X1 G7282 (.A1(W5637), .A2(W22407), .ZN(W30125));
  NOR2X1 G7283 (.A1(W8492), .A2(W942), .ZN(W20656));
  NOR2X1 G7284 (.A1(W4902), .A2(W11939), .ZN(W30124));
  NOR2X1 G7285 (.A1(W2015), .A2(W10743), .ZN(W20658));
  NOR2X1 G7286 (.A1(W30555), .A2(W2490), .ZN(O8529));
  NOR2X1 G7287 (.A1(W28423), .A2(I1480), .ZN(W36661));
  NOR2X1 G7288 (.A1(W12474), .A2(W27126), .ZN(O5196));
  NOR2X1 G7289 (.A1(W4167), .A2(W1020), .ZN(W14192));
  NOR2X1 G7290 (.A1(W8775), .A2(W16709), .ZN(O2048));
  NOR2X1 G7291 (.A1(W16475), .A2(W12806), .ZN(O8512));
  NOR2X1 G7292 (.A1(W5919), .A2(W5695), .ZN(W14199));
  NOR2X1 G7293 (.A1(W8375), .A2(W28400), .ZN(W36628));
  NOR2X1 G7294 (.A1(W17852), .A2(W24064), .ZN(O8514));
  NOR2X1 G7295 (.A1(W8458), .A2(W2263), .ZN(W14195));
  NOR2X1 G7296 (.A1(W57), .A2(W18590), .ZN(W36631));
  NOR2X1 G7297 (.A1(W1468), .A2(W1615), .ZN(W14193));
  NOR2X1 G7298 (.A1(W899), .A2(W18188), .ZN(W20660));
  NOR2X1 G7299 (.A1(I1861), .A2(W12861), .ZN(O839));
  NOR2X1 G7300 (.A1(W18691), .A2(W882), .ZN(W36633));
  NOR2X1 G7301 (.A1(W12625), .A2(W5255), .ZN(W14189));
  NOR2X1 G7302 (.A1(I1786), .A2(W10922), .ZN(O838));
  NOR2X1 G7303 (.A1(W9854), .A2(W8909), .ZN(O2050));
  NOR2X1 G7304 (.A1(W17153), .A2(W21763), .ZN(W36635));
  NOR2X1 G7305 (.A1(W20795), .A2(W3223), .ZN(O5199));
  NOR2X1 G7306 (.A1(W2184), .A2(W13128), .ZN(O828));
  NOR2X1 G7307 (.A1(W10026), .A2(W21872), .ZN(O8543));
  NOR2X1 G7308 (.A1(W5780), .A2(W8428), .ZN(W36690));
  NOR2X1 G7309 (.A1(W17027), .A2(W10501), .ZN(W20667));
  NOR2X1 G7310 (.A1(W25488), .A2(W26605), .ZN(O8545));
  NOR2X1 G7311 (.A1(W3904), .A2(W9681), .ZN(W14138));
  NOR2X1 G7312 (.A1(W19942), .A2(W17386), .ZN(O5193));
  NOR2X1 G7313 (.A1(I429), .A2(W396), .ZN(W14136));
  NOR2X1 G7314 (.A1(W5517), .A2(W3330), .ZN(W14135));
  NOR2X1 G7315 (.A1(W7047), .A2(W315), .ZN(W14143));
  NOR2X1 G7316 (.A1(I1339), .A2(W7775), .ZN(W14133));
  NOR2X1 G7317 (.A1(W30574), .A2(W17446), .ZN(O8547));
  NOR2X1 G7318 (.A1(W11518), .A2(W10880), .ZN(W14131));
  NOR2X1 G7319 (.A1(W7022), .A2(W21478), .ZN(O8548));
  NOR2X1 G7320 (.A1(W22967), .A2(W14989), .ZN(W36697));
  NOR2X1 G7321 (.A1(W18270), .A2(W11505), .ZN(W20669));
  NOR2X1 G7322 (.A1(W3483), .A2(W5850), .ZN(W14126));
  NOR2X1 G7323 (.A1(W29943), .A2(W20748), .ZN(W36702));
  NOR2X1 G7324 (.A1(W17579), .A2(W25681), .ZN(O8535));
  NOR2X1 G7325 (.A1(W5060), .A2(W9674), .ZN(O833));
  NOR2X1 G7326 (.A1(W8081), .A2(W10864), .ZN(W20662));
  NOR2X1 G7327 (.A1(W13324), .A2(W26780), .ZN(O8531));
  NOR2X1 G7328 (.A1(W2298), .A2(W22633), .ZN(W36670));
  NOR2X1 G7329 (.A1(W6808), .A2(W6204), .ZN(W14157));
  NOR2X1 G7330 (.A1(W3613), .A2(W7608), .ZN(W36673));
  NOR2X1 G7331 (.A1(W32204), .A2(W35823), .ZN(W36675));
  NOR2X1 G7332 (.A1(W5810), .A2(W13366), .ZN(W14153));
  NOR2X1 G7333 (.A1(W5559), .A2(W2642), .ZN(O842));
  NOR2X1 G7334 (.A1(I358), .A2(W2357), .ZN(W36679));
  NOR2X1 G7335 (.A1(W16611), .A2(W12596), .ZN(W36680));
  NOR2X1 G7336 (.A1(W5370), .A2(W7012), .ZN(O2052));
  NOR2X1 G7337 (.A1(W20992), .A2(W15823), .ZN(W30114));
  NOR2X1 G7338 (.A1(W22047), .A2(W14011), .ZN(O8540));
  NOR2X1 G7339 (.A1(W569), .A2(W11184), .ZN(W14145));
  NOR2X1 G7340 (.A1(W2558), .A2(W20263), .ZN(O8541));
  NOR2X1 G7341 (.A1(W35733), .A2(W6030), .ZN(O8481));
  NOR2X1 G7342 (.A1(W35995), .A2(W9569), .ZN(W36558));
  NOR2X1 G7343 (.A1(I1320), .A2(W26767), .ZN(W36561));
  NOR2X1 G7344 (.A1(W730), .A2(W25868), .ZN(O5212));
  NOR2X1 G7345 (.A1(W2056), .A2(W16094), .ZN(W20621));
  NOR2X1 G7346 (.A1(W35963), .A2(W14588), .ZN(O8476));
  NOR2X1 G7347 (.A1(W20603), .A2(W8509), .ZN(O2044));
  NOR2X1 G7348 (.A1(W35284), .A2(W30873), .ZN(O8479));
  NOR2X1 G7349 (.A1(W9237), .A2(W2977), .ZN(W14257));
  NOR2X1 G7350 (.A1(W51), .A2(I1160), .ZN(W14268));
  NOR2X1 G7351 (.A1(W27136), .A2(W32405), .ZN(O8482));
  NOR2X1 G7352 (.A1(W8220), .A2(W18034), .ZN(O5209));
  NOR2X1 G7353 (.A1(I1725), .A2(W4119), .ZN(W14253));
  NOR2X1 G7354 (.A1(W13324), .A2(W23224), .ZN(W30160));
  NOR2X1 G7355 (.A1(I1416), .A2(W6899), .ZN(W14251));
  NOR2X1 G7356 (.A1(W4929), .A2(W28088), .ZN(W30159));
  NOR2X1 G7357 (.A1(W22919), .A2(W30115), .ZN(W36576));
  NOR2X1 G7358 (.A1(W21145), .A2(W29981), .ZN(O5208));
  NOR2X1 G7359 (.A1(W8195), .A2(W16270), .ZN(W20615));
  NOR2X1 G7360 (.A1(W9618), .A2(W3515), .ZN(W14286));
  NOR2X1 G7361 (.A1(W7779), .A2(W518), .ZN(W20613));
  NOR2X1 G7362 (.A1(I1614), .A2(W16307), .ZN(O8459));
  NOR2X1 G7363 (.A1(W6942), .A2(W2480), .ZN(W14283));
  NOR2X1 G7364 (.A1(W420), .A2(W8131), .ZN(W14282));
  NOR2X1 G7365 (.A1(W13255), .A2(W4986), .ZN(W36543));
  NOR2X1 G7366 (.A1(W20624), .A2(I1934), .ZN(O8460));
  NOR2X1 G7367 (.A1(W2503), .A2(W2758), .ZN(W14279));
  NOR2X1 G7368 (.A1(W24717), .A2(W19833), .ZN(W30155));
  NOR2X1 G7369 (.A1(W2413), .A2(W15551), .ZN(O8463));
  NOR2X1 G7370 (.A1(W710), .A2(W7602), .ZN(W14275));
  NOR2X1 G7371 (.A1(W25049), .A2(W24182), .ZN(W30173));
  NOR2X1 G7372 (.A1(W10566), .A2(W2155), .ZN(W14272));
  NOR2X1 G7373 (.A1(W7584), .A2(W9776), .ZN(W14271));
  NOR2X1 G7374 (.A1(W14605), .A2(W27189), .ZN(O8469));
  NOR2X1 G7375 (.A1(W26455), .A2(W26037), .ZN(O8470));
  NOR2X1 G7376 (.A1(W5031), .A2(W5210), .ZN(W14214));
  NOR2X1 G7377 (.A1(I1478), .A2(W36417), .ZN(W36605));
  NOR2X1 G7378 (.A1(W2914), .A2(W13121), .ZN(W14221));
  NOR2X1 G7379 (.A1(W17738), .A2(W28319), .ZN(W36608));
  NOR2X1 G7380 (.A1(W12960), .A2(W17671), .ZN(W20639));
  NOR2X1 G7381 (.A1(W20550), .A2(I198), .ZN(W20640));
  NOR2X1 G7382 (.A1(W1473), .A2(W3064), .ZN(W14217));
  NOR2X1 G7383 (.A1(W35662), .A2(W17389), .ZN(O8502));
  NOR2X1 G7384 (.A1(W11941), .A2(W2292), .ZN(W14215));
  NOR2X1 G7385 (.A1(W9683), .A2(W3935), .ZN(W36602));
  NOR2X1 G7386 (.A1(W2391), .A2(W13756), .ZN(W14213));
  NOR2X1 G7387 (.A1(W6338), .A2(W13528), .ZN(W14212));
  NOR2X1 G7388 (.A1(W13691), .A2(W8884), .ZN(W20641));
  NOR2X1 G7389 (.A1(W12172), .A2(W17831), .ZN(O8506));
  NOR2X1 G7390 (.A1(W28497), .A2(W14951), .ZN(O8507));
  NOR2X1 G7391 (.A1(W27122), .A2(W12338), .ZN(O8509));
  NOR2X1 G7392 (.A1(W1864), .A2(W5956), .ZN(W14205));
  NOR2X1 G7393 (.A1(W128), .A2(W11184), .ZN(W14204));
  NOR2X1 G7394 (.A1(W950), .A2(W8641), .ZN(W20633));
  NOR2X1 G7395 (.A1(W9433), .A2(W11119), .ZN(W36582));
  NOR2X1 G7396 (.A1(W8357), .A2(W28256), .ZN(W30152));
  NOR2X1 G7397 (.A1(I1777), .A2(W14120), .ZN(W14243));
  NOR2X1 G7398 (.A1(W11892), .A2(W5933), .ZN(W14242));
  NOR2X1 G7399 (.A1(W33989), .A2(W10880), .ZN(O8488));
  NOR2X1 G7400 (.A1(W16678), .A2(W27544), .ZN(W30150));
  NOR2X1 G7401 (.A1(W9346), .A2(W28794), .ZN(O8489));
  NOR2X1 G7402 (.A1(W29391), .A2(W27726), .ZN(W36589));
  NOR2X1 G7403 (.A1(W10980), .A2(W12748), .ZN(W14124));
  NOR2X1 G7404 (.A1(I726), .A2(W10525), .ZN(W14235));
  NOR2X1 G7405 (.A1(W34033), .A2(W17440), .ZN(W36592));
  NOR2X1 G7406 (.A1(W30214), .A2(W27629), .ZN(W36595));
  NOR2X1 G7407 (.A1(W14336), .A2(W26403), .ZN(O8493));
  NOR2X1 G7408 (.A1(W13465), .A2(W14260), .ZN(W36599));
  NOR2X1 G7409 (.A1(W3392), .A2(W8053), .ZN(O8494));
  NOR2X1 G7410 (.A1(W11805), .A2(W5084), .ZN(O845));
  NOR2X1 G7411 (.A1(W2747), .A2(I1030), .ZN(W14006));
  NOR2X1 G7412 (.A1(W16053), .A2(W2947), .ZN(O5173));
  NOR2X1 G7413 (.A1(W10708), .A2(W13173), .ZN(O816));
  NOR2X1 G7414 (.A1(W12292), .A2(W1484), .ZN(W14012));
  NOR2X1 G7415 (.A1(W13547), .A2(W13900), .ZN(W14011));
  NOR2X1 G7416 (.A1(W13612), .A2(W22433), .ZN(W36807));
  NOR2X1 G7417 (.A1(I331), .A2(W4163), .ZN(O815));
  NOR2X1 G7418 (.A1(W16119), .A2(W2018), .ZN(W20716));
  NOR2X1 G7419 (.A1(W26705), .A2(W23843), .ZN(W36810));
  NOR2X1 G7420 (.A1(W2517), .A2(W726), .ZN(W14015));
  NOR2X1 G7421 (.A1(W29621), .A2(W26311), .ZN(W36814));
  NOR2X1 G7422 (.A1(W11635), .A2(W4715), .ZN(W14004));
  NOR2X1 G7423 (.A1(W23288), .A2(W18733), .ZN(O5172));
  NOR2X1 G7424 (.A1(W27595), .A2(W17963), .ZN(W30053));
  NOR2X1 G7425 (.A1(W647), .A2(W3881), .ZN(W14000));
  NOR2X1 G7426 (.A1(W9400), .A2(W3550), .ZN(W20720));
  NOR2X1 G7427 (.A1(W5875), .A2(W21407), .ZN(O8615));
  NOR2X1 G7428 (.A1(W3216), .A2(W10439), .ZN(W13997));
  NOR2X1 G7429 (.A1(W9681), .A2(W5608), .ZN(O2063));
  NOR2X1 G7430 (.A1(W24594), .A2(W2236), .ZN(W36791));
  NOR2X1 G7431 (.A1(W3706), .A2(W4075), .ZN(W14032));
  NOR2X1 G7432 (.A1(W13692), .A2(I839), .ZN(W14031));
  NOR2X1 G7433 (.A1(W11739), .A2(W13487), .ZN(W14030));
  NOR2X1 G7434 (.A1(W9938), .A2(W7524), .ZN(W30063));
  NOR2X1 G7435 (.A1(W6364), .A2(W8179), .ZN(W14028));
  NOR2X1 G7436 (.A1(W1903), .A2(W2791), .ZN(W14027));
  NOR2X1 G7437 (.A1(W8451), .A2(W7912), .ZN(W14026));
  NOR2X1 G7438 (.A1(W17496), .A2(W6893), .ZN(W30050));
  NOR2X1 G7439 (.A1(W5095), .A2(W19428), .ZN(W36796));
  NOR2X1 G7440 (.A1(W12036), .A2(W8497), .ZN(W20712));
  NOR2X1 G7441 (.A1(W828), .A2(W3994), .ZN(W14020));
  NOR2X1 G7442 (.A1(W12738), .A2(W2041), .ZN(W14019));
  NOR2X1 G7443 (.A1(W30180), .A2(W25711), .ZN(O8604));
  NOR2X1 G7444 (.A1(W3019), .A2(W16137), .ZN(O8605));
  NOR2X1 G7445 (.A1(W7134), .A2(W933), .ZN(W20714));
  NOR2X1 G7446 (.A1(W12994), .A2(W9207), .ZN(W13968));
  NOR2X1 G7447 (.A1(W7537), .A2(W423), .ZN(W13976));
  NOR2X1 G7448 (.A1(W22820), .A2(W6082), .ZN(O8630));
  NOR2X1 G7449 (.A1(I393), .A2(W13098), .ZN(W13974));
  NOR2X1 G7450 (.A1(W20326), .A2(W496), .ZN(W30046));
  NOR2X1 G7451 (.A1(W9818), .A2(W828), .ZN(W13972));
  NOR2X1 G7452 (.A1(W28931), .A2(W34251), .ZN(O8631));
  NOR2X1 G7453 (.A1(W8659), .A2(W11447), .ZN(O812));
  NOR2X1 G7454 (.A1(W2487), .A2(W6601), .ZN(W36848));
  NOR2X1 G7455 (.A1(W20036), .A2(W6668), .ZN(W36841));
  NOR2X1 G7456 (.A1(W3466), .A2(W7588), .ZN(W13967));
  NOR2X1 G7457 (.A1(W2479), .A2(W3461), .ZN(W13966));
  NOR2X1 G7458 (.A1(W1003), .A2(W3628), .ZN(W13965));
  NOR2X1 G7459 (.A1(W881), .A2(I705), .ZN(O811));
  NOR2X1 G7460 (.A1(W1650), .A2(W28699), .ZN(W36849));
  NOR2X1 G7461 (.A1(I694), .A2(W16457), .ZN(W36850));
  NOR2X1 G7462 (.A1(W16078), .A2(W29844), .ZN(O8632));
  NOR2X1 G7463 (.A1(W6186), .A2(W9894), .ZN(O8633));
  NOR2X1 G7464 (.A1(W9402), .A2(W549), .ZN(W13986));
  NOR2X1 G7465 (.A1(W2899), .A2(I337), .ZN(W13995));
  NOR2X1 G7466 (.A1(W2419), .A2(W636), .ZN(W13994));
  NOR2X1 G7467 (.A1(W11801), .A2(W18952), .ZN(W36825));
  NOR2X1 G7468 (.A1(W25025), .A2(W10431), .ZN(O8619));
  NOR2X1 G7469 (.A1(W18580), .A2(W18288), .ZN(W20722));
  NOR2X1 G7470 (.A1(W10800), .A2(W12243), .ZN(W13989));
  NOR2X1 G7471 (.A1(W11893), .A2(W10224), .ZN(W13988));
  NOR2X1 G7472 (.A1(W23717), .A2(W36216), .ZN(O8621));
  NOR2X1 G7473 (.A1(W6551), .A2(W5959), .ZN(W30065));
  NOR2X1 G7474 (.A1(W702), .A2(W20912), .ZN(O8623));
  NOR2X1 G7475 (.A1(W12393), .A2(W12360), .ZN(W13984));
  NOR2X1 G7476 (.A1(W20160), .A2(W32507), .ZN(O8626));
  NOR2X1 G7477 (.A1(W6524), .A2(I474), .ZN(W13982));
  NOR2X1 G7478 (.A1(W7064), .A2(I442), .ZN(W13981));
  NOR2X1 G7479 (.A1(W6216), .A2(W6159), .ZN(O8628));
  NOR2X1 G7480 (.A1(W9084), .A2(W1874), .ZN(W13979));
  NOR2X1 G7481 (.A1(W28729), .A2(W25476), .ZN(O8566));
  NOR2X1 G7482 (.A1(W18010), .A2(W15587), .ZN(W20678));
  NOR2X1 G7483 (.A1(W23820), .A2(W5310), .ZN(W30103));
  NOR2X1 G7484 (.A1(W10223), .A2(W2597), .ZN(W14101));
  NOR2X1 G7485 (.A1(W12506), .A2(I1287), .ZN(W14100));
  NOR2X1 G7486 (.A1(I1253), .A2(W13414), .ZN(O826));
  NOR2X1 G7487 (.A1(W8505), .A2(W1451), .ZN(O825));
  NOR2X1 G7488 (.A1(W3271), .A2(W12407), .ZN(W14096));
  NOR2X1 G7489 (.A1(W4189), .A2(W11394), .ZN(W14095));
  NOR2X1 G7490 (.A1(W10052), .A2(W8785), .ZN(W14104));
  NOR2X1 G7491 (.A1(W10932), .A2(W959), .ZN(O2055));
  NOR2X1 G7492 (.A1(W26261), .A2(W13032), .ZN(W36735));
  NOR2X1 G7493 (.A1(W28011), .A2(W30818), .ZN(W36736));
  NOR2X1 G7494 (.A1(W1058), .A2(W7265), .ZN(W36737));
  NOR2X1 G7495 (.A1(W32771), .A2(W20802), .ZN(W36738));
  NOR2X1 G7496 (.A1(I1200), .A2(W3097), .ZN(W14087));
  NOR2X1 G7497 (.A1(W12538), .A2(W894), .ZN(O2056));
  NOR2X1 G7498 (.A1(W7986), .A2(W19220), .ZN(W30094));
  NOR2X1 G7499 (.A1(W343), .A2(W8513), .ZN(W14113));
  NOR2X1 G7500 (.A1(W32164), .A2(W952), .ZN(W36704));
  NOR2X1 G7501 (.A1(W13199), .A2(W13312), .ZN(W14122));
  NOR2X1 G7502 (.A1(W20872), .A2(W29240), .ZN(W30109));
  NOR2X1 G7503 (.A1(W8197), .A2(W10769), .ZN(O8555));
  NOR2X1 G7504 (.A1(I603), .A2(W4829), .ZN(O2054));
  NOR2X1 G7505 (.A1(W29579), .A2(W35855), .ZN(O8556));
  NOR2X1 G7506 (.A1(W22088), .A2(W13771), .ZN(O5192));
  NOR2X1 G7507 (.A1(W18653), .A2(W28676), .ZN(O8558));
  NOR2X1 G7508 (.A1(W7971), .A2(W3705), .ZN(W14083));
  NOR2X1 G7509 (.A1(W9874), .A2(W2824), .ZN(W14112));
  NOR2X1 G7510 (.A1(W5032), .A2(W9152), .ZN(W14111));
  NOR2X1 G7511 (.A1(W1900), .A2(W36642), .ZN(W36716));
  NOR2X1 G7512 (.A1(W12157), .A2(W15161), .ZN(W20677));
  NOR2X1 G7513 (.A1(W36186), .A2(W9073), .ZN(O8561));
  NOR2X1 G7514 (.A1(I1952), .A2(W13913), .ZN(W14106));
  NOR2X1 G7515 (.A1(W28584), .A2(W5190), .ZN(W36721));
  NOR2X1 G7516 (.A1(W569), .A2(W13749), .ZN(W20704));
  NOR2X1 G7517 (.A1(W18154), .A2(W20928), .ZN(O8589));
  NOR2X1 G7518 (.A1(W2856), .A2(W3906), .ZN(O820));
  NOR2X1 G7519 (.A1(W8102), .A2(W6476), .ZN(W14050));
  NOR2X1 G7520 (.A1(W8562), .A2(W12858), .ZN(W14049));
  NOR2X1 G7521 (.A1(W6038), .A2(W879), .ZN(W20702));
  NOR2X1 G7522 (.A1(W327), .A2(W4831), .ZN(W14047));
  NOR2X1 G7523 (.A1(W21720), .A2(W34877), .ZN(W36778));
  NOR2X1 G7524 (.A1(W17340), .A2(W8591), .ZN(W20703));
  NOR2X1 G7525 (.A1(W22565), .A2(W35939), .ZN(W36774));
  NOR2X1 G7526 (.A1(W2258), .A2(I558), .ZN(W14043));
  NOR2X1 G7527 (.A1(W4706), .A2(W16483), .ZN(O8592));
  NOR2X1 G7528 (.A1(W17880), .A2(W20909), .ZN(O8593));
  NOR2X1 G7529 (.A1(W8737), .A2(W7873), .ZN(W20705));
  NOR2X1 G7530 (.A1(W24061), .A2(W26054), .ZN(O8595));
  NOR2X1 G7531 (.A1(W13753), .A2(W2749), .ZN(O819));
  NOR2X1 G7532 (.A1(W17045), .A2(W28087), .ZN(W30068));
  NOR2X1 G7533 (.A1(W5644), .A2(W5221), .ZN(W14036));
  NOR2X1 G7534 (.A1(W2857), .A2(W34167), .ZN(W36754));
  NOR2X1 G7535 (.A1(W7844), .A2(W11364), .ZN(O2058));
  NOR2X1 G7536 (.A1(W35), .A2(W6383), .ZN(W14077));
  NOR2X1 G7537 (.A1(W3099), .A2(W11140), .ZN(W14076));
  NOR2X1 G7538 (.A1(W19202), .A2(W12400), .ZN(O5185));
  NOR2X1 G7539 (.A1(W9814), .A2(W24465), .ZN(O8577));
  NOR2X1 G7540 (.A1(W2943), .A2(W4581), .ZN(W14073));
  NOR2X1 G7541 (.A1(W1943), .A2(W4797), .ZN(W14072));
  NOR2X1 G7542 (.A1(I928), .A2(W4058), .ZN(W14071));
  NOR2X1 G7543 (.A1(I1018), .A2(W9787), .ZN(W14287));
  NOR2X1 G7544 (.A1(W27090), .A2(W22581), .ZN(W36758));
  NOR2X1 G7545 (.A1(I1863), .A2(W7524), .ZN(W36760));
  NOR2X1 G7546 (.A1(W7107), .A2(W1120), .ZN(W14065));
  NOR2X1 G7547 (.A1(W7040), .A2(W11111), .ZN(O8586));
  NOR2X1 G7548 (.A1(W27229), .A2(W27164), .ZN(O5179));
  NOR2X1 G7549 (.A1(W1451), .A2(W10852), .ZN(W14058));
  NOR2X1 G7550 (.A1(W5044), .A2(W9593), .ZN(W14055));
  NOR2X1 G7551 (.A1(W13646), .A2(W8280), .ZN(W14494));
  NOR2X1 G7552 (.A1(W4256), .A2(W1657), .ZN(O878));
  NOR2X1 G7553 (.A1(W3491), .A2(W9441), .ZN(W14502));
  NOR2X1 G7554 (.A1(W2773), .A2(W11841), .ZN(O8318));
  NOR2X1 G7555 (.A1(W11140), .A2(W12780), .ZN(W14500));
  NOR2X1 G7556 (.A1(I1854), .A2(W4286), .ZN(W14498));
  NOR2X1 G7557 (.A1(W21717), .A2(W22291), .ZN(O8320));
  NOR2X1 G7558 (.A1(W3766), .A2(W33694), .ZN(O8322));
  NOR2X1 G7559 (.A1(W27929), .A2(W31348), .ZN(O8323));
  NOR2X1 G7560 (.A1(W6801), .A2(W25917), .ZN(O8315));
  NOR2X1 G7561 (.A1(W11585), .A2(W10900), .ZN(O8324));
  NOR2X1 G7562 (.A1(W16342), .A2(W10567), .ZN(O8326));
  NOR2X1 G7563 (.A1(I1638), .A2(W19561), .ZN(W20548));
  NOR2X1 G7564 (.A1(W7610), .A2(W10521), .ZN(W14489));
  NOR2X1 G7565 (.A1(W388), .A2(W14747), .ZN(O8329));
  NOR2X1 G7566 (.A1(W10674), .A2(W12489), .ZN(W14487));
  NOR2X1 G7567 (.A1(W10843), .A2(W17863), .ZN(O8331));
  NOR2X1 G7568 (.A1(W30086), .A2(W36067), .ZN(W36325));
  NOR2X1 G7569 (.A1(W6784), .A2(W4716), .ZN(W14513));
  NOR2X1 G7570 (.A1(W22252), .A2(W5368), .ZN(O8303));
  NOR2X1 G7571 (.A1(W4296), .A2(W13910), .ZN(W14524));
  NOR2X1 G7572 (.A1(W8078), .A2(W5315), .ZN(W14523));
  NOR2X1 G7573 (.A1(W34592), .A2(W32397), .ZN(O8308));
  NOR2X1 G7574 (.A1(W201), .A2(W9193), .ZN(W14520));
  NOR2X1 G7575 (.A1(W11833), .A2(W29171), .ZN(O5255));
  NOR2X1 G7576 (.A1(W9360), .A2(W9337), .ZN(W14516));
  NOR2X1 G7577 (.A1(I393), .A2(W10686), .ZN(W30249));
  NOR2X1 G7578 (.A1(W10397), .A2(W511), .ZN(O2027));
  NOR2X1 G7579 (.A1(I1003), .A2(W3765), .ZN(W14512));
  NOR2X1 G7580 (.A1(W2378), .A2(I752), .ZN(W14511));
  NOR2X1 G7581 (.A1(W5102), .A2(W2574), .ZN(O5253));
  NOR2X1 G7582 (.A1(W12617), .A2(W2116), .ZN(W14509));
  NOR2X1 G7583 (.A1(W12063), .A2(I1662), .ZN(W14508));
  NOR2X1 G7584 (.A1(I770), .A2(W8768), .ZN(O5252));
  NOR2X1 G7585 (.A1(W12042), .A2(W24086), .ZN(O5251));
  NOR2X1 G7586 (.A1(W29207), .A2(W21698), .ZN(O5246));
  NOR2X1 G7587 (.A1(W12549), .A2(I572), .ZN(W36344));
  NOR2X1 G7588 (.A1(W17207), .A2(W17910), .ZN(W20552));
  NOR2X1 G7589 (.A1(W26973), .A2(W10085), .ZN(W30238));
  NOR2X1 G7590 (.A1(W25350), .A2(W20882), .ZN(W36347));
  NOR2X1 G7591 (.A1(W10088), .A2(W2381), .ZN(W14462));
  NOR2X1 G7592 (.A1(W20002), .A2(W4202), .ZN(O8340));
  NOR2X1 G7593 (.A1(W2254), .A2(W13696), .ZN(W36351));
  NOR2X1 G7594 (.A1(W3818), .A2(W2739), .ZN(O8341));
  NOR2X1 G7595 (.A1(W29209), .A2(W17732), .ZN(O8337));
  NOR2X1 G7596 (.A1(W13861), .A2(I68), .ZN(W14457));
  NOR2X1 G7597 (.A1(W16167), .A2(W23931), .ZN(W36355));
  NOR2X1 G7598 (.A1(W2091), .A2(W33319), .ZN(O8343));
  NOR2X1 G7599 (.A1(W2777), .A2(W17444), .ZN(O5245));
  NOR2X1 G7600 (.A1(W17603), .A2(I1959), .ZN(W20556));
  NOR2X1 G7601 (.A1(W1398), .A2(W31299), .ZN(W36361));
  NOR2X1 G7602 (.A1(W11651), .A2(W3871), .ZN(W14450));
  NOR2X1 G7603 (.A1(W11470), .A2(W608), .ZN(W14448));
  NOR2X1 G7604 (.A1(W32906), .A2(W9508), .ZN(W36335));
  NOR2X1 G7605 (.A1(W911), .A2(W11719), .ZN(W14483));
  NOR2X1 G7606 (.A1(W34877), .A2(W2280), .ZN(W36328));
  NOR2X1 G7607 (.A1(W10302), .A2(I1534), .ZN(O5248));
  NOR2X1 G7608 (.A1(W369), .A2(W6568), .ZN(W14480));
  NOR2X1 G7609 (.A1(W5545), .A2(W27717), .ZN(O8332));
  NOR2X1 G7610 (.A1(W6831), .A2(W26265), .ZN(W36332));
  NOR2X1 G7611 (.A1(W18140), .A2(I570), .ZN(O8334));
  NOR2X1 G7612 (.A1(W4492), .A2(W35369), .ZN(O8335));
  NOR2X1 G7613 (.A1(W16372), .A2(W15074), .ZN(W20535));
  NOR2X1 G7614 (.A1(W14791), .A2(W21561), .ZN(O8336));
  NOR2X1 G7615 (.A1(W26502), .A2(W7420), .ZN(W36340));
  NOR2X1 G7616 (.A1(W23600), .A2(W36135), .ZN(W36341));
  NOR2X1 G7617 (.A1(W4694), .A2(W1440), .ZN(W14471));
  NOR2X1 G7618 (.A1(W8132), .A2(W12185), .ZN(W14470));
  NOR2X1 G7619 (.A1(W11390), .A2(W54), .ZN(W14469));
  NOR2X1 G7620 (.A1(W725), .A2(W8438), .ZN(W30239));
  NOR2X1 G7621 (.A1(W12427), .A2(W14205), .ZN(W14574));
  NOR2X1 G7622 (.A1(W15246), .A2(W1460), .ZN(W20519));
  NOR2X1 G7623 (.A1(W4987), .A2(W1044), .ZN(W14581));
  NOR2X1 G7624 (.A1(W9304), .A2(I1427), .ZN(O885));
  NOR2X1 G7625 (.A1(W8686), .A2(W2286), .ZN(W14579));
  NOR2X1 G7626 (.A1(W12122), .A2(W15227), .ZN(O2022));
  NOR2X1 G7627 (.A1(W27127), .A2(W34092), .ZN(O8277));
  NOR2X1 G7628 (.A1(W7721), .A2(W4396), .ZN(W14576));
  NOR2X1 G7629 (.A1(W8974), .A2(W4592), .ZN(W14575));
  NOR2X1 G7630 (.A1(W5129), .A2(W6049), .ZN(O8275));
  NOR2X1 G7631 (.A1(W14516), .A2(W4614), .ZN(W36239));
  NOR2X1 G7632 (.A1(W11693), .A2(W19568), .ZN(W20521));
  NOR2X1 G7633 (.A1(W1434), .A2(W8434), .ZN(W14571));
  NOR2X1 G7634 (.A1(W11421), .A2(I414), .ZN(W36241));
  NOR2X1 G7635 (.A1(W29053), .A2(W32397), .ZN(O8280));
  NOR2X1 G7636 (.A1(W19067), .A2(W2967), .ZN(W20522));
  NOR2X1 G7637 (.A1(W7456), .A2(W3342), .ZN(W14567));
  NOR2X1 G7638 (.A1(W14209), .A2(W10644), .ZN(W14566));
  NOR2X1 G7639 (.A1(W1155), .A2(W11867), .ZN(W14591));
  NOR2X1 G7640 (.A1(W6844), .A2(I1599), .ZN(W14599));
  NOR2X1 G7641 (.A1(W12876), .A2(W547), .ZN(W14598));
  NOR2X1 G7642 (.A1(W31822), .A2(W23916), .ZN(W36215));
  NOR2X1 G7643 (.A1(W5011), .A2(W29727), .ZN(O8264));
  NOR2X1 G7644 (.A1(W30360), .A2(W17232), .ZN(O8265));
  NOR2X1 G7645 (.A1(W7534), .A2(W19813), .ZN(W36220));
  NOR2X1 G7646 (.A1(W13220), .A2(W19762), .ZN(O8266));
  NOR2X1 G7647 (.A1(I549), .A2(W4329), .ZN(O887));
  NOR2X1 G7648 (.A1(W7349), .A2(W10638), .ZN(O2023));
  NOR2X1 G7649 (.A1(W20923), .A2(W6868), .ZN(W36222));
  NOR2X1 G7650 (.A1(W14880), .A2(W17004), .ZN(O2021));
  NOR2X1 G7651 (.A1(W34192), .A2(W13617), .ZN(O8270));
  NOR2X1 G7652 (.A1(W12345), .A2(W18788), .ZN(W36229));
  NOR2X1 G7653 (.A1(W28371), .A2(W19887), .ZN(O5262));
  NOR2X1 G7654 (.A1(W9948), .A2(W24420), .ZN(O8274));
  NOR2X1 G7655 (.A1(W29011), .A2(W26146), .ZN(W36233));
  NOR2X1 G7656 (.A1(W31494), .A2(W14080), .ZN(W36274));
  NOR2X1 G7657 (.A1(I1134), .A2(W8443), .ZN(W14544));
  NOR2X1 G7658 (.A1(W571), .A2(W27647), .ZN(W36266));
  NOR2X1 G7659 (.A1(I890), .A2(W3222), .ZN(W14542));
  NOR2X1 G7660 (.A1(W16002), .A2(W14451), .ZN(W30263));
  NOR2X1 G7661 (.A1(W19173), .A2(W3650), .ZN(W20530));
  NOR2X1 G7662 (.A1(W17453), .A2(W7305), .ZN(W20531));
  NOR2X1 G7663 (.A1(W4445), .A2(W14415), .ZN(W14538));
  NOR2X1 G7664 (.A1(W7717), .A2(W13290), .ZN(W14537));
  NOR2X1 G7665 (.A1(W27393), .A2(W17123), .ZN(O5259));
  NOR2X1 G7666 (.A1(W21979), .A2(W24726), .ZN(W36278));
  NOR2X1 G7667 (.A1(W28508), .A2(W12951), .ZN(W36279));
  NOR2X1 G7668 (.A1(W1332), .A2(W6302), .ZN(O8298));
  NOR2X1 G7669 (.A1(W23959), .A2(W6620), .ZN(W30262));
  NOR2X1 G7670 (.A1(W6971), .A2(W24946), .ZN(W36282));
  NOR2X1 G7671 (.A1(W7462), .A2(W10922), .ZN(W14530));
  NOR2X1 G7672 (.A1(W9363), .A2(W11626), .ZN(W36284));
  NOR2X1 G7673 (.A1(W17010), .A2(W26331), .ZN(W30259));
  NOR2X1 G7674 (.A1(W20492), .A2(W3624), .ZN(W36254));
  NOR2X1 G7675 (.A1(W2435), .A2(W13714), .ZN(W14564));
  NOR2X1 G7676 (.A1(I1042), .A2(I1684), .ZN(W14563));
  NOR2X1 G7677 (.A1(W11203), .A2(W13924), .ZN(W14562));
  NOR2X1 G7678 (.A1(W35807), .A2(W27927), .ZN(W36249));
  NOR2X1 G7679 (.A1(W10666), .A2(W21159), .ZN(O8282));
  NOR2X1 G7680 (.A1(W28293), .A2(W16209), .ZN(O5261));
  NOR2X1 G7681 (.A1(W11583), .A2(W974), .ZN(W14558));
  NOR2X1 G7682 (.A1(W1806), .A2(W9169), .ZN(W14557));
  NOR2X1 G7683 (.A1(W19376), .A2(W8544), .ZN(W36365));
  NOR2X1 G7684 (.A1(W995), .A2(W8956), .ZN(W14553));
  NOR2X1 G7685 (.A1(W19421), .A2(W34400), .ZN(O8285));
  NOR2X1 G7686 (.A1(W24593), .A2(W20843), .ZN(O8286));
  NOR2X1 G7687 (.A1(W31444), .A2(W11248), .ZN(O8287));
  NOR2X1 G7688 (.A1(W25553), .A2(W4254), .ZN(W36260));
  NOR2X1 G7689 (.A1(W3013), .A2(W6586), .ZN(W14548));
  NOR2X1 G7690 (.A1(W8549), .A2(W4674), .ZN(W36263));
  NOR2X1 G7691 (.A1(W32232), .A2(W23403), .ZN(O8432));
  NOR2X1 G7692 (.A1(W12877), .A2(W7903), .ZN(W36484));
  NOR2X1 G7693 (.A1(W7359), .A2(W2152), .ZN(W14346));
  NOR2X1 G7694 (.A1(W15945), .A2(W29665), .ZN(W36485));
  NOR2X1 G7695 (.A1(W15296), .A2(W13917), .ZN(W30194));
  NOR2X1 G7696 (.A1(I392), .A2(I1512), .ZN(O855));
  NOR2X1 G7697 (.A1(W17947), .A2(W35235), .ZN(W36487));
  NOR2X1 G7698 (.A1(W15542), .A2(W9668), .ZN(W36488));
  NOR2X1 G7699 (.A1(W13430), .A2(W8439), .ZN(O5224));
  NOR2X1 G7700 (.A1(W8704), .A2(W5577), .ZN(O8424));
  NOR2X1 G7701 (.A1(W24818), .A2(W6863), .ZN(O5223));
  NOR2X1 G7702 (.A1(W6586), .A2(W8260), .ZN(W14336));
  NOR2X1 G7703 (.A1(W32209), .A2(W7057), .ZN(W36504));
  NOR2X1 G7704 (.A1(W10174), .A2(W34488), .ZN(W36505));
  NOR2X1 G7705 (.A1(W10892), .A2(W10833), .ZN(W14330));
  NOR2X1 G7706 (.A1(W7097), .A2(W1754), .ZN(W14329));
  NOR2X1 G7707 (.A1(W12453), .A2(I1888), .ZN(W14328));
  NOR2X1 G7708 (.A1(W30980), .A2(W3530), .ZN(W36506));
  NOR2X1 G7709 (.A1(W10817), .A2(W18567), .ZN(O5227));
  NOR2X1 G7710 (.A1(I1305), .A2(W11464), .ZN(O857));
  NOR2X1 G7711 (.A1(W27278), .A2(W30024), .ZN(O8411));
  NOR2X1 G7712 (.A1(W4046), .A2(W20297), .ZN(O8412));
  NOR2X1 G7713 (.A1(W4270), .A2(W3723), .ZN(W14363));
  NOR2X1 G7714 (.A1(W2520), .A2(W774), .ZN(W14362));
  NOR2X1 G7715 (.A1(W9757), .A2(W12400), .ZN(O8413));
  NOR2X1 G7716 (.A1(W22850), .A2(W22034), .ZN(W36467));
  NOR2X1 G7717 (.A1(W24690), .A2(W24695), .ZN(W36469));
  NOR2X1 G7718 (.A1(W4957), .A2(I661), .ZN(W14326));
  NOR2X1 G7719 (.A1(W12155), .A2(W13611), .ZN(W20593));
  NOR2X1 G7720 (.A1(W18112), .A2(W16049), .ZN(W20594));
  NOR2X1 G7721 (.A1(W14174), .A2(I1409), .ZN(W30199));
  NOR2X1 G7722 (.A1(W29047), .A2(W16172), .ZN(O8421));
  NOR2X1 G7723 (.A1(W3440), .A2(W10521), .ZN(W14353));
  NOR2X1 G7724 (.A1(W2019), .A2(W6508), .ZN(W14352));
  NOR2X1 G7725 (.A1(W10428), .A2(W9064), .ZN(W14350));
  NOR2X1 G7726 (.A1(W27239), .A2(W25715), .ZN(W30178));
  NOR2X1 G7727 (.A1(W14048), .A2(W8354), .ZN(W14307));
  NOR2X1 G7728 (.A1(W3463), .A2(W23766), .ZN(O8444));
  NOR2X1 G7729 (.A1(I402), .A2(W7735), .ZN(W14305));
  NOR2X1 G7730 (.A1(W8511), .A2(W3179), .ZN(W14304));
  NOR2X1 G7731 (.A1(W32349), .A2(W17911), .ZN(W36518));
  NOR2X1 G7732 (.A1(W13365), .A2(W15944), .ZN(W20610));
  NOR2X1 G7733 (.A1(W31812), .A2(W20889), .ZN(O8450));
  NOR2X1 G7734 (.A1(W2113), .A2(W30304), .ZN(O8453));
  NOR2X1 G7735 (.A1(I85), .A2(W8409), .ZN(W14308));
  NOR2X1 G7736 (.A1(W1475), .A2(W10604), .ZN(W36533));
  NOR2X1 G7737 (.A1(W11950), .A2(W8235), .ZN(O853));
  NOR2X1 G7738 (.A1(W15603), .A2(W633), .ZN(O8456));
  NOR2X1 G7739 (.A1(W4130), .A2(W10547), .ZN(W14293));
  NOR2X1 G7740 (.A1(W2276), .A2(I326), .ZN(W14292));
  NOR2X1 G7741 (.A1(W12252), .A2(W2198), .ZN(W36535));
  NOR2X1 G7742 (.A1(W28183), .A2(W23770), .ZN(W36537));
  NOR2X1 G7743 (.A1(W6642), .A2(W20176), .ZN(O8458));
  NOR2X1 G7744 (.A1(I895), .A2(I235), .ZN(W14317));
  NOR2X1 G7745 (.A1(W9989), .A2(W11981), .ZN(W14325));
  NOR2X1 G7746 (.A1(I1697), .A2(W6664), .ZN(W14324));
  NOR2X1 G7747 (.A1(W10847), .A2(I116), .ZN(W14323));
  NOR2X1 G7748 (.A1(W1865), .A2(W22852), .ZN(O8437));
  NOR2X1 G7749 (.A1(W684), .A2(W264), .ZN(W14321));
  NOR2X1 G7750 (.A1(W1761), .A2(W4636), .ZN(W14320));
  NOR2X1 G7751 (.A1(W12400), .A2(W4087), .ZN(W14319));
  NOR2X1 G7752 (.A1(W17758), .A2(W24776), .ZN(O8438));
  NOR2X1 G7753 (.A1(W22686), .A2(W25547), .ZN(O8410));
  NOR2X1 G7754 (.A1(W27426), .A2(W6786), .ZN(W36509));
  NOR2X1 G7755 (.A1(W14371), .A2(W22078), .ZN(O5220));
  NOR2X1 G7756 (.A1(W7554), .A2(W6394), .ZN(W14314));
  NOR2X1 G7757 (.A1(W10768), .A2(W9167), .ZN(W14313));
  NOR2X1 G7758 (.A1(W14293), .A2(W14627), .ZN(O5219));
  NOR2X1 G7759 (.A1(W35465), .A2(W12051), .ZN(W36514));
  NOR2X1 G7760 (.A1(W9222), .A2(W9607), .ZN(W14309));
  NOR2X1 G7761 (.A1(W15523), .A2(W19830), .ZN(W30215));
  NOR2X1 G7762 (.A1(W3934), .A2(W2790), .ZN(W14426));
  NOR2X1 G7763 (.A1(W7430), .A2(W12880), .ZN(W30221));
  NOR2X1 G7764 (.A1(W15359), .A2(W25078), .ZN(O8371));
  NOR2X1 G7765 (.A1(W12773), .A2(W16156), .ZN(O5238));
  NOR2X1 G7766 (.A1(W8126), .A2(W9353), .ZN(W14421));
  NOR2X1 G7767 (.A1(I493), .A2(W1182), .ZN(W14420));
  NOR2X1 G7768 (.A1(W23636), .A2(W15879), .ZN(W36397));
  NOR2X1 G7769 (.A1(W14382), .A2(W13137), .ZN(O8375));
  NOR2X1 G7770 (.A1(W6119), .A2(W563), .ZN(W14427));
  NOR2X1 G7771 (.A1(W7399), .A2(W9336), .ZN(W14414));
  NOR2X1 G7772 (.A1(W1629), .A2(W3140), .ZN(W14413));
  NOR2X1 G7773 (.A1(W20140), .A2(W25530), .ZN(O8376));
  NOR2X1 G7774 (.A1(W8389), .A2(W3613), .ZN(W20575));
  NOR2X1 G7775 (.A1(W30139), .A2(W25160), .ZN(O5235));
  NOR2X1 G7776 (.A1(W20515), .A2(W377), .ZN(W20577));
  NOR2X1 G7777 (.A1(W1998), .A2(I259), .ZN(W20578));
  NOR2X1 G7778 (.A1(W28734), .A2(W14347), .ZN(W36412));
  NOR2X1 G7779 (.A1(W2102), .A2(W2539), .ZN(W14437));
  NOR2X1 G7780 (.A1(W15594), .A2(W24638), .ZN(W30231));
  NOR2X1 G7781 (.A1(W27326), .A2(W28980), .ZN(W30230));
  NOR2X1 G7782 (.A1(I559), .A2(W20153), .ZN(O8354));
  NOR2X1 G7783 (.A1(W35999), .A2(W2167), .ZN(W36372));
  NOR2X1 G7784 (.A1(W5202), .A2(W2196), .ZN(W14441));
  NOR2X1 G7785 (.A1(W8698), .A2(W28243), .ZN(O8359));
  NOR2X1 G7786 (.A1(W14813), .A2(W19895), .ZN(W20562));
  NOR2X1 G7787 (.A1(W6273), .A2(W12642), .ZN(W20563));
  NOR2X1 G7788 (.A1(W10257), .A2(I29), .ZN(O2037));
  NOR2X1 G7789 (.A1(W1107), .A2(W355), .ZN(W36381));
  NOR2X1 G7790 (.A1(W10776), .A2(W13493), .ZN(O8363));
  NOR2X1 G7791 (.A1(W28425), .A2(W7888), .ZN(O5242));
  NOR2X1 G7792 (.A1(W9140), .A2(W12350), .ZN(W14433));
  NOR2X1 G7793 (.A1(W5889), .A2(W165), .ZN(W14432));
  NOR2X1 G7794 (.A1(W11612), .A2(I1763), .ZN(W14430));
  NOR2X1 G7795 (.A1(W14697), .A2(W7870), .ZN(W30224));
  NOR2X1 G7796 (.A1(W34768), .A2(W9136), .ZN(O8406));
  NOR2X1 G7797 (.A1(W36089), .A2(W17159), .ZN(O8398));
  NOR2X1 G7798 (.A1(W9143), .A2(W15914), .ZN(O2039));
  NOR2X1 G7799 (.A1(W32529), .A2(W8756), .ZN(O8400));
  NOR2X1 G7800 (.A1(W14961), .A2(W5745), .ZN(O8403));
  NOR2X1 G7801 (.A1(W24859), .A2(W9208), .ZN(O8404));
  NOR2X1 G7802 (.A1(W8872), .A2(W8980), .ZN(W14380));
  NOR2X1 G7803 (.A1(W23294), .A2(W28354), .ZN(W36451));
  NOR2X1 G7804 (.A1(W4544), .A2(W9520), .ZN(W20587));
  NOR2X1 G7805 (.A1(W26257), .A2(I454), .ZN(W36435));
  NOR2X1 G7806 (.A1(W5997), .A2(W12457), .ZN(W14376));
  NOR2X1 G7807 (.A1(W3594), .A2(W19539), .ZN(O5229));
  NOR2X1 G7808 (.A1(W1621), .A2(W19387), .ZN(W30203));
  NOR2X1 G7809 (.A1(W13059), .A2(W12134), .ZN(W14372));
  NOR2X1 G7810 (.A1(W251), .A2(W1806), .ZN(W14371));
  NOR2X1 G7811 (.A1(W9322), .A2(W11930), .ZN(O8409));
  NOR2X1 G7812 (.A1(W8174), .A2(W13831), .ZN(O859));
  NOR2X1 G7813 (.A1(W10908), .A2(I641), .ZN(O865));
  NOR2X1 G7814 (.A1(W6747), .A2(I648), .ZN(O866));
  NOR2X1 G7815 (.A1(W2361), .A2(W11095), .ZN(W14403));
  NOR2X1 G7816 (.A1(I206), .A2(W360), .ZN(W14402));
  NOR2X1 G7817 (.A1(W28957), .A2(W15298), .ZN(W36417));
  NOR2X1 G7818 (.A1(W5885), .A2(W21455), .ZN(O5233));
  NOR2X1 G7819 (.A1(W7151), .A2(W13915), .ZN(W14399));
  NOR2X1 G7820 (.A1(W35664), .A2(W15406), .ZN(O8384));
  NOR2X1 G7821 (.A1(W18075), .A2(W892), .ZN(O8385));
  NOR2X1 G7822 (.A1(W3861), .A2(I210), .ZN(W15241));
  NOR2X1 G7823 (.A1(W18744), .A2(W11337), .ZN(W30210));
  NOR2X1 G7824 (.A1(W14280), .A2(I409), .ZN(O8389));
  NOR2X1 G7825 (.A1(W3045), .A2(W25573), .ZN(O8390));
  NOR2X1 G7826 (.A1(W15784), .A2(W24821), .ZN(W36428));
  NOR2X1 G7827 (.A1(W1707), .A2(W3267), .ZN(O8391));
  NOR2X1 G7828 (.A1(W403), .A2(W5842), .ZN(W20583));
  NOR2X1 G7829 (.A1(W24187), .A2(W16108), .ZN(O5231));
  NOR2X1 G7830 (.A1(W3153), .A2(W12945), .ZN(O5501));
  NOR2X1 G7831 (.A1(I1590), .A2(W9406), .ZN(W16078));
  NOR2X1 G7832 (.A1(W11575), .A2(W5093), .ZN(O1117));
  NOR2X1 G7833 (.A1(W15641), .A2(W5120), .ZN(W16076));
  NOR2X1 G7834 (.A1(W15591), .A2(W15288), .ZN(W16075));
  NOR2X1 G7835 (.A1(W9863), .A2(W8978), .ZN(O5502));
  NOR2X1 G7836 (.A1(W16452), .A2(W9366), .ZN(O7425));
  NOR2X1 G7837 (.A1(W15183), .A2(W6726), .ZN(O7427));
  NOR2X1 G7838 (.A1(W12640), .A2(W12030), .ZN(O7428));
  NOR2X1 G7839 (.A1(W2550), .A2(W2887), .ZN(W16079));
  NOR2X1 G7840 (.A1(W25972), .A2(W27217), .ZN(O7431));
  NOR2X1 G7841 (.A1(W34363), .A2(W16424), .ZN(W34757));
  NOR2X1 G7842 (.A1(W12598), .A2(W783), .ZN(W16067));
  NOR2X1 G7843 (.A1(W10829), .A2(W5182), .ZN(W16066));
  NOR2X1 G7844 (.A1(W29362), .A2(W11137), .ZN(W34761));
  NOR2X1 G7845 (.A1(W15696), .A2(W24539), .ZN(W34762));
  NOR2X1 G7846 (.A1(W16128), .A2(W24104), .ZN(O7436));
  NOR2X1 G7847 (.A1(W12005), .A2(W6040), .ZN(W16059));
  NOR2X1 G7848 (.A1(W4787), .A2(W9253), .ZN(W16089));
  NOR2X1 G7849 (.A1(I258), .A2(W14300), .ZN(O7410));
  NOR2X1 G7850 (.A1(W12362), .A2(W4879), .ZN(W16096));
  NOR2X1 G7851 (.A1(W13753), .A2(W26924), .ZN(O7411));
  NOR2X1 G7852 (.A1(W21682), .A2(W28339), .ZN(W34726));
  NOR2X1 G7853 (.A1(W2932), .A2(W1724), .ZN(O7413));
  NOR2X1 G7854 (.A1(W32442), .A2(W6061), .ZN(W34729));
  NOR2X1 G7855 (.A1(W19849), .A2(W8185), .ZN(O7414));
  NOR2X1 G7856 (.A1(W29995), .A2(W22452), .ZN(O7415));
  NOR2X1 G7857 (.A1(W10988), .A2(W13742), .ZN(W34764));
  NOR2X1 G7858 (.A1(W5389), .A2(W428), .ZN(W16088));
  NOR2X1 G7859 (.A1(W720), .A2(I1094), .ZN(W16086));
  NOR2X1 G7860 (.A1(W31949), .A2(W29290), .ZN(O7417));
  NOR2X1 G7861 (.A1(W15373), .A2(W4745), .ZN(W30814));
  NOR2X1 G7862 (.A1(W2853), .A2(W3397), .ZN(W16083));
  NOR2X1 G7863 (.A1(W6668), .A2(W30801), .ZN(O7419));
  NOR2X1 G7864 (.A1(W15819), .A2(I566), .ZN(O7422));
  NOR2X1 G7865 (.A1(W5843), .A2(W9321), .ZN(O1108));
  NOR2X1 G7866 (.A1(W7286), .A2(W13356), .ZN(W30790));
  NOR2X1 G7867 (.A1(W3341), .A2(W9306), .ZN(W20021));
  NOR2X1 G7868 (.A1(W5642), .A2(W7839), .ZN(O1111));
  NOR2X1 G7869 (.A1(W3147), .A2(W13011), .ZN(W16032));
  NOR2X1 G7870 (.A1(W7196), .A2(W11860), .ZN(W20024));
  NOR2X1 G7871 (.A1(W24735), .A2(W25956), .ZN(O7453));
  NOR2X1 G7872 (.A1(W9213), .A2(W15382), .ZN(W16028));
  NOR2X1 G7873 (.A1(I1936), .A2(W4066), .ZN(W16027));
  NOR2X1 G7874 (.A1(W9376), .A2(W13013), .ZN(W34786));
  NOR2X1 G7875 (.A1(W966), .A2(W4786), .ZN(O1107));
  NOR2X1 G7876 (.A1(W1179), .A2(W11255), .ZN(O1106));
  NOR2X1 G7877 (.A1(I1836), .A2(W10934), .ZN(W16021));
  NOR2X1 G7878 (.A1(W14837), .A2(W5603), .ZN(O1105));
  NOR2X1 G7879 (.A1(I1846), .A2(W7631), .ZN(W16019));
  NOR2X1 G7880 (.A1(W11259), .A2(W13028), .ZN(O7456));
  NOR2X1 G7881 (.A1(W328), .A2(W12094), .ZN(W16017));
  NOR2X1 G7882 (.A1(W12911), .A2(W3719), .ZN(O5489));
  NOR2X1 G7883 (.A1(W7018), .A2(W28198), .ZN(O5493));
  NOR2X1 G7884 (.A1(W15108), .A2(W7263), .ZN(W16056));
  NOR2X1 G7885 (.A1(W5180), .A2(W2162), .ZN(W16055));
  NOR2X1 G7886 (.A1(W29059), .A2(W18601), .ZN(O7437));
  NOR2X1 G7887 (.A1(W10396), .A2(I1065), .ZN(W16052));
  NOR2X1 G7888 (.A1(W13782), .A2(W21989), .ZN(W34770));
  NOR2X1 G7889 (.A1(W4898), .A2(W1141), .ZN(O1114));
  NOR2X1 G7890 (.A1(W7399), .A2(W12587), .ZN(O5494));
  NOR2X1 G7891 (.A1(W29047), .A2(W23399), .ZN(O7439));
  NOR2X1 G7892 (.A1(W15040), .A2(W15638), .ZN(W16098));
  NOR2X1 G7893 (.A1(W1677), .A2(W3316), .ZN(O7443));
  NOR2X1 G7894 (.A1(W6565), .A2(W7130), .ZN(W16045));
  NOR2X1 G7895 (.A1(W11941), .A2(W17568), .ZN(W30794));
  NOR2X1 G7896 (.A1(W12729), .A2(W11383), .ZN(W16043));
  NOR2X1 G7897 (.A1(W21464), .A2(W18106), .ZN(W34779));
  NOR2X1 G7898 (.A1(W1843), .A2(W27709), .ZN(W34782));
  NOR2X1 G7899 (.A1(W2005), .A2(W9763), .ZN(W16038));
  NOR2X1 G7900 (.A1(W10901), .A2(W12084), .ZN(W16146));
  NOR2X1 G7901 (.A1(W4765), .A2(W6167), .ZN(W16157));
  NOR2X1 G7902 (.A1(W8023), .A2(W816), .ZN(W16155));
  NOR2X1 G7903 (.A1(W11947), .A2(I1110), .ZN(W16153));
  NOR2X1 G7904 (.A1(W4723), .A2(W11727), .ZN(W16152));
  NOR2X1 G7905 (.A1(W14751), .A2(W1655), .ZN(O7383));
  NOR2X1 G7906 (.A1(W26958), .A2(W22582), .ZN(O7384));
  NOR2X1 G7907 (.A1(W10014), .A2(W10442), .ZN(O7386));
  NOR2X1 G7908 (.A1(W15489), .A2(I1783), .ZN(W19991));
  NOR2X1 G7909 (.A1(W4352), .A2(W3270), .ZN(W16158));
  NOR2X1 G7910 (.A1(I1482), .A2(W2408), .ZN(O1131));
  NOR2X1 G7911 (.A1(W3950), .A2(W6795), .ZN(O5509));
  NOR2X1 G7912 (.A1(W30380), .A2(W5692), .ZN(W30825));
  NOR2X1 G7913 (.A1(W4603), .A2(W25558), .ZN(W34676));
  NOR2X1 G7914 (.A1(W15722), .A2(W17849), .ZN(W19994));
  NOR2X1 G7915 (.A1(W831), .A2(W13754), .ZN(W16140));
  NOR2X1 G7916 (.A1(W17934), .A2(W24891), .ZN(W34678));
  NOR2X1 G7917 (.A1(W28280), .A2(W23953), .ZN(W34679));
  NOR2X1 G7918 (.A1(W2429), .A2(W8385), .ZN(W16167));
  NOR2X1 G7919 (.A1(W3916), .A2(W27765), .ZN(O7375));
  NOR2X1 G7920 (.A1(W17331), .A2(W10273), .ZN(O7376));
  NOR2X1 G7921 (.A1(W13264), .A2(W14911), .ZN(W16174));
  NOR2X1 G7922 (.A1(W9459), .A2(W1533), .ZN(W16173));
  NOR2X1 G7923 (.A1(W31535), .A2(W5805), .ZN(O7377));
  NOR2X1 G7924 (.A1(W8939), .A2(W6265), .ZN(W16170));
  NOR2X1 G7925 (.A1(W7100), .A2(W11823), .ZN(O1135));
  NOR2X1 G7926 (.A1(W966), .A2(W12179), .ZN(O1134));
  NOR2X1 G7927 (.A1(W1162), .A2(W7351), .ZN(W16137));
  NOR2X1 G7928 (.A1(W5639), .A2(W11977), .ZN(W16166));
  NOR2X1 G7929 (.A1(W10099), .A2(W2819), .ZN(W16164));
  NOR2X1 G7930 (.A1(W5263), .A2(W10390), .ZN(O1133));
  NOR2X1 G7931 (.A1(W13533), .A2(W14835), .ZN(W16162));
  NOR2X1 G7932 (.A1(W8571), .A2(W10256), .ZN(W16161));
  NOR2X1 G7933 (.A1(W13357), .A2(W26586), .ZN(W34662));
  NOR2X1 G7934 (.A1(W2646), .A2(W11486), .ZN(W16159));
  NOR2X1 G7935 (.A1(W10662), .A2(W18376), .ZN(O7406));
  NOR2X1 G7936 (.A1(W14927), .A2(W5562), .ZN(O1124));
  NOR2X1 G7937 (.A1(W5397), .A2(W7921), .ZN(W16116));
  NOR2X1 G7938 (.A1(W8127), .A2(W6817), .ZN(O7401));
  NOR2X1 G7939 (.A1(W8333), .A2(W4219), .ZN(W20001));
  NOR2X1 G7940 (.A1(W12066), .A2(W7858), .ZN(O1123));
  NOR2X1 G7941 (.A1(W12653), .A2(W6981), .ZN(O1122));
  NOR2X1 G7942 (.A1(W854), .A2(I526), .ZN(W16111));
  NOR2X1 G7943 (.A1(W13279), .A2(W22297), .ZN(W34707));
  NOR2X1 G7944 (.A1(W6420), .A2(W12510), .ZN(W16119));
  NOR2X1 G7945 (.A1(W28889), .A2(W25516), .ZN(W34713));
  NOR2X1 G7946 (.A1(W15326), .A2(W2961), .ZN(W16106));
  NOR2X1 G7947 (.A1(W7490), .A2(W6503), .ZN(W34714));
  NOR2X1 G7948 (.A1(W1511), .A2(W14603), .ZN(W16104));
  NOR2X1 G7949 (.A1(W13571), .A2(W29334), .ZN(W30817));
  NOR2X1 G7950 (.A1(W9930), .A2(W15690), .ZN(W16102));
  NOR2X1 G7951 (.A1(W25358), .A2(W21637), .ZN(W34717));
  NOR2X1 G7952 (.A1(W13191), .A2(W13667), .ZN(W16099));
  NOR2X1 G7953 (.A1(W13365), .A2(W30606), .ZN(W30824));
  NOR2X1 G7954 (.A1(W8065), .A2(W8932), .ZN(W16136));
  NOR2X1 G7955 (.A1(W3226), .A2(W24828), .ZN(O7392));
  NOR2X1 G7956 (.A1(W26644), .A2(W6570), .ZN(W34683));
  NOR2X1 G7957 (.A1(W11975), .A2(W23932), .ZN(W34684));
  NOR2X1 G7958 (.A1(W31632), .A2(W34337), .ZN(W34687));
  NOR2X1 G7959 (.A1(W985), .A2(W4119), .ZN(W19995));
  NOR2X1 G7960 (.A1(W15330), .A2(W6403), .ZN(O1127));
  NOR2X1 G7961 (.A1(W9279), .A2(W8564), .ZN(O7394));
  NOR2X1 G7962 (.A1(W12356), .A2(W3447), .ZN(O5488));
  NOR2X1 G7963 (.A1(W17571), .A2(W4065), .ZN(W34693));
  NOR2X1 G7964 (.A1(W12867), .A2(W8250), .ZN(O1126));
  NOR2X1 G7965 (.A1(I592), .A2(W13543), .ZN(W16124));
  NOR2X1 G7966 (.A1(W10165), .A2(W17716), .ZN(W19998));
  NOR2X1 G7967 (.A1(W30960), .A2(W28361), .ZN(O7398));
  NOR2X1 G7968 (.A1(W18718), .A2(I1206), .ZN(W19999));
  NOR2X1 G7969 (.A1(W10769), .A2(I480), .ZN(O7400));
  NOR2X1 G7970 (.A1(W8961), .A2(W8572), .ZN(O5475));
  NOR2X1 G7971 (.A1(W9183), .A2(W26109), .ZN(W34916));
  NOR2X1 G7972 (.A1(W19556), .A2(I1367), .ZN(W34917));
  NOR2X1 G7973 (.A1(W7285), .A2(I1390), .ZN(W15916));
  NOR2X1 G7974 (.A1(W5774), .A2(W32809), .ZN(O7513));
  NOR2X1 G7975 (.A1(W12241), .A2(W426), .ZN(W15914));
  NOR2X1 G7976 (.A1(W34003), .A2(W23634), .ZN(O7514));
  NOR2X1 G7977 (.A1(W7190), .A2(W20924), .ZN(O7515));
  NOR2X1 G7978 (.A1(W20791), .A2(W25179), .ZN(O5476));
  NOR2X1 G7979 (.A1(W5243), .A2(W4242), .ZN(W15919));
  NOR2X1 G7980 (.A1(I462), .A2(W3894), .ZN(O1089));
  NOR2X1 G7981 (.A1(W18071), .A2(W6339), .ZN(O7519));
  NOR2X1 G7982 (.A1(W10464), .A2(W18706), .ZN(W20060));
  NOR2X1 G7983 (.A1(W1138), .A2(W4387), .ZN(O1919));
  NOR2X1 G7984 (.A1(W11737), .A2(W11117), .ZN(O7524));
  NOR2X1 G7985 (.A1(W7157), .A2(W12826), .ZN(W15903));
  NOR2X1 G7986 (.A1(W14331), .A2(W6244), .ZN(W30747));
  NOR2X1 G7987 (.A1(W17848), .A2(W4734), .ZN(W20064));
  NOR2X1 G7988 (.A1(W5812), .A2(W13994), .ZN(W20055));
  NOR2X1 G7989 (.A1(W12320), .A2(W7052), .ZN(W15936));
  NOR2X1 G7990 (.A1(W12620), .A2(W21489), .ZN(O7501));
  NOR2X1 G7991 (.A1(W12151), .A2(I1477), .ZN(W15934));
  NOR2X1 G7992 (.A1(W9113), .A2(W18005), .ZN(W34899));
  NOR2X1 G7993 (.A1(W12275), .A2(W11290), .ZN(W15932));
  NOR2X1 G7994 (.A1(W14548), .A2(W8166), .ZN(O5479));
  NOR2X1 G7995 (.A1(W15320), .A2(W15599), .ZN(O7505));
  NOR2X1 G7996 (.A1(W21811), .A2(W3944), .ZN(W30755));
  NOR2X1 G7997 (.A1(W5074), .A2(W2281), .ZN(W15900));
  NOR2X1 G7998 (.A1(W3314), .A2(W13887), .ZN(W15927));
  NOR2X1 G7999 (.A1(W10788), .A2(W1854), .ZN(W34909));
  NOR2X1 G8000 (.A1(W11429), .A2(W21448), .ZN(W34912));
  NOR2X1 G8001 (.A1(I853), .A2(W14055), .ZN(O1094));
  NOR2X1 G8002 (.A1(I436), .A2(W13344), .ZN(W15923));
  NOR2X1 G8003 (.A1(I117), .A2(I509), .ZN(O1093));
  NOR2X1 G8004 (.A1(W6889), .A2(W11893), .ZN(W20057));
  NOR2X1 G8005 (.A1(W13436), .A2(W2874), .ZN(W15868));
  NOR2X1 G8006 (.A1(W20258), .A2(W21341), .ZN(O7533));
  NOR2X1 G8007 (.A1(W17991), .A2(W11898), .ZN(W20073));
  NOR2X1 G8008 (.A1(W6910), .A2(I1026), .ZN(W15875));
  NOR2X1 G8009 (.A1(W12384), .A2(W3627), .ZN(O1082));
  NOR2X1 G8010 (.A1(W1203), .A2(W2638), .ZN(W20075));
  NOR2X1 G8011 (.A1(I1069), .A2(W10958), .ZN(W15872));
  NOR2X1 G8012 (.A1(W3125), .A2(W9182), .ZN(W20077));
  NOR2X1 G8013 (.A1(I1134), .A2(W17782), .ZN(W34958));
  NOR2X1 G8014 (.A1(W32967), .A2(W23421), .ZN(W34949));
  NOR2X1 G8015 (.A1(W33144), .A2(W1205), .ZN(W34960));
  NOR2X1 G8016 (.A1(W383), .A2(W9364), .ZN(W15866));
  NOR2X1 G8017 (.A1(W6983), .A2(W2581), .ZN(W15865));
  NOR2X1 G8018 (.A1(W3695), .A2(W17325), .ZN(O7537));
  NOR2X1 G8019 (.A1(W14759), .A2(W7196), .ZN(O5469));
  NOR2X1 G8020 (.A1(W13692), .A2(W435), .ZN(O1078));
  NOR2X1 G8021 (.A1(W33005), .A2(W2488), .ZN(O7540));
  NOR2X1 G8022 (.A1(W6356), .A2(W593), .ZN(W15858));
  NOR2X1 G8023 (.A1(W14622), .A2(W7307), .ZN(W15890));
  NOR2X1 G8024 (.A1(W18247), .A2(W28560), .ZN(W34936));
  NOR2X1 G8025 (.A1(W12554), .A2(W3348), .ZN(O5473));
  NOR2X1 G8026 (.A1(W10095), .A2(W7550), .ZN(O1087));
  NOR2X1 G8027 (.A1(W19771), .A2(W18650), .ZN(O7527));
  NOR2X1 G8028 (.A1(W1316), .A2(W6212), .ZN(W15895));
  NOR2X1 G8029 (.A1(W17422), .A2(W20598), .ZN(O5472));
  NOR2X1 G8030 (.A1(W16923), .A2(W28553), .ZN(O5471));
  NOR2X1 G8031 (.A1(W14598), .A2(W4957), .ZN(W15892));
  NOR2X1 G8032 (.A1(W8521), .A2(W21942), .ZN(W34895));
  NOR2X1 G8033 (.A1(W18535), .A2(W3757), .ZN(O7530));
  NOR2X1 G8034 (.A1(W31735), .A2(W33435), .ZN(W34944));
  NOR2X1 G8035 (.A1(W3215), .A2(W11425), .ZN(W15887));
  NOR2X1 G8036 (.A1(W1956), .A2(W13168), .ZN(W15885));
  NOR2X1 G8037 (.A1(W1012), .A2(I1074), .ZN(W15884));
  NOR2X1 G8038 (.A1(W9353), .A2(W3455), .ZN(O1084));
  NOR2X1 G8039 (.A1(W14787), .A2(W16376), .ZN(W20070));
  NOR2X1 G8040 (.A1(W23589), .A2(W9436), .ZN(W34837));
  NOR2X1 G8041 (.A1(W20214), .A2(W15177), .ZN(W30779));
  NOR2X1 G8042 (.A1(W12496), .A2(W4154), .ZN(O1911));
  NOR2X1 G8043 (.A1(I849), .A2(W24482), .ZN(O7470));
  NOR2X1 G8044 (.A1(W5025), .A2(W12217), .ZN(W15993));
  NOR2X1 G8045 (.A1(W4847), .A2(W8253), .ZN(W15992));
  NOR2X1 G8046 (.A1(W11639), .A2(W113), .ZN(O7471));
  NOR2X1 G8047 (.A1(W1915), .A2(W4598), .ZN(W34833));
  NOR2X1 G8048 (.A1(W21152), .A2(W22984), .ZN(W30775));
  NOR2X1 G8049 (.A1(W22949), .A2(W23451), .ZN(O7467));
  NOR2X1 G8050 (.A1(W29635), .A2(W12926), .ZN(W34838));
  NOR2X1 G8051 (.A1(W8007), .A2(W4781), .ZN(O1099));
  NOR2X1 G8052 (.A1(I1226), .A2(W31300), .ZN(O7475));
  NOR2X1 G8053 (.A1(W18039), .A2(W6869), .ZN(W34843));
  NOR2X1 G8054 (.A1(W17734), .A2(W18307), .ZN(W20038));
  NOR2X1 G8055 (.A1(W32779), .A2(W10822), .ZN(O7476));
  NOR2X1 G8056 (.A1(W4413), .A2(I297), .ZN(O7477));
  NOR2X1 G8057 (.A1(W8127), .A2(I625), .ZN(W15977));
  NOR2X1 G8058 (.A1(W34447), .A2(W31480), .ZN(O7461));
  NOR2X1 G8059 (.A1(W1662), .A2(W541), .ZN(W34809));
  NOR2X1 G8060 (.A1(W5496), .A2(I779), .ZN(W16013));
  NOR2X1 G8061 (.A1(W14786), .A2(W9974), .ZN(W16012));
  NOR2X1 G8062 (.A1(W22801), .A2(W27239), .ZN(W30782));
  NOR2X1 G8063 (.A1(W16164), .A2(W9715), .ZN(W34811));
  NOR2X1 G8064 (.A1(W29666), .A2(W18203), .ZN(W34812));
  NOR2X1 G8065 (.A1(W15932), .A2(W11717), .ZN(W16008));
  NOR2X1 G8066 (.A1(I124), .A2(W13295), .ZN(O7460));
  NOR2X1 G8067 (.A1(W5210), .A2(W19644), .ZN(O5483));
  NOR2X1 G8068 (.A1(W8456), .A2(W4578), .ZN(W16004));
  NOR2X1 G8069 (.A1(W24644), .A2(W15220), .ZN(O7463));
  NOR2X1 G8070 (.A1(W11058), .A2(W5473), .ZN(W16002));
  NOR2X1 G8071 (.A1(W9851), .A2(W19223), .ZN(W20031));
  NOR2X1 G8072 (.A1(W25327), .A2(W24808), .ZN(W30780));
  NOR2X1 G8073 (.A1(W9600), .A2(W655), .ZN(W15999));
  NOR2X1 G8074 (.A1(W22845), .A2(W7911), .ZN(O7466));
  NOR2X1 G8075 (.A1(W13835), .A2(W1950), .ZN(O7495));
  NOR2X1 G8076 (.A1(W28586), .A2(W5096), .ZN(W30766));
  NOR2X1 G8077 (.A1(W30183), .A2(I858), .ZN(W34874));
  NOR2X1 G8078 (.A1(W20320), .A2(W31617), .ZN(W34875));
  NOR2X1 G8079 (.A1(W8852), .A2(W8865), .ZN(W15954));
  NOR2X1 G8080 (.A1(W23876), .A2(W31586), .ZN(W34876));
  NOR2X1 G8081 (.A1(W18127), .A2(W31246), .ZN(O7492));
  NOR2X1 G8082 (.A1(W10695), .A2(W1927), .ZN(O1095));
  NOR2X1 G8083 (.A1(W19980), .A2(W17589), .ZN(O7494));
  NOR2X1 G8084 (.A1(W29534), .A2(W8756), .ZN(W30767));
  NOR2X1 G8085 (.A1(W18898), .A2(W5559), .ZN(O1916));
  NOR2X1 G8086 (.A1(W13017), .A2(W21433), .ZN(W34887));
  NOR2X1 G8087 (.A1(W25688), .A2(W32756), .ZN(O7497));
  NOR2X1 G8088 (.A1(W3906), .A2(W6232), .ZN(W15943));
  NOR2X1 G8089 (.A1(W10827), .A2(W18209), .ZN(W20051));
  NOR2X1 G8090 (.A1(W23739), .A2(W12798), .ZN(W30760));
  NOR2X1 G8091 (.A1(W3760), .A2(W3883), .ZN(O7499));
  NOR2X1 G8092 (.A1(W13775), .A2(W9579), .ZN(W15938));
  NOR2X1 G8093 (.A1(W5942), .A2(W6627), .ZN(W15967));
  NOR2X1 G8094 (.A1(W25618), .A2(W31559), .ZN(O7480));
  NOR2X1 G8095 (.A1(W164), .A2(W2366), .ZN(W15974));
  NOR2X1 G8096 (.A1(W24699), .A2(W32910), .ZN(W34852));
  NOR2X1 G8097 (.A1(W15156), .A2(W1684), .ZN(O7482));
  NOR2X1 G8098 (.A1(W3740), .A2(W13503), .ZN(O7483));
  NOR2X1 G8099 (.A1(W11675), .A2(W2264), .ZN(W15970));
  NOR2X1 G8100 (.A1(W24154), .A2(W20960), .ZN(W30770));
  NOR2X1 G8101 (.A1(W28142), .A2(W22101), .ZN(W34857));
  NOR2X1 G8102 (.A1(W16152), .A2(I1880), .ZN(O1137));
  NOR2X1 G8103 (.A1(W10230), .A2(I1480), .ZN(W15966));
  NOR2X1 G8104 (.A1(W9574), .A2(W8049), .ZN(W34859));
  NOR2X1 G8105 (.A1(W12861), .A2(W13779), .ZN(W20043));
  NOR2X1 G8106 (.A1(W19932), .A2(W21471), .ZN(W34863));
  NOR2X1 G8107 (.A1(W7478), .A2(W1779), .ZN(W15961));
  NOR2X1 G8108 (.A1(W6287), .A2(W2327), .ZN(W30768));
  NOR2X1 G8109 (.A1(W18231), .A2(W32599), .ZN(W34867));
  NOR2X1 G8110 (.A1(W2639), .A2(W10565), .ZN(W16380));
  NOR2X1 G8111 (.A1(W13626), .A2(W712), .ZN(W16390));
  NOR2X1 G8112 (.A1(W18614), .A2(W4128), .ZN(O5551));
  NOR2X1 G8113 (.A1(W4760), .A2(I467), .ZN(W16388));
  NOR2X1 G8114 (.A1(W7716), .A2(W1532), .ZN(W16385));
  NOR2X1 G8115 (.A1(W4090), .A2(W3953), .ZN(O1171));
  NOR2X1 G8116 (.A1(W6270), .A2(W7114), .ZN(W16383));
  NOR2X1 G8117 (.A1(W6844), .A2(W9831), .ZN(W19917));
  NOR2X1 G8118 (.A1(W9896), .A2(W4448), .ZN(W19918));
  NOR2X1 G8119 (.A1(W8881), .A2(W4565), .ZN(O7273));
  NOR2X1 G8120 (.A1(W9232), .A2(W20534), .ZN(O7281));
  NOR2X1 G8121 (.A1(W11323), .A2(W28682), .ZN(O5545));
  NOR2X1 G8122 (.A1(I362), .A2(W4424), .ZN(O1884));
  NOR2X1 G8123 (.A1(W12509), .A2(W10811), .ZN(W16375));
  NOR2X1 G8124 (.A1(W27068), .A2(W2019), .ZN(W30899));
  NOR2X1 G8125 (.A1(W31005), .A2(W31178), .ZN(O7284));
  NOR2X1 G8126 (.A1(W22878), .A2(W7773), .ZN(W34487));
  NOR2X1 G8127 (.A1(I555), .A2(W5243), .ZN(W16370));
  NOR2X1 G8128 (.A1(W24397), .A2(W34361), .ZN(W34459));
  NOR2X1 G8129 (.A1(W9), .A2(W11599), .ZN(W16410));
  NOR2X1 G8130 (.A1(W1098), .A2(W25956), .ZN(O7265));
  NOR2X1 G8131 (.A1(W8583), .A2(W14931), .ZN(W16408));
  NOR2X1 G8132 (.A1(W3977), .A2(W12537), .ZN(O5553));
  NOR2X1 G8133 (.A1(W13881), .A2(W289), .ZN(W16405));
  NOR2X1 G8134 (.A1(W11439), .A2(W10087), .ZN(O1173));
  NOR2X1 G8135 (.A1(W11695), .A2(W2993), .ZN(W16403));
  NOR2X1 G8136 (.A1(W25682), .A2(W6469), .ZN(W34458));
  NOR2X1 G8137 (.A1(W28500), .A2(W20399), .ZN(W34488));
  NOR2X1 G8138 (.A1(W4473), .A2(W5095), .ZN(W16399));
  NOR2X1 G8139 (.A1(W33292), .A2(W5864), .ZN(W34461));
  NOR2X1 G8140 (.A1(W21476), .A2(I719), .ZN(O7269));
  NOR2X1 G8141 (.A1(W4765), .A2(W9251), .ZN(O7271));
  NOR2X1 G8142 (.A1(W2163), .A2(W1926), .ZN(W16394));
  NOR2X1 G8143 (.A1(W4898), .A2(W20638), .ZN(W30916));
  NOR2X1 G8144 (.A1(W10564), .A2(W3059), .ZN(W19913));
  NOR2X1 G8145 (.A1(W2332), .A2(W10826), .ZN(W16342));
  NOR2X1 G8146 (.A1(W2856), .A2(I787), .ZN(W16351));
  NOR2X1 G8147 (.A1(W9402), .A2(W14288), .ZN(O1886));
  NOR2X1 G8148 (.A1(W10487), .A2(W34220), .ZN(O7296));
  NOR2X1 G8149 (.A1(W10894), .A2(W11342), .ZN(W34506));
  NOR2X1 G8150 (.A1(W12853), .A2(W9500), .ZN(W16347));
  NOR2X1 G8151 (.A1(W14378), .A2(W4792), .ZN(W16346));
  NOR2X1 G8152 (.A1(W20313), .A2(W31618), .ZN(W34507));
  NOR2X1 G8153 (.A1(W13407), .A2(I124), .ZN(W16344));
  NOR2X1 G8154 (.A1(W7031), .A2(W2478), .ZN(W16352));
  NOR2X1 G8155 (.A1(W3945), .A2(W11415), .ZN(W16341));
  NOR2X1 G8156 (.A1(W20468), .A2(W24400), .ZN(W34511));
  NOR2X1 G8157 (.A1(W4333), .A2(W30683), .ZN(O7301));
  NOR2X1 G8158 (.A1(I348), .A2(W246), .ZN(W19931));
  NOR2X1 G8159 (.A1(W13693), .A2(W6931), .ZN(W16337));
  NOR2X1 G8160 (.A1(I1975), .A2(W6774), .ZN(W19932));
  NOR2X1 G8161 (.A1(W2343), .A2(W8003), .ZN(W16335));
  NOR2X1 G8162 (.A1(W17357), .A2(I1542), .ZN(O1887));
  NOR2X1 G8163 (.A1(I866), .A2(W24560), .ZN(O7289));
  NOR2X1 G8164 (.A1(W4680), .A2(W13074), .ZN(O1169));
  NOR2X1 G8165 (.A1(W8250), .A2(W6200), .ZN(W16367));
  NOR2X1 G8166 (.A1(I1058), .A2(W15781), .ZN(W16366));
  NOR2X1 G8167 (.A1(W315), .A2(W17072), .ZN(W19924));
  NOR2X1 G8168 (.A1(W5325), .A2(W2828), .ZN(W16364));
  NOR2X1 G8169 (.A1(W28377), .A2(W15162), .ZN(O5541));
  NOR2X1 G8170 (.A1(W18163), .A2(W17272), .ZN(W19926));
  NOR2X1 G8171 (.A1(W23425), .A2(W12987), .ZN(W30895));
  NOR2X1 G8172 (.A1(W9192), .A2(I1128), .ZN(W16411));
  NOR2X1 G8173 (.A1(W8474), .A2(W8451), .ZN(W19928));
  NOR2X1 G8174 (.A1(W9705), .A2(W23529), .ZN(O7291));
  NOR2X1 G8175 (.A1(W15302), .A2(W8175), .ZN(W16357));
  NOR2X1 G8176 (.A1(W14556), .A2(W2340), .ZN(O1164));
  NOR2X1 G8177 (.A1(W31054), .A2(W29173), .ZN(O7292));
  NOR2X1 G8178 (.A1(W2002), .A2(W5830), .ZN(W16354));
  NOR2X1 G8179 (.A1(W31652), .A2(W6513), .ZN(O7293));
  NOR2X1 G8180 (.A1(W2685), .A2(W4700), .ZN(W16464));
  NOR2X1 G8181 (.A1(I1909), .A2(W4882), .ZN(W16474));
  NOR2X1 G8182 (.A1(W3986), .A2(W16019), .ZN(W34402));
  NOR2X1 G8183 (.A1(W11960), .A2(W6572), .ZN(W16472));
  NOR2X1 G8184 (.A1(W3858), .A2(W19708), .ZN(W19887));
  NOR2X1 G8185 (.A1(W10773), .A2(W19577), .ZN(O7236));
  NOR2X1 G8186 (.A1(W31088), .A2(W33369), .ZN(O7238));
  NOR2X1 G8187 (.A1(W7054), .A2(W9815), .ZN(W16466));
  NOR2X1 G8188 (.A1(W5812), .A2(W16103), .ZN(W16465));
  NOR2X1 G8189 (.A1(W2286), .A2(W1136), .ZN(W16475));
  NOR2X1 G8190 (.A1(W15105), .A2(W18306), .ZN(O5563));
  NOR2X1 G8191 (.A1(W18936), .A2(W11476), .ZN(O7239));
  NOR2X1 G8192 (.A1(W6136), .A2(W14833), .ZN(W16460));
  NOR2X1 G8193 (.A1(W12692), .A2(W14280), .ZN(W19893));
  NOR2X1 G8194 (.A1(W13965), .A2(W4582), .ZN(W16457));
  NOR2X1 G8195 (.A1(W581), .A2(W1617), .ZN(W16456));
  NOR2X1 G8196 (.A1(W8121), .A2(W14897), .ZN(W16455));
  NOR2X1 G8197 (.A1(W15313), .A2(W4446), .ZN(W30937));
  NOR2X1 G8198 (.A1(W17332), .A2(W15203), .ZN(W30945));
  NOR2X1 G8199 (.A1(W421), .A2(W29503), .ZN(W34388));
  NOR2X1 G8200 (.A1(W12542), .A2(W30330), .ZN(O7225));
  NOR2X1 G8201 (.A1(W16276), .A2(W6233), .ZN(W16491));
  NOR2X1 G8202 (.A1(I1911), .A2(W27312), .ZN(O7226));
  NOR2X1 G8203 (.A1(W6316), .A2(W19857), .ZN(O5566));
  NOR2X1 G8204 (.A1(W5354), .A2(W3469), .ZN(W16487));
  NOR2X1 G8205 (.A1(W14952), .A2(W33764), .ZN(O7228));
  NOR2X1 G8206 (.A1(W23853), .A2(W16188), .ZN(W30946));
  NOR2X1 G8207 (.A1(W10065), .A2(I20), .ZN(O5560));
  NOR2X1 G8208 (.A1(I356), .A2(W4353), .ZN(W16483));
  NOR2X1 G8209 (.A1(W4643), .A2(W10827), .ZN(W16482));
  NOR2X1 G8210 (.A1(W27323), .A2(W3255), .ZN(O7231));
  NOR2X1 G8211 (.A1(W18473), .A2(W22843), .ZN(O7232));
  NOR2X1 G8212 (.A1(W4830), .A2(W19590), .ZN(W19884));
  NOR2X1 G8213 (.A1(W14733), .A2(I296), .ZN(W19886));
  NOR2X1 G8214 (.A1(W14111), .A2(I1770), .ZN(O1182));
  NOR2X1 G8215 (.A1(W23432), .A2(W26944), .ZN(W34443));
  NOR2X1 G8216 (.A1(W12984), .A2(W11960), .ZN(W30930));
  NOR2X1 G8217 (.A1(W4754), .A2(W9878), .ZN(O1880));
  NOR2X1 G8218 (.A1(W27391), .A2(W21675), .ZN(O7256));
  NOR2X1 G8219 (.A1(W4989), .A2(W14414), .ZN(W19901));
  NOR2X1 G8220 (.A1(W20258), .A2(W27059), .ZN(W34439));
  NOR2X1 G8221 (.A1(W1878), .A2(W11915), .ZN(O1178));
  NOR2X1 G8222 (.A1(W88), .A2(W29332), .ZN(W34441));
  NOR2X1 G8223 (.A1(W4711), .A2(W11128), .ZN(W16424));
  NOR2X1 G8224 (.A1(I1592), .A2(W457), .ZN(W16434));
  NOR2X1 G8225 (.A1(W2674), .A2(W6575), .ZN(W16422));
  NOR2X1 G8226 (.A1(W6953), .A2(W10169), .ZN(W16420));
  NOR2X1 G8227 (.A1(W11114), .A2(W22802), .ZN(O7262));
  NOR2X1 G8228 (.A1(W26930), .A2(W7193), .ZN(W34448));
  NOR2X1 G8229 (.A1(W31678), .A2(W424), .ZN(W34449));
  NOR2X1 G8230 (.A1(W6154), .A2(W9476), .ZN(W16415));
  NOR2X1 G8231 (.A1(W10609), .A2(W13593), .ZN(W16413));
  NOR2X1 G8232 (.A1(W8042), .A2(W22835), .ZN(W30922));
  NOR2X1 G8233 (.A1(W12750), .A2(W15356), .ZN(O1879));
  NOR2X1 G8234 (.A1(W13122), .A2(W1330), .ZN(W16451));
  NOR2X1 G8235 (.A1(W15419), .A2(W1819), .ZN(W16450));
  NOR2X1 G8236 (.A1(W30554), .A2(W12371), .ZN(W34419));
  NOR2X1 G8237 (.A1(W3733), .A2(I1008), .ZN(O7246));
  NOR2X1 G8238 (.A1(W91), .A2(W652), .ZN(W16446));
  NOR2X1 G8239 (.A1(W14659), .A2(W7936), .ZN(O1180));
  NOR2X1 G8240 (.A1(W9674), .A2(W14514), .ZN(W16444));
  NOR2X1 G8241 (.A1(W16773), .A2(W884), .ZN(O7247));
  NOR2X1 G8242 (.A1(W155), .A2(W20435), .ZN(O7307));
  NOR2X1 G8243 (.A1(W10784), .A2(W5113), .ZN(W16441));
  NOR2X1 G8244 (.A1(W33896), .A2(W24995), .ZN(W34426));
  NOR2X1 G8245 (.A1(W8667), .A2(W9694), .ZN(O7252));
  NOR2X1 G8246 (.A1(W7963), .A2(W13932), .ZN(W16438));
  NOR2X1 G8247 (.A1(W9182), .A2(W3270), .ZN(W16437));
  NOR2X1 G8248 (.A1(W34232), .A2(W19594), .ZN(W34430));
  NOR2X1 G8249 (.A1(W10624), .A2(W714), .ZN(W16435));
  NOR2X1 G8250 (.A1(W13653), .A2(W17034), .ZN(O7354));
  NOR2X1 G8251 (.A1(W13175), .A2(W9708), .ZN(O1143));
  NOR2X1 G8252 (.A1(W8472), .A2(W22487), .ZN(O7348));
  NOR2X1 G8253 (.A1(W4976), .A2(I1731), .ZN(W16235));
  NOR2X1 G8254 (.A1(W29550), .A2(W32111), .ZN(O7350));
  NOR2X1 G8255 (.A1(W5988), .A2(W7195), .ZN(W16233));
  NOR2X1 G8256 (.A1(W32120), .A2(W29575), .ZN(O7351));
  NOR2X1 G8257 (.A1(W9252), .A2(W25005), .ZN(W34611));
  NOR2X1 G8258 (.A1(W5204), .A2(I624), .ZN(W19963));
  NOR2X1 G8259 (.A1(I1075), .A2(W6064), .ZN(W16238));
  NOR2X1 G8260 (.A1(W8076), .A2(W11701), .ZN(O7355));
  NOR2X1 G8261 (.A1(W7281), .A2(W18771), .ZN(W19965));
  NOR2X1 G8262 (.A1(W8519), .A2(W11658), .ZN(W16225));
  NOR2X1 G8263 (.A1(W5553), .A2(W3247), .ZN(O1142));
  NOR2X1 G8264 (.A1(W5302), .A2(W8025), .ZN(W16222));
  NOR2X1 G8265 (.A1(W25479), .A2(W6541), .ZN(W34620));
  NOR2X1 G8266 (.A1(W3006), .A2(W2048), .ZN(W16220));
  NOR2X1 G8267 (.A1(W11418), .A2(W9939), .ZN(O1141));
  NOR2X1 G8268 (.A1(W15551), .A2(W2808), .ZN(W34598));
  NOR2X1 G8269 (.A1(W7607), .A2(W30508), .ZN(W34591));
  NOR2X1 G8270 (.A1(W5448), .A2(W584), .ZN(W34592));
  NOR2X1 G8271 (.A1(W2645), .A2(W9991), .ZN(W16254));
  NOR2X1 G8272 (.A1(W15806), .A2(W14182), .ZN(W16252));
  NOR2X1 G8273 (.A1(I27), .A2(W6248), .ZN(O5525));
  NOR2X1 G8274 (.A1(I246), .A2(W10690), .ZN(W16249));
  NOR2X1 G8275 (.A1(W14192), .A2(W13558), .ZN(W16248));
  NOR2X1 G8276 (.A1(W18450), .A2(W15190), .ZN(O1898));
  NOR2X1 G8277 (.A1(W8067), .A2(W894), .ZN(W30856));
  NOR2X1 G8278 (.A1(W10046), .A2(W13524), .ZN(O1145));
  NOR2X1 G8279 (.A1(W27514), .A2(W8135), .ZN(W30860));
  NOR2X1 G8280 (.A1(W4570), .A2(W14864), .ZN(W16243));
  NOR2X1 G8281 (.A1(W12033), .A2(W6198), .ZN(W16242));
  NOR2X1 G8282 (.A1(W19303), .A2(W18388), .ZN(W34600));
  NOR2X1 G8283 (.A1(W10059), .A2(W8844), .ZN(W16240));
  NOR2X1 G8284 (.A1(W498), .A2(I1138), .ZN(W16239));
  NOR2X1 G8285 (.A1(W3004), .A2(W13419), .ZN(W16188));
  NOR2X1 G8286 (.A1(W3170), .A2(W8706), .ZN(W16199));
  NOR2X1 G8287 (.A1(W14482), .A2(W4950), .ZN(W16197));
  NOR2X1 G8288 (.A1(W6528), .A2(W5629), .ZN(W16195));
  NOR2X1 G8289 (.A1(W9116), .A2(W25595), .ZN(O7370));
  NOR2X1 G8290 (.A1(W9242), .A2(W19152), .ZN(W19979));
  NOR2X1 G8291 (.A1(W18340), .A2(W14869), .ZN(W19980));
  NOR2X1 G8292 (.A1(W10852), .A2(W2557), .ZN(W30843));
  NOR2X1 G8293 (.A1(I880), .A2(W7184), .ZN(W16189));
  NOR2X1 G8294 (.A1(W27850), .A2(W2429), .ZN(O7368));
  NOR2X1 G8295 (.A1(W1981), .A2(W14156), .ZN(W16187));
  NOR2X1 G8296 (.A1(W13065), .A2(W2329), .ZN(W34648));
  NOR2X1 G8297 (.A1(W12927), .A2(I1312), .ZN(W16185));
  NOR2X1 G8298 (.A1(W130), .A2(I76), .ZN(O5518));
  NOR2X1 G8299 (.A1(W11742), .A2(W4765), .ZN(O5515));
  NOR2X1 G8300 (.A1(I644), .A2(W4168), .ZN(W16182));
  NOR2X1 G8301 (.A1(W10086), .A2(W15822), .ZN(W16181));
  NOR2X1 G8302 (.A1(I562), .A2(W29283), .ZN(O7372));
  NOR2X1 G8303 (.A1(W10198), .A2(I1640), .ZN(W16209));
  NOR2X1 G8304 (.A1(I394), .A2(W5329), .ZN(W16217));
  NOR2X1 G8305 (.A1(W1065), .A2(W10640), .ZN(W30855));
  NOR2X1 G8306 (.A1(W383), .A2(W2048), .ZN(W34623));
  NOR2X1 G8307 (.A1(W13505), .A2(W12404), .ZN(W34624));
  NOR2X1 G8308 (.A1(W13253), .A2(W10775), .ZN(W19969));
  NOR2X1 G8309 (.A1(W21244), .A2(W10705), .ZN(W30854));
  NOR2X1 G8310 (.A1(W29185), .A2(W1327), .ZN(O7361));
  NOR2X1 G8311 (.A1(W3699), .A2(W9340), .ZN(W16210));
  NOR2X1 G8312 (.A1(W13327), .A2(W22809), .ZN(O5527));
  NOR2X1 G8313 (.A1(W25613), .A2(W5907), .ZN(W30852));
  NOR2X1 G8314 (.A1(W15225), .A2(W9548), .ZN(W16207));
  NOR2X1 G8315 (.A1(W6607), .A2(W10457), .ZN(W19972));
  NOR2X1 G8316 (.A1(W553), .A2(W16642), .ZN(O5523));
  NOR2X1 G8317 (.A1(W3661), .A2(W3216), .ZN(O1138));
  NOR2X1 G8318 (.A1(W13725), .A2(W2236), .ZN(W16203));
  NOR2X1 G8319 (.A1(W1533), .A2(W7655), .ZN(W19975));
  NOR2X1 G8320 (.A1(W1106), .A2(W809), .ZN(W30885));
  NOR2X1 G8321 (.A1(W2790), .A2(W16704), .ZN(W34537));
  NOR2X1 G8322 (.A1(I622), .A2(W5644), .ZN(W16314));
  NOR2X1 G8323 (.A1(W16602), .A2(W17536), .ZN(O1890));
  NOR2X1 G8324 (.A1(W5174), .A2(W3153), .ZN(W16312));
  NOR2X1 G8325 (.A1(W14771), .A2(W4985), .ZN(O7317));
  NOR2X1 G8326 (.A1(W3101), .A2(W10557), .ZN(W16310));
  NOR2X1 G8327 (.A1(W25406), .A2(W31796), .ZN(O7318));
  NOR2X1 G8328 (.A1(W10289), .A2(W14513), .ZN(W16308));
  NOR2X1 G8329 (.A1(W11178), .A2(W13967), .ZN(W16316));
  NOR2X1 G8330 (.A1(W11744), .A2(W32804), .ZN(O7319));
  NOR2X1 G8331 (.A1(W11121), .A2(W12902), .ZN(W16305));
  NOR2X1 G8332 (.A1(W10178), .A2(W14533), .ZN(W16304));
  NOR2X1 G8333 (.A1(W1439), .A2(W5168), .ZN(W16303));
  NOR2X1 G8334 (.A1(W8962), .A2(W9704), .ZN(W16302));
  NOR2X1 G8335 (.A1(W16225), .A2(W2830), .ZN(W16301));
  NOR2X1 G8336 (.A1(W33667), .A2(W20324), .ZN(O7320));
  NOR2X1 G8337 (.A1(W11747), .A2(W2843), .ZN(O1156));
  NOR2X1 G8338 (.A1(W16386), .A2(W1947), .ZN(W34531));
  NOR2X1 G8339 (.A1(W16990), .A2(W7845), .ZN(O7308));
  NOR2X1 G8340 (.A1(W2795), .A2(W21817), .ZN(O7309));
  NOR2X1 G8341 (.A1(W8426), .A2(W18716), .ZN(W30892));
  NOR2X1 G8342 (.A1(W11772), .A2(W9126), .ZN(W16329));
  NOR2X1 G8343 (.A1(W13492), .A2(W5239), .ZN(O1159));
  NOR2X1 G8344 (.A1(W5524), .A2(W20158), .ZN(O7310));
  NOR2X1 G8345 (.A1(W27650), .A2(W7017), .ZN(O5536));
  NOR2X1 G8346 (.A1(W11371), .A2(W30673), .ZN(W34530));
  NOR2X1 G8347 (.A1(W11020), .A2(W10165), .ZN(W16297));
  NOR2X1 G8348 (.A1(W18203), .A2(W11343), .ZN(O1888));
  NOR2X1 G8349 (.A1(W19310), .A2(W27324), .ZN(W34533));
  NOR2X1 G8350 (.A1(I1632), .A2(W1373), .ZN(O5535));
  NOR2X1 G8351 (.A1(W11068), .A2(W9126), .ZN(O1158));
  NOR2X1 G8352 (.A1(W22758), .A2(W1558), .ZN(O7313));
  NOR2X1 G8353 (.A1(W5834), .A2(W7838), .ZN(W16318));
  NOR2X1 G8354 (.A1(W24669), .A2(W12684), .ZN(W30886));
  NOR2X1 G8355 (.A1(W14568), .A2(W402), .ZN(W34580));
  NOR2X1 G8356 (.A1(W15433), .A2(W11996), .ZN(W34572));
  NOR2X1 G8357 (.A1(W10754), .A2(W11881), .ZN(W16272));
  NOR2X1 G8358 (.A1(W5449), .A2(W19601), .ZN(W34573));
  NOR2X1 G8359 (.A1(W8094), .A2(W23537), .ZN(W34574));
  NOR2X1 G8360 (.A1(W22846), .A2(W5957), .ZN(O7335));
  NOR2X1 G8361 (.A1(W25293), .A2(W13316), .ZN(O7336));
  NOR2X1 G8362 (.A1(W12175), .A2(W14869), .ZN(O1149));
  NOR2X1 G8363 (.A1(W2192), .A2(W5063), .ZN(O1894));
  NOR2X1 G8364 (.A1(W10055), .A2(W5469), .ZN(O1151));
  NOR2X1 G8365 (.A1(W6046), .A2(W11869), .ZN(W19953));
  NOR2X1 G8366 (.A1(W15545), .A2(I1317), .ZN(W30868));
  NOR2X1 G8367 (.A1(W6992), .A2(W9279), .ZN(W19955));
  NOR2X1 G8368 (.A1(W17855), .A2(W3665), .ZN(O7342));
  NOR2X1 G8369 (.A1(W18620), .A2(W11676), .ZN(W30867));
  NOR2X1 G8370 (.A1(W16071), .A2(W23183), .ZN(W34589));
  NOR2X1 G8371 (.A1(W10359), .A2(W14522), .ZN(W16258));
  NOR2X1 G8372 (.A1(W25346), .A2(W26034), .ZN(W34561));
  NOR2X1 G8373 (.A1(W24864), .A2(W6246), .ZN(W30883));
  NOR2X1 G8374 (.A1(W15908), .A2(W7232), .ZN(W16295));
  NOR2X1 G8375 (.A1(W31621), .A2(W25184), .ZN(W34552));
  NOR2X1 G8376 (.A1(W9275), .A2(W34482), .ZN(O7326));
  NOR2X1 G8377 (.A1(W5163), .A2(I1730), .ZN(O1892));
  NOR2X1 G8378 (.A1(W11450), .A2(W7487), .ZN(O7328));
  NOR2X1 G8379 (.A1(W15163), .A2(W1525), .ZN(O1155));
  NOR2X1 G8380 (.A1(W17308), .A2(W25881), .ZN(W34559));
  NOR2X1 G8381 (.A1(W12984), .A2(W24858), .ZN(O7541));
  NOR2X1 G8382 (.A1(W12204), .A2(W9654), .ZN(W16284));
  NOR2X1 G8383 (.A1(W6097), .A2(W16109), .ZN(W30877));
  NOR2X1 G8384 (.A1(W31363), .A2(W2590), .ZN(W34565));
  NOR2X1 G8385 (.A1(W3851), .A2(W19050), .ZN(O7330));
  NOR2X1 G8386 (.A1(W18178), .A2(W3076), .ZN(O7331));
  NOR2X1 G8387 (.A1(W19033), .A2(W13808), .ZN(W30869));
  NOR2X1 G8388 (.A1(W32460), .A2(W12704), .ZN(O7333));
  NOR2X1 G8389 (.A1(W2514), .A2(W42), .ZN(O7754));
  NOR2X1 G8390 (.A1(W5660), .A2(W12367), .ZN(O1007));
  NOR2X1 G8391 (.A1(W31831), .A2(W12127), .ZN(O7750));
  NOR2X1 G8392 (.A1(W1208), .A2(W19503), .ZN(O5405));
  NOR2X1 G8393 (.A1(W20273), .A2(W6547), .ZN(W35344));
  NOR2X1 G8394 (.A1(W14211), .A2(I764), .ZN(O1956));
  NOR2X1 G8395 (.A1(W6212), .A2(W2528), .ZN(W15448));
  NOR2X1 G8396 (.A1(W3050), .A2(W13766), .ZN(W15447));
  NOR2X1 G8397 (.A1(W9521), .A2(W5509), .ZN(W15446));
  NOR2X1 G8398 (.A1(W10338), .A2(W4192), .ZN(O1008));
  NOR2X1 G8399 (.A1(I1638), .A2(W12459), .ZN(W15444));
  NOR2X1 G8400 (.A1(W3569), .A2(W3655), .ZN(W15443));
  NOR2X1 G8401 (.A1(W9681), .A2(W12473), .ZN(W15442));
  NOR2X1 G8402 (.A1(W22681), .A2(W5184), .ZN(W30583));
  NOR2X1 G8403 (.A1(W15558), .A2(W4928), .ZN(O7756));
  NOR2X1 G8404 (.A1(W7658), .A2(I1139), .ZN(W30582));
  NOR2X1 G8405 (.A1(W2546), .A2(W1369), .ZN(W15438));
  NOR2X1 G8406 (.A1(W11845), .A2(W6753), .ZN(W15437));
  NOR2X1 G8407 (.A1(W8668), .A2(W15545), .ZN(O1954));
  NOR2X1 G8408 (.A1(W6912), .A2(W7230), .ZN(W15474));
  NOR2X1 G8409 (.A1(W216), .A2(W5994), .ZN(W20203));
  NOR2X1 G8410 (.A1(W7519), .A2(W10331), .ZN(W15472));
  NOR2X1 G8411 (.A1(W1177), .A2(W9667), .ZN(W35331));
  NOR2X1 G8412 (.A1(W28998), .A2(W30166), .ZN(O7743));
  NOR2X1 G8413 (.A1(W8261), .A2(W13300), .ZN(O1012));
  NOR2X1 G8414 (.A1(W8905), .A2(W13289), .ZN(W15467));
  NOR2X1 G8415 (.A1(W4629), .A2(W15782), .ZN(W35333));
  NOR2X1 G8416 (.A1(W13348), .A2(W8045), .ZN(W15436));
  NOR2X1 G8417 (.A1(W13718), .A2(W3910), .ZN(W15463));
  NOR2X1 G8418 (.A1(W13231), .A2(W1706), .ZN(W15462));
  NOR2X1 G8419 (.A1(W21363), .A2(W6613), .ZN(O7746));
  NOR2X1 G8420 (.A1(I365), .A2(W6442), .ZN(W30591));
  NOR2X1 G8421 (.A1(W9018), .A2(W5456), .ZN(W15459));
  NOR2X1 G8422 (.A1(W11584), .A2(W7956), .ZN(W15458));
  NOR2X1 G8423 (.A1(I188), .A2(W7768), .ZN(W20208));
  NOR2X1 G8424 (.A1(W1281), .A2(W14864), .ZN(W20226));
  NOR2X1 G8425 (.A1(W463), .A2(W6927), .ZN(W35369));
  NOR2X1 G8426 (.A1(W6880), .A2(W19367), .ZN(W20220));
  NOR2X1 G8427 (.A1(W11001), .A2(W18024), .ZN(W35371));
  NOR2X1 G8428 (.A1(W22002), .A2(W25137), .ZN(W35381));
  NOR2X1 G8429 (.A1(W7622), .A2(W14480), .ZN(O1001));
  NOR2X1 G8430 (.A1(W26483), .A2(W20883), .ZN(W30576));
  NOR2X1 G8431 (.A1(W16276), .A2(W18923), .ZN(O5400));
  NOR2X1 G8432 (.A1(W9557), .A2(W2044), .ZN(W15407));
  NOR2X1 G8433 (.A1(W4879), .A2(W9225), .ZN(W15418));
  NOR2X1 G8434 (.A1(W2964), .A2(W13951), .ZN(O7777));
  NOR2X1 G8435 (.A1(W4771), .A2(I778), .ZN(W15404));
  NOR2X1 G8436 (.A1(W4752), .A2(W13802), .ZN(W15403));
  NOR2X1 G8437 (.A1(W7225), .A2(W3910), .ZN(W15402));
  NOR2X1 G8438 (.A1(W5144), .A2(W6363), .ZN(O7778));
  NOR2X1 G8439 (.A1(W22494), .A2(W22617), .ZN(O7780));
  NOR2X1 G8440 (.A1(I744), .A2(W1581), .ZN(W20227));
  NOR2X1 G8441 (.A1(W4624), .A2(W31228), .ZN(W35400));
  NOR2X1 G8442 (.A1(W2921), .A2(W8525), .ZN(W15426));
  NOR2X1 G8443 (.A1(W16203), .A2(W8024), .ZN(W30581));
  NOR2X1 G8444 (.A1(W11630), .A2(W19631), .ZN(W20216));
  NOR2X1 G8445 (.A1(W10349), .A2(W3035), .ZN(W35360));
  NOR2X1 G8446 (.A1(W6871), .A2(I1541), .ZN(O1005));
  NOR2X1 G8447 (.A1(W1625), .A2(I1052), .ZN(W15431));
  NOR2X1 G8448 (.A1(W10522), .A2(W742), .ZN(W20218));
  NOR2X1 G8449 (.A1(W14457), .A2(W8625), .ZN(O7761));
  NOR2X1 G8450 (.A1(W3585), .A2(W6290), .ZN(W15427));
  NOR2X1 G8451 (.A1(I1476), .A2(W18465), .ZN(O7741));
  NOR2X1 G8452 (.A1(W29190), .A2(I1533), .ZN(O7762));
  NOR2X1 G8453 (.A1(W28748), .A2(I1421), .ZN(W30579));
  NOR2X1 G8454 (.A1(W9334), .A2(W14943), .ZN(O1004));
  NOR2X1 G8455 (.A1(W9800), .A2(W22198), .ZN(O7764));
  NOR2X1 G8456 (.A1(W8605), .A2(I266), .ZN(O1003));
  NOR2X1 G8457 (.A1(W28721), .A2(W8236), .ZN(W35367));
  NOR2X1 G8458 (.A1(W12792), .A2(W17685), .ZN(O7765));
  NOR2X1 G8459 (.A1(W14255), .A2(W19415), .ZN(O7716));
  NOR2X1 G8460 (.A1(W29276), .A2(W17699), .ZN(W30610));
  NOR2X1 G8461 (.A1(W17370), .A2(W11414), .ZN(W20192));
  NOR2X1 G8462 (.A1(W1714), .A2(W13894), .ZN(O1022));
  NOR2X1 G8463 (.A1(W8053), .A2(W13119), .ZN(O5414));
  NOR2X1 G8464 (.A1(W25778), .A2(W10713), .ZN(W35283));
  NOR2X1 G8465 (.A1(W25225), .A2(W21529), .ZN(W35285));
  NOR2X1 G8466 (.A1(W1288), .A2(W1413), .ZN(W15523));
  NOR2X1 G8467 (.A1(W198), .A2(W14620), .ZN(W15522));
  NOR2X1 G8468 (.A1(W576), .A2(W437), .ZN(W15532));
  NOR2X1 G8469 (.A1(W1421), .A2(W21825), .ZN(O5409));
  NOR2X1 G8470 (.A1(W18037), .A2(W27060), .ZN(O7719));
  NOR2X1 G8471 (.A1(W7360), .A2(W14615), .ZN(O7720));
  NOR2X1 G8472 (.A1(I297), .A2(W33781), .ZN(W35293));
  NOR2X1 G8473 (.A1(W1322), .A2(W14509), .ZN(W15515));
  NOR2X1 G8474 (.A1(W8288), .A2(W4150), .ZN(W15514));
  NOR2X1 G8475 (.A1(W19845), .A2(W17400), .ZN(O7721));
  NOR2X1 G8476 (.A1(I901), .A2(W11395), .ZN(O1019));
  NOR2X1 G8477 (.A1(W5382), .A2(W15379), .ZN(W15541));
  NOR2X1 G8478 (.A1(W31073), .A2(W29898), .ZN(O7701));
  NOR2X1 G8479 (.A1(W3095), .A2(W21130), .ZN(W30618));
  NOR2X1 G8480 (.A1(W24546), .A2(W22612), .ZN(W35264));
  NOR2X1 G8481 (.A1(W14748), .A2(W4373), .ZN(W15547));
  NOR2X1 G8482 (.A1(W2225), .A2(W9614), .ZN(W30615));
  NOR2X1 G8483 (.A1(W29743), .A2(W6096), .ZN(W35267));
  NOR2X1 G8484 (.A1(W11043), .A2(W9513), .ZN(W20186));
  NOR2X1 G8485 (.A1(W15128), .A2(W24986), .ZN(W35270));
  NOR2X1 G8486 (.A1(W676), .A2(W11836), .ZN(W15511));
  NOR2X1 G8487 (.A1(W3394), .A2(W14470), .ZN(O5415));
  NOR2X1 G8488 (.A1(W16636), .A2(I1211), .ZN(W30613));
  NOR2X1 G8489 (.A1(W10307), .A2(W13558), .ZN(O1025));
  NOR2X1 G8490 (.A1(I1877), .A2(W18973), .ZN(O7709));
  NOR2X1 G8491 (.A1(W8814), .A2(W15406), .ZN(W15535));
  NOR2X1 G8492 (.A1(W4540), .A2(W1578), .ZN(O7710));
  NOR2X1 G8493 (.A1(W12924), .A2(W24497), .ZN(W30611));
  NOR2X1 G8494 (.A1(W23075), .A2(W27725), .ZN(O7733));
  NOR2X1 G8495 (.A1(W4995), .A2(W13687), .ZN(W30598));
  NOR2X1 G8496 (.A1(W3211), .A2(I1542), .ZN(W15492));
  NOR2X1 G8497 (.A1(W13910), .A2(W21078), .ZN(W35308));
  NOR2X1 G8498 (.A1(W32531), .A2(W11490), .ZN(O7729));
  NOR2X1 G8499 (.A1(W6635), .A2(W12863), .ZN(W15489));
  NOR2X1 G8500 (.A1(W29385), .A2(W5116), .ZN(W30596));
  NOR2X1 G8501 (.A1(W10276), .A2(W3743), .ZN(O7730));
  NOR2X1 G8502 (.A1(W14846), .A2(W7360), .ZN(W15486));
  NOR2X1 G8503 (.A1(W11487), .A2(W9232), .ZN(W15494));
  NOR2X1 G8504 (.A1(W4277), .A2(W3053), .ZN(O1016));
  NOR2X1 G8505 (.A1(W21955), .A2(W11141), .ZN(O7735));
  NOR2X1 G8506 (.A1(W29612), .A2(W32132), .ZN(O7737));
  NOR2X1 G8507 (.A1(W10430), .A2(W30974), .ZN(O7738));
  NOR2X1 G8508 (.A1(W15202), .A2(W5061), .ZN(W15480));
  NOR2X1 G8509 (.A1(W27278), .A2(W29164), .ZN(O7739));
  NOR2X1 G8510 (.A1(W5247), .A2(W14205), .ZN(W15477));
  NOR2X1 G8511 (.A1(W12590), .A2(W10019), .ZN(W15476));
  NOR2X1 G8512 (.A1(W3174), .A2(I459), .ZN(W35300));
  NOR2X1 G8513 (.A1(W5888), .A2(W14293), .ZN(O1018));
  NOR2X1 G8514 (.A1(W8610), .A2(W3839), .ZN(W35295));
  NOR2X1 G8515 (.A1(W21987), .A2(W3291), .ZN(W30600));
  NOR2X1 G8516 (.A1(W28583), .A2(W26714), .ZN(O5408));
  NOR2X1 G8517 (.A1(W10183), .A2(W6728), .ZN(W15506));
  NOR2X1 G8518 (.A1(W20683), .A2(W13775), .ZN(W35298));
  NOR2X1 G8519 (.A1(W4528), .A2(W30165), .ZN(O7724));
  NOR2X1 G8520 (.A1(W6367), .A2(W3842), .ZN(O1017));
  NOR2X1 G8521 (.A1(W10115), .A2(W9842), .ZN(O1000));
  NOR2X1 G8522 (.A1(W27956), .A2(W2329), .ZN(W35301));
  NOR2X1 G8523 (.A1(I1116), .A2(W64), .ZN(O7725));
  NOR2X1 G8524 (.A1(W11920), .A2(W7483), .ZN(W15499));
  NOR2X1 G8525 (.A1(W12716), .A2(W8976), .ZN(W15498));
  NOR2X1 G8526 (.A1(W19706), .A2(W34746), .ZN(O7726));
  NOR2X1 G8527 (.A1(W393), .A2(W11646), .ZN(W15496));
  NOR2X1 G8528 (.A1(W2944), .A2(W16343), .ZN(O7727));
  NOR2X1 G8529 (.A1(W32630), .A2(W24306), .ZN(O7846));
  NOR2X1 G8530 (.A1(W10624), .A2(W3993), .ZN(W15300));
  NOR2X1 G8531 (.A1(W23345), .A2(W1328), .ZN(O7841));
  NOR2X1 G8532 (.A1(W4404), .A2(W12592), .ZN(W15298));
  NOR2X1 G8533 (.A1(W4627), .A2(W5713), .ZN(O988));
  NOR2X1 G8534 (.A1(W4432), .A2(W17528), .ZN(O7842));
  NOR2X1 G8535 (.A1(W11346), .A2(W20755), .ZN(O7843));
  NOR2X1 G8536 (.A1(W11144), .A2(W13692), .ZN(W15294));
  NOR2X1 G8537 (.A1(W212), .A2(W26532), .ZN(W35503));
  NOR2X1 G8538 (.A1(W14846), .A2(W8733), .ZN(O5388));
  NOR2X1 G8539 (.A1(W31989), .A2(W27565), .ZN(O7847));
  NOR2X1 G8540 (.A1(W10727), .A2(W20620), .ZN(O5387));
  NOR2X1 G8541 (.A1(W15332), .A2(W5500), .ZN(O1965));
  NOR2X1 G8542 (.A1(W16388), .A2(W6027), .ZN(W20258));
  NOR2X1 G8543 (.A1(W23348), .A2(W31160), .ZN(W35510));
  NOR2X1 G8544 (.A1(W16136), .A2(W6684), .ZN(O5384));
  NOR2X1 G8545 (.A1(W20847), .A2(W1475), .ZN(O7852));
  NOR2X1 G8546 (.A1(W27729), .A2(W32585), .ZN(W35515));
  NOR2X1 G8547 (.A1(W14796), .A2(W6462), .ZN(W15310));
  NOR2X1 G8548 (.A1(W2763), .A2(W785), .ZN(W15318));
  NOR2X1 G8549 (.A1(W9657), .A2(W9923), .ZN(O7826));
  NOR2X1 G8550 (.A1(W10521), .A2(W2211), .ZN(W15316));
  NOR2X1 G8551 (.A1(W21746), .A2(W25800), .ZN(W35482));
  NOR2X1 G8552 (.A1(W5615), .A2(W7653), .ZN(O1962));
  NOR2X1 G8553 (.A1(W10083), .A2(W112), .ZN(W15313));
  NOR2X1 G8554 (.A1(W9893), .A2(W13082), .ZN(W15312));
  NOR2X1 G8555 (.A1(W4094), .A2(W2477), .ZN(W15311));
  NOR2X1 G8556 (.A1(W13775), .A2(W9716), .ZN(W15281));
  NOR2X1 G8557 (.A1(W12261), .A2(W15028), .ZN(O7832));
  NOR2X1 G8558 (.A1(W10528), .A2(W12761), .ZN(W15308));
  NOR2X1 G8559 (.A1(W27986), .A2(W23213), .ZN(W35486));
  NOR2X1 G8560 (.A1(W3785), .A2(W5242), .ZN(W15306));
  NOR2X1 G8561 (.A1(W26209), .A2(W521), .ZN(O7838));
  NOR2X1 G8562 (.A1(W27893), .A2(W8273), .ZN(O5389));
  NOR2X1 G8563 (.A1(W14576), .A2(W6117), .ZN(W15302));
  NOR2X1 G8564 (.A1(W10222), .A2(W19018), .ZN(W30525));
  NOR2X1 G8565 (.A1(W5317), .A2(W11556), .ZN(O7867));
  NOR2X1 G8566 (.A1(W28182), .A2(W25261), .ZN(W30528));
  NOR2X1 G8567 (.A1(W18991), .A2(W29890), .ZN(O7869));
  NOR2X1 G8568 (.A1(W5910), .A2(W5370), .ZN(W20268));
  NOR2X1 G8569 (.A1(W31139), .A2(W34604), .ZN(W35547));
  NOR2X1 G8570 (.A1(W3490), .A2(W16450), .ZN(W20269));
  NOR2X1 G8571 (.A1(W4706), .A2(W20724), .ZN(W35551));
  NOR2X1 G8572 (.A1(W10138), .A2(W2540), .ZN(O979));
  NOR2X1 G8573 (.A1(W16285), .A2(W10599), .ZN(W20266));
  NOR2X1 G8574 (.A1(W4590), .A2(W135), .ZN(W15250));
  NOR2X1 G8575 (.A1(W12142), .A2(W10768), .ZN(O978));
  NOR2X1 G8576 (.A1(W1979), .A2(W14016), .ZN(W15247));
  NOR2X1 G8577 (.A1(W16321), .A2(W984), .ZN(W35556));
  NOR2X1 G8578 (.A1(W1423), .A2(W4817), .ZN(O7881));
  NOR2X1 G8579 (.A1(W22860), .A2(W2750), .ZN(O7882));
  NOR2X1 G8580 (.A1(W14472), .A2(W16880), .ZN(O5376));
  NOR2X1 G8581 (.A1(W9363), .A2(W16668), .ZN(O5375));
  NOR2X1 G8582 (.A1(W12309), .A2(W15205), .ZN(W35530));
  NOR2X1 G8583 (.A1(W2681), .A2(W6170), .ZN(W15280));
  NOR2X1 G8584 (.A1(W17804), .A2(W13379), .ZN(W20262));
  NOR2X1 G8585 (.A1(W18967), .A2(W6378), .ZN(O7858));
  NOR2X1 G8586 (.A1(W30244), .A2(W32263), .ZN(W35522));
  NOR2X1 G8587 (.A1(W7920), .A2(W10116), .ZN(W15274));
  NOR2X1 G8588 (.A1(W33575), .A2(W565), .ZN(O7859));
  NOR2X1 G8589 (.A1(W5400), .A2(W12378), .ZN(W35526));
  NOR2X1 G8590 (.A1(W25528), .A2(W14962), .ZN(W35528));
  NOR2X1 G8591 (.A1(W11274), .A2(W22179), .ZN(W35475));
  NOR2X1 G8592 (.A1(W1358), .A2(W495), .ZN(W15268));
  NOR2X1 G8593 (.A1(W23076), .A2(W21119), .ZN(O5381));
  NOR2X1 G8594 (.A1(W15938), .A2(W16281), .ZN(O7862));
  NOR2X1 G8595 (.A1(W14170), .A2(I193), .ZN(O5380));
  NOR2X1 G8596 (.A1(W34866), .A2(W13961), .ZN(O7864));
  NOR2X1 G8597 (.A1(W35234), .A2(W8731), .ZN(O7865));
  NOR2X1 G8598 (.A1(W8056), .A2(W20227), .ZN(O7866));
  NOR2X1 G8599 (.A1(W24515), .A2(W22617), .ZN(W35429));
  NOR2X1 G8600 (.A1(W32055), .A2(W769), .ZN(W35421));
  NOR2X1 G8601 (.A1(W21544), .A2(W9685), .ZN(W35422));
  NOR2X1 G8602 (.A1(W9379), .A2(I1860), .ZN(O7797));
  NOR2X1 G8603 (.A1(W6649), .A2(W5848), .ZN(W15375));
  NOR2X1 G8604 (.A1(W12413), .A2(W710), .ZN(W15374));
  NOR2X1 G8605 (.A1(W14292), .A2(W4450), .ZN(W35426));
  NOR2X1 G8606 (.A1(W108), .A2(W5723), .ZN(W15371));
  NOR2X1 G8607 (.A1(I1200), .A2(W13509), .ZN(W15370));
  NOR2X1 G8608 (.A1(W13921), .A2(W13546), .ZN(W15379));
  NOR2X1 G8609 (.A1(W24302), .A2(W24016), .ZN(W35431));
  NOR2X1 G8610 (.A1(W10661), .A2(W4459), .ZN(W20234));
  NOR2X1 G8611 (.A1(W33870), .A2(W17647), .ZN(W35433));
  NOR2X1 G8612 (.A1(I1520), .A2(W11264), .ZN(W15364));
  NOR2X1 G8613 (.A1(W3470), .A2(W6095), .ZN(W15363));
  NOR2X1 G8614 (.A1(W4630), .A2(W13897), .ZN(W15362));
  NOR2X1 G8615 (.A1(W8101), .A2(W13003), .ZN(W15360));
  NOR2X1 G8616 (.A1(W12331), .A2(W25254), .ZN(O7803));
  NOR2X1 G8617 (.A1(W8177), .A2(W23026), .ZN(O7793));
  NOR2X1 G8618 (.A1(W7400), .A2(W5740), .ZN(W15396));
  NOR2X1 G8619 (.A1(W8882), .A2(W5506), .ZN(W15395));
  NOR2X1 G8620 (.A1(W9171), .A2(W8825), .ZN(O7783));
  NOR2X1 G8621 (.A1(I1103), .A2(W7715), .ZN(O7787));
  NOR2X1 G8622 (.A1(W4311), .A2(W10048), .ZN(O1957));
  NOR2X1 G8623 (.A1(W16420), .A2(W25720), .ZN(O7791));
  NOR2X1 G8624 (.A1(W9428), .A2(W19456), .ZN(O7792));
  NOR2X1 G8625 (.A1(W4267), .A2(W14146), .ZN(W15388));
  NOR2X1 G8626 (.A1(W13316), .A2(W14884), .ZN(O7804));
  NOR2X1 G8627 (.A1(I43), .A2(W15362), .ZN(O998));
  NOR2X1 G8628 (.A1(W7661), .A2(W1299), .ZN(O5398));
  NOR2X1 G8629 (.A1(W19190), .A2(W31616), .ZN(W35415));
  NOR2X1 G8630 (.A1(I0), .A2(W7747), .ZN(W15383));
  NOR2X1 G8631 (.A1(W7378), .A2(W6944), .ZN(W20231));
  NOR2X1 G8632 (.A1(W29287), .A2(W3721), .ZN(W35417));
  NOR2X1 G8633 (.A1(W3686), .A2(W20459), .ZN(W35420));
  NOR2X1 G8634 (.A1(W5645), .A2(W6529), .ZN(O1961));
  NOR2X1 G8635 (.A1(W715), .A2(W3037), .ZN(O1960));
  NOR2X1 G8636 (.A1(W1040), .A2(W3014), .ZN(W15336));
  NOR2X1 G8637 (.A1(I1431), .A2(W636), .ZN(O993));
  NOR2X1 G8638 (.A1(W34791), .A2(W22789), .ZN(O7819));
  NOR2X1 G8639 (.A1(W12892), .A2(W29622), .ZN(O5392));
  NOR2X1 G8640 (.A1(W14329), .A2(W14691), .ZN(W15332));
  NOR2X1 G8641 (.A1(W198), .A2(W11004), .ZN(W20245));
  NOR2X1 G8642 (.A1(W6186), .A2(W10685), .ZN(W15330));
  NOR2X1 G8643 (.A1(W16260), .A2(W4631), .ZN(W35459));
  NOR2X1 G8644 (.A1(I246), .A2(W5006), .ZN(W15327));
  NOR2X1 G8645 (.A1(I289), .A2(W12830), .ZN(W15326));
  NOR2X1 G8646 (.A1(W12064), .A2(W27512), .ZN(O5390));
  NOR2X1 G8647 (.A1(W13318), .A2(W8997), .ZN(W15324));
  NOR2X1 G8648 (.A1(W4806), .A2(W31154), .ZN(O7821));
  NOR2X1 G8649 (.A1(W6506), .A2(W10803), .ZN(W15322));
  NOR2X1 G8650 (.A1(W19620), .A2(W18726), .ZN(W20249));
  NOR2X1 G8651 (.A1(W8927), .A2(W9620), .ZN(W15320));
  NOR2X1 G8652 (.A1(W8407), .A2(W9339), .ZN(O7812));
  NOR2X1 G8653 (.A1(W12949), .A2(W11176), .ZN(O7805));
  NOR2X1 G8654 (.A1(W12994), .A2(W13992), .ZN(W35440));
  NOR2X1 G8655 (.A1(W4548), .A2(W848), .ZN(W15355));
  NOR2X1 G8656 (.A1(W9249), .A2(W2228), .ZN(W15354));
  NOR2X1 G8657 (.A1(W1465), .A2(W11777), .ZN(W15353));
  NOR2X1 G8658 (.A1(W17142), .A2(W30618), .ZN(O7810));
  NOR2X1 G8659 (.A1(W2216), .A2(W2689), .ZN(W30556));
  NOR2X1 G8660 (.A1(W881), .A2(W28615), .ZN(W30555));
  NOR2X1 G8661 (.A1(W20189), .A2(W29664), .ZN(O5416));
  NOR2X1 G8662 (.A1(W35181), .A2(W27211), .ZN(O7813));
  NOR2X1 G8663 (.A1(W5417), .A2(W3142), .ZN(W20241));
  NOR2X1 G8664 (.A1(W19556), .A2(W25594), .ZN(O5393));
  NOR2X1 G8665 (.A1(W4397), .A2(W19417), .ZN(W35456));
  NOR2X1 G8666 (.A1(W22808), .A2(W19655), .ZN(W35457));
  NOR2X1 G8667 (.A1(W13959), .A2(W2397), .ZN(W15340));
  NOR2X1 G8668 (.A1(W29730), .A2(W14927), .ZN(O7815));
  NOR2X1 G8669 (.A1(W5742), .A2(W11470), .ZN(O7607));
  NOR2X1 G8670 (.A1(W9340), .A2(W9432), .ZN(W30685));
  NOR2X1 G8671 (.A1(W3557), .A2(W3316), .ZN(W35065));
  NOR2X1 G8672 (.A1(W13617), .A2(W14872), .ZN(W15757));
  NOR2X1 G8673 (.A1(W5117), .A2(W9330), .ZN(O7604));
  NOR2X1 G8674 (.A1(W17723), .A2(W21704), .ZN(O7606));
  NOR2X1 G8675 (.A1(W21670), .A2(W16367), .ZN(W35069));
  NOR2X1 G8676 (.A1(W6089), .A2(W9338), .ZN(W15753));
  NOR2X1 G8677 (.A1(W19010), .A2(W11346), .ZN(W35070));
  NOR2X1 G8678 (.A1(I1151), .A2(I235), .ZN(W15760));
  NOR2X1 G8679 (.A1(W9749), .A2(W3571), .ZN(W20116));
  NOR2X1 G8680 (.A1(W364), .A2(W3316), .ZN(W35076));
  NOR2X1 G8681 (.A1(W33021), .A2(W9419), .ZN(O7612));
  NOR2X1 G8682 (.A1(W17370), .A2(W3984), .ZN(W30679));
  NOR2X1 G8683 (.A1(W2358), .A2(W13883), .ZN(O1060));
  NOR2X1 G8684 (.A1(W22463), .A2(I1322), .ZN(O7614));
  NOR2X1 G8685 (.A1(W33695), .A2(W8973), .ZN(O7615));
  NOR2X1 G8686 (.A1(W6361), .A2(W664), .ZN(W15742));
  NOR2X1 G8687 (.A1(W5119), .A2(W11891), .ZN(W15770));
  NOR2X1 G8688 (.A1(W15714), .A2(W13516), .ZN(O1928));
  NOR2X1 G8689 (.A1(W17704), .A2(W5187), .ZN(W30697));
  NOR2X1 G8690 (.A1(I435), .A2(W11097), .ZN(W15776));
  NOR2X1 G8691 (.A1(W7756), .A2(W9247), .ZN(W20108));
  NOR2X1 G8692 (.A1(W35021), .A2(W19807), .ZN(W35050));
  NOR2X1 G8693 (.A1(W11165), .A2(W34730), .ZN(O7594));
  NOR2X1 G8694 (.A1(W3512), .A2(W1218), .ZN(W35053));
  NOR2X1 G8695 (.A1(W5346), .A2(W10535), .ZN(W20109));
  NOR2X1 G8696 (.A1(W11966), .A2(W9782), .ZN(O1929));
  NOR2X1 G8697 (.A1(W27972), .A2(W6876), .ZN(O7597));
  NOR2X1 G8698 (.A1(W3100), .A2(W14550), .ZN(O5455));
  NOR2X1 G8699 (.A1(W2187), .A2(W16663), .ZN(O5453));
  NOR2X1 G8700 (.A1(W8012), .A2(W13973), .ZN(W20112));
  NOR2X1 G8701 (.A1(W12637), .A2(W20188), .ZN(O7601));
  NOR2X1 G8702 (.A1(W12520), .A2(W10057), .ZN(W15764));
  NOR2X1 G8703 (.A1(W11026), .A2(W9004), .ZN(W15763));
  NOR2X1 G8704 (.A1(W13035), .A2(W7418), .ZN(W15711));
  NOR2X1 G8705 (.A1(W2577), .A2(W4781), .ZN(W15723));
  NOR2X1 G8706 (.A1(W28671), .A2(W15978), .ZN(W35096));
  NOR2X1 G8707 (.A1(W2167), .A2(W24490), .ZN(W35098));
  NOR2X1 G8708 (.A1(W26196), .A2(I786), .ZN(O5446));
  NOR2X1 G8709 (.A1(W13499), .A2(W5565), .ZN(W20128));
  NOR2X1 G8710 (.A1(I230), .A2(W21578), .ZN(O7628));
  NOR2X1 G8711 (.A1(W4642), .A2(W9769), .ZN(O1054));
  NOR2X1 G8712 (.A1(W7310), .A2(W4505), .ZN(O7629));
  NOR2X1 G8713 (.A1(W26201), .A2(W10697), .ZN(O7621));
  NOR2X1 G8714 (.A1(W10495), .A2(W18937), .ZN(O7630));
  NOR2X1 G8715 (.A1(W6838), .A2(W3064), .ZN(W15709));
  NOR2X1 G8716 (.A1(W31172), .A2(W19686), .ZN(O7631));
  NOR2X1 G8717 (.A1(W9289), .A2(W3705), .ZN(W15707));
  NOR2X1 G8718 (.A1(W16774), .A2(W16563), .ZN(W20130));
  NOR2X1 G8719 (.A1(W7171), .A2(W1866), .ZN(O7633));
  NOR2X1 G8720 (.A1(I875), .A2(W10717), .ZN(W15704));
  NOR2X1 G8721 (.A1(W4336), .A2(W2822), .ZN(W15703));
  NOR2X1 G8722 (.A1(W7901), .A2(I1746), .ZN(O1057));
  NOR2X1 G8723 (.A1(W1682), .A2(W13024), .ZN(W15740));
  NOR2X1 G8724 (.A1(W15790), .A2(W11704), .ZN(O1930));
  NOR2X1 G8725 (.A1(W7690), .A2(W2212), .ZN(O1058));
  NOR2X1 G8726 (.A1(W11868), .A2(W11586), .ZN(O1931));
  NOR2X1 G8727 (.A1(W5383), .A2(W29447), .ZN(O5449));
  NOR2X1 G8728 (.A1(W10441), .A2(W20489), .ZN(O5447));
  NOR2X1 G8729 (.A1(W15426), .A2(W8201), .ZN(W35089));
  NOR2X1 G8730 (.A1(W22205), .A2(W30971), .ZN(W35090));
  NOR2X1 G8731 (.A1(W14321), .A2(W11205), .ZN(W15779));
  NOR2X1 G8732 (.A1(W6089), .A2(W4091), .ZN(W15731));
  NOR2X1 G8733 (.A1(W686), .A2(I1424), .ZN(W15730));
  NOR2X1 G8734 (.A1(W7797), .A2(W518), .ZN(O7618));
  NOR2X1 G8735 (.A1(W13825), .A2(W30402), .ZN(W35092));
  NOR2X1 G8736 (.A1(W10299), .A2(W1110), .ZN(W15727));
  NOR2X1 G8737 (.A1(W5821), .A2(W315), .ZN(O7619));
  NOR2X1 G8738 (.A1(W32720), .A2(W13974), .ZN(O7620));
  NOR2X1 G8739 (.A1(W20695), .A2(W9827), .ZN(W34992));
  NOR2X1 G8740 (.A1(W1349), .A2(W19167), .ZN(O7553));
  NOR2X1 G8741 (.A1(W3098), .A2(W4297), .ZN(W15838));
  NOR2X1 G8742 (.A1(W14757), .A2(W14535), .ZN(O1073));
  NOR2X1 G8743 (.A1(W12486), .A2(W11917), .ZN(W15836));
  NOR2X1 G8744 (.A1(W8370), .A2(W942), .ZN(W30728));
  NOR2X1 G8745 (.A1(W3687), .A2(W1892), .ZN(W15834));
  NOR2X1 G8746 (.A1(W19101), .A2(I842), .ZN(O7555));
  NOR2X1 G8747 (.A1(W10559), .A2(W2821), .ZN(W15831));
  NOR2X1 G8748 (.A1(W11202), .A2(W6666), .ZN(O7552));
  NOR2X1 G8749 (.A1(W12080), .A2(W21385), .ZN(O7560));
  NOR2X1 G8750 (.A1(W34378), .A2(W27346), .ZN(O7561));
  NOR2X1 G8751 (.A1(W12879), .A2(W7498), .ZN(W15827));
  NOR2X1 G8752 (.A1(W26495), .A2(W3879), .ZN(O7562));
  NOR2X1 G8753 (.A1(W1653), .A2(W12935), .ZN(W15825));
  NOR2X1 G8754 (.A1(W4532), .A2(W4504), .ZN(W15824));
  NOR2X1 G8755 (.A1(W10920), .A2(W19698), .ZN(W30725));
  NOR2X1 G8756 (.A1(W11350), .A2(W24672), .ZN(O7563));
  NOR2X1 G8757 (.A1(W14158), .A2(W33418), .ZN(O7546));
  NOR2X1 G8758 (.A1(W17775), .A2(W31841), .ZN(O7542));
  NOR2X1 G8759 (.A1(W4193), .A2(W15066), .ZN(W15855));
  NOR2X1 G8760 (.A1(W18505), .A2(W15135), .ZN(O1922));
  NOR2X1 G8761 (.A1(W14004), .A2(W31724), .ZN(O7543));
  NOR2X1 G8762 (.A1(W12858), .A2(W16456), .ZN(W20082));
  NOR2X1 G8763 (.A1(W14438), .A2(W26819), .ZN(O7545));
  NOR2X1 G8764 (.A1(W26506), .A2(W12431), .ZN(W34974));
  NOR2X1 G8765 (.A1(W7607), .A2(W1918), .ZN(W15849));
  NOR2X1 G8766 (.A1(W6097), .A2(W10555), .ZN(W15821));
  NOR2X1 G8767 (.A1(W2937), .A2(W10252), .ZN(O1074));
  NOR2X1 G8768 (.A1(W15417), .A2(W10070), .ZN(W15846));
  NOR2X1 G8769 (.A1(W20090), .A2(W11972), .ZN(O7547));
  NOR2X1 G8770 (.A1(W110), .A2(W20431), .ZN(O7550));
  NOR2X1 G8771 (.A1(W10181), .A2(W23838), .ZN(W30729));
  NOR2X1 G8772 (.A1(W2304), .A2(W10650), .ZN(W15842));
  NOR2X1 G8773 (.A1(W12175), .A2(W14694), .ZN(W15841));
  NOR2X1 G8774 (.A1(W732), .A2(W5601), .ZN(W15791));
  NOR2X1 G8775 (.A1(W27421), .A2(W25285), .ZN(W30716));
  NOR2X1 G8776 (.A1(W21925), .A2(W26485), .ZN(W30713));
  NOR2X1 G8777 (.A1(W13922), .A2(W26135), .ZN(O5460));
  NOR2X1 G8778 (.A1(W2438), .A2(I610), .ZN(W15798));
  NOR2X1 G8779 (.A1(W28023), .A2(W17345), .ZN(W35028));
  NOR2X1 G8780 (.A1(W8446), .A2(W14662), .ZN(W15795));
  NOR2X1 G8781 (.A1(W7592), .A2(I38), .ZN(W15794));
  NOR2X1 G8782 (.A1(W14724), .A2(W24289), .ZN(W35030));
  NOR2X1 G8783 (.A1(W8015), .A2(W3619), .ZN(W15802));
  NOR2X1 G8784 (.A1(W2275), .A2(W14711), .ZN(W15790));
  NOR2X1 G8785 (.A1(W10982), .A2(I1835), .ZN(O7585));
  NOR2X1 G8786 (.A1(W7275), .A2(W15414), .ZN(O5459));
  NOR2X1 G8787 (.A1(W28588), .A2(I480), .ZN(W30705));
  NOR2X1 G8788 (.A1(W1958), .A2(W14657), .ZN(W15785));
  NOR2X1 G8789 (.A1(I206), .A2(W1515), .ZN(W20102));
  NOR2X1 G8790 (.A1(W32903), .A2(W13914), .ZN(O7588));
  NOR2X1 G8791 (.A1(W7569), .A2(W3987), .ZN(W30701));
  NOR2X1 G8792 (.A1(W32183), .A2(W6536), .ZN(W35011));
  NOR2X1 G8793 (.A1(W23125), .A2(W31711), .ZN(O7564));
  NOR2X1 G8794 (.A1(W6906), .A2(W9350), .ZN(O1925));
  NOR2X1 G8795 (.A1(W14597), .A2(W13237), .ZN(W15818));
  NOR2X1 G8796 (.A1(W5274), .A2(W12354), .ZN(W20088));
  NOR2X1 G8797 (.A1(W24710), .A2(W19810), .ZN(O7567));
  NOR2X1 G8798 (.A1(W4528), .A2(W8479), .ZN(W15815));
  NOR2X1 G8799 (.A1(W13571), .A2(W9231), .ZN(W15813));
  NOR2X1 G8800 (.A1(I1536), .A2(W2328), .ZN(W15811));
  NOR2X1 G8801 (.A1(W9774), .A2(W205), .ZN(O1053));
  NOR2X1 G8802 (.A1(W31191), .A2(W13209), .ZN(W35012));
  NOR2X1 G8803 (.A1(I698), .A2(W21971), .ZN(W30718));
  NOR2X1 G8804 (.A1(W11232), .A2(W6451), .ZN(O5462));
  NOR2X1 G8805 (.A1(W20505), .A2(W23097), .ZN(O7576));
  NOR2X1 G8806 (.A1(W1791), .A2(W18949), .ZN(W20093));
  NOR2X1 G8807 (.A1(W8721), .A2(W33122), .ZN(O7577));
  NOR2X1 G8808 (.A1(W14850), .A2(W2615), .ZN(O7578));
  NOR2X1 G8809 (.A1(W14351), .A2(W10307), .ZN(W15596));
  NOR2X1 G8810 (.A1(W8254), .A2(W5987), .ZN(W30635));
  NOR2X1 G8811 (.A1(W24666), .A2(W22968), .ZN(W35209));
  NOR2X1 G8812 (.A1(W11447), .A2(W4077), .ZN(O5422));
  NOR2X1 G8813 (.A1(W2554), .A2(I1141), .ZN(W15601));
  NOR2X1 G8814 (.A1(W10650), .A2(W14007), .ZN(W20169));
  NOR2X1 G8815 (.A1(W10643), .A2(W1825), .ZN(W15599));
  NOR2X1 G8816 (.A1(W1918), .A2(W15415), .ZN(W15598));
  NOR2X1 G8817 (.A1(W3082), .A2(W24080), .ZN(O7680));
  NOR2X1 G8818 (.A1(W11847), .A2(W8522), .ZN(W35206));
  NOR2X1 G8819 (.A1(W32194), .A2(W12416), .ZN(W35214));
  NOR2X1 G8820 (.A1(W20451), .A2(W24166), .ZN(W30633));
  NOR2X1 G8821 (.A1(W9132), .A2(W18456), .ZN(O7681));
  NOR2X1 G8822 (.A1(W17179), .A2(W25999), .ZN(O7682));
  NOR2X1 G8823 (.A1(W14976), .A2(W28183), .ZN(W35222));
  NOR2X1 G8824 (.A1(I540), .A2(W405), .ZN(W15590));
  NOR2X1 G8825 (.A1(W3766), .A2(W2949), .ZN(W15589));
  NOR2X1 G8826 (.A1(W13254), .A2(I145), .ZN(W15588));
  NOR2X1 G8827 (.A1(W1080), .A2(W9015), .ZN(W15614));
  NOR2X1 G8828 (.A1(W17304), .A2(W8303), .ZN(O1943));
  NOR2X1 G8829 (.A1(W16871), .A2(W34435), .ZN(W35196));
  NOR2X1 G8830 (.A1(I774), .A2(W3897), .ZN(O1944));
  NOR2X1 G8831 (.A1(W14504), .A2(W191), .ZN(O5424));
  NOR2X1 G8832 (.A1(W10263), .A2(W15236), .ZN(W15618));
  NOR2X1 G8833 (.A1(W15367), .A2(W7960), .ZN(O1038));
  NOR2X1 G8834 (.A1(W16015), .A2(W30946), .ZN(W35201));
  NOR2X1 G8835 (.A1(W13479), .A2(W19113), .ZN(O7675));
  NOR2X1 G8836 (.A1(W19383), .A2(W3640), .ZN(O7684));
  NOR2X1 G8837 (.A1(W4023), .A2(W12242), .ZN(W15613));
  NOR2X1 G8838 (.A1(W10621), .A2(W15884), .ZN(W35203));
  NOR2X1 G8839 (.A1(W9249), .A2(W8625), .ZN(W15610));
  NOR2X1 G8840 (.A1(W8127), .A2(W3079), .ZN(O1035));
  NOR2X1 G8841 (.A1(W23460), .A2(W28947), .ZN(O7676));
  NOR2X1 G8842 (.A1(W10346), .A2(W4616), .ZN(W15607));
  NOR2X1 G8843 (.A1(W6763), .A2(I693), .ZN(W15606));
  NOR2X1 G8844 (.A1(W26768), .A2(W6973), .ZN(W35251));
  NOR2X1 G8845 (.A1(W27055), .A2(W16586), .ZN(W35238));
  NOR2X1 G8846 (.A1(W24109), .A2(W22038), .ZN(O7691));
  NOR2X1 G8847 (.A1(W17323), .A2(W18686), .ZN(W35242));
  NOR2X1 G8848 (.A1(W25370), .A2(W17097), .ZN(O5421));
  NOR2X1 G8849 (.A1(I1318), .A2(W10891), .ZN(W30627));
  NOR2X1 G8850 (.A1(W34899), .A2(W27057), .ZN(O7693));
  NOR2X1 G8851 (.A1(W7120), .A2(W22494), .ZN(W35249));
  NOR2X1 G8852 (.A1(W19085), .A2(W1874), .ZN(O7695));
  NOR2X1 G8853 (.A1(I300), .A2(W33173), .ZN(W35236));
  NOR2X1 G8854 (.A1(W29002), .A2(W25430), .ZN(O5419));
  NOR2X1 G8855 (.A1(W12359), .A2(W7340), .ZN(W30622));
  NOR2X1 G8856 (.A1(W4231), .A2(W20213), .ZN(O7698));
  NOR2X1 G8857 (.A1(W13935), .A2(W8076), .ZN(W15556));
  NOR2X1 G8858 (.A1(W3173), .A2(W25376), .ZN(O5417));
  NOR2X1 G8859 (.A1(W33010), .A2(W22920), .ZN(O7700));
  NOR2X1 G8860 (.A1(W2850), .A2(W8774), .ZN(O1028));
  NOR2X1 G8861 (.A1(W25021), .A2(W1711), .ZN(W35259));
  NOR2X1 G8862 (.A1(W4076), .A2(W8181), .ZN(W20174));
  NOR2X1 G8863 (.A1(W8203), .A2(W3890), .ZN(W15586));
  NOR2X1 G8864 (.A1(W20692), .A2(W18206), .ZN(W30632));
  NOR2X1 G8865 (.A1(W11258), .A2(W9063), .ZN(W15584));
  NOR2X1 G8866 (.A1(W3245), .A2(W18822), .ZN(W20172));
  NOR2X1 G8867 (.A1(W8388), .A2(W4272), .ZN(W15582));
  NOR2X1 G8868 (.A1(W13064), .A2(W9818), .ZN(W15581));
  NOR2X1 G8869 (.A1(W20687), .A2(W6404), .ZN(W30630));
  NOR2X1 G8870 (.A1(W8426), .A2(W12385), .ZN(W15579));
  NOR2X1 G8871 (.A1(W12711), .A2(W6813), .ZN(W15624));
  NOR2X1 G8872 (.A1(W33858), .A2(W13537), .ZN(W35230));
  NOR2X1 G8873 (.A1(W14272), .A2(W16616), .ZN(O7686));
  NOR2X1 G8874 (.A1(W435), .A2(W10995), .ZN(W20175));
  NOR2X1 G8875 (.A1(W17909), .A2(W17756), .ZN(W35235));
  NOR2X1 G8876 (.A1(W5096), .A2(W450), .ZN(W15573));
  NOR2X1 G8877 (.A1(W15188), .A2(W8023), .ZN(O1030));
  NOR2X1 G8878 (.A1(W11698), .A2(W11523), .ZN(O1029));
  NOR2X1 G8879 (.A1(W12531), .A2(W26345), .ZN(W30662));
  NOR2X1 G8880 (.A1(W5070), .A2(W11689), .ZN(W15682));
  NOR2X1 G8881 (.A1(W25137), .A2(W17879), .ZN(O5440));
  NOR2X1 G8882 (.A1(W13984), .A2(W15588), .ZN(W15680));
  NOR2X1 G8883 (.A1(W7436), .A2(W22904), .ZN(W35135));
  NOR2X1 G8884 (.A1(W14639), .A2(W5712), .ZN(O7644));
  NOR2X1 G8885 (.A1(W16000), .A2(W31317), .ZN(O7645));
  NOR2X1 G8886 (.A1(W6653), .A2(W12071), .ZN(W30663));
  NOR2X1 G8887 (.A1(W15443), .A2(W12510), .ZN(W15675));
  NOR2X1 G8888 (.A1(W8704), .A2(W9842), .ZN(W20138));
  NOR2X1 G8889 (.A1(W31740), .A2(W557), .ZN(W35140));
  NOR2X1 G8890 (.A1(W24655), .A2(W26067), .ZN(W35141));
  NOR2X1 G8891 (.A1(W32442), .A2(W6345), .ZN(W35143));
  NOR2X1 G8892 (.A1(W1845), .A2(W29573), .ZN(W30661));
  NOR2X1 G8893 (.A1(W13535), .A2(W28462), .ZN(W35145));
  NOR2X1 G8894 (.A1(W10027), .A2(W11132), .ZN(W20143));
  NOR2X1 G8895 (.A1(W24928), .A2(W26822), .ZN(O5439));
  NOR2X1 G8896 (.A1(I941), .A2(I1365), .ZN(W15666));
  NOR2X1 G8897 (.A1(W29861), .A2(W3090), .ZN(W35125));
  NOR2X1 G8898 (.A1(W3526), .A2(W10270), .ZN(O1935));
  NOR2X1 G8899 (.A1(W14692), .A2(W29117), .ZN(W35117));
  NOR2X1 G8900 (.A1(W11907), .A2(W2074), .ZN(W15699));
  NOR2X1 G8901 (.A1(I162), .A2(W12703), .ZN(W15698));
  NOR2X1 G8902 (.A1(W21436), .A2(W33455), .ZN(O7635));
  NOR2X1 G8903 (.A1(W14449), .A2(W1856), .ZN(W20133));
  NOR2X1 G8904 (.A1(I1464), .A2(W27230), .ZN(O5442));
  NOR2X1 G8905 (.A1(W11261), .A2(W11052), .ZN(O7641));
  NOR2X1 G8906 (.A1(W1660), .A2(W19965), .ZN(O1939));
  NOR2X1 G8907 (.A1(W3810), .A2(W12929), .ZN(W20135));
  NOR2X1 G8908 (.A1(W32904), .A2(W3150), .ZN(O7643));
  NOR2X1 G8909 (.A1(W2665), .A2(W26715), .ZN(O5441));
  NOR2X1 G8910 (.A1(W14316), .A2(W3482), .ZN(W15687));
  NOR2X1 G8911 (.A1(W4958), .A2(W7438), .ZN(W15686));
  NOR2X1 G8912 (.A1(W8337), .A2(W32303), .ZN(W35131));
  NOR2X1 G8913 (.A1(W27041), .A2(W1875), .ZN(W35132));
  NOR2X1 G8914 (.A1(W17934), .A2(W7648), .ZN(O5429));
  NOR2X1 G8915 (.A1(W847), .A2(W1010), .ZN(W35173));
  NOR2X1 G8916 (.A1(W3979), .A2(W8757), .ZN(W15643));
  NOR2X1 G8917 (.A1(W17703), .A2(W17728), .ZN(W35175));
  NOR2X1 G8918 (.A1(W22518), .A2(W22223), .ZN(O5431));
  NOR2X1 G8919 (.A1(W15298), .A2(W34366), .ZN(O7664));
  NOR2X1 G8920 (.A1(W19442), .A2(W12910), .ZN(W35182));
  NOR2X1 G8921 (.A1(W18919), .A2(W6260), .ZN(O7665));
  NOR2X1 G8922 (.A1(W12608), .A2(W8137), .ZN(W15635));
  NOR2X1 G8923 (.A1(W7988), .A2(W11890), .ZN(O5433));
  NOR2X1 G8924 (.A1(W28227), .A2(W4239), .ZN(O5427));
  NOR2X1 G8925 (.A1(W8397), .A2(W10791), .ZN(W20160));
  NOR2X1 G8926 (.A1(W22628), .A2(W23579), .ZN(O7669));
  NOR2X1 G8927 (.A1(I1760), .A2(W27410), .ZN(W35189));
  NOR2X1 G8928 (.A1(W8364), .A2(I1783), .ZN(O7670));
  NOR2X1 G8929 (.A1(W10487), .A2(W6080), .ZN(W15627));
  NOR2X1 G8930 (.A1(I1019), .A2(W63), .ZN(W15625));
  NOR2X1 G8931 (.A1(W35076), .A2(W26106), .ZN(O7651));
  NOR2X1 G8932 (.A1(W14897), .A2(W7285), .ZN(W15664));
  NOR2X1 G8933 (.A1(W27786), .A2(W24864), .ZN(W35149));
  NOR2X1 G8934 (.A1(W3357), .A2(W33316), .ZN(O7649));
  NOR2X1 G8935 (.A1(W2900), .A2(W5962), .ZN(O1046));
  NOR2X1 G8936 (.A1(W17689), .A2(W19562), .ZN(O7650));
  NOR2X1 G8937 (.A1(W6209), .A2(W4549), .ZN(W15659));
  NOR2X1 G8938 (.A1(W12783), .A2(W12493), .ZN(W15657));
  NOR2X1 G8939 (.A1(W8821), .A2(W17620), .ZN(W35156));
  NOR2X1 G8940 (.A1(W9966), .A2(W10350), .ZN(O2432));
  NOR2X1 G8941 (.A1(W3406), .A2(W2062), .ZN(O5438));
  NOR2X1 G8942 (.A1(W7609), .A2(W162), .ZN(W15653));
  NOR2X1 G8943 (.A1(W16302), .A2(W3283), .ZN(O5437));
  NOR2X1 G8944 (.A1(W8928), .A2(W7132), .ZN(O7655));
  NOR2X1 G8945 (.A1(W815), .A2(W16148), .ZN(W20149));
  NOR2X1 G8946 (.A1(W6949), .A2(W15699), .ZN(O7657));
  NOR2X1 G8947 (.A1(W5826), .A2(W14058), .ZN(O5435));
  NOR2X1 G8948 (.A1(W159), .A2(I288), .ZN(O32));
  NOR2X1 G8949 (.A1(W31912), .A2(W24140), .ZN(O16575));
  NOR2X1 G8950 (.A1(W19850), .A2(W9347), .ZN(O3778));
  NOR2X1 G8951 (.A1(W2501), .A2(I1830), .ZN(W3342));
  NOR2X1 G8952 (.A1(W15815), .A2(W15350), .ZN(O3012));
  NOR2X1 G8953 (.A1(W11846), .A2(W32748), .ZN(O16578));
  NOR2X1 G8954 (.A1(I662), .A2(I762), .ZN(W3338));
  NOR2X1 G8955 (.A1(W35620), .A2(W3220), .ZN(O16579));
  NOR2X1 G8956 (.A1(W9749), .A2(W22154), .ZN(O3013));
  NOR2X1 G8957 (.A1(W19757), .A2(W37570), .ZN(O16573));
  NOR2X1 G8958 (.A1(I1504), .A2(W28763), .ZN(W47631));
  NOR2X1 G8959 (.A1(W58), .A2(W313), .ZN(W3333));
  NOR2X1 G8960 (.A1(W267), .A2(I1868), .ZN(W3332));
  NOR2X1 G8961 (.A1(W23763), .A2(W38449), .ZN(O16583));
  NOR2X1 G8962 (.A1(I563), .A2(I1538), .ZN(W3329));
  NOR2X1 G8963 (.A1(I740), .A2(W1962), .ZN(W3328));
  NOR2X1 G8964 (.A1(W11345), .A2(W9048), .ZN(O3777));
  NOR2X1 G8965 (.A1(W29823), .A2(W25750), .ZN(O16586));
  NOR2X1 G8966 (.A1(I1031), .A2(I1473), .ZN(W3353));
  NOR2X1 G8967 (.A1(W20961), .A2(W39319), .ZN(O16557));
  NOR2X1 G8968 (.A1(W35627), .A2(W12095), .ZN(O16558));
  NOR2X1 G8969 (.A1(W4560), .A2(I242), .ZN(O16559));
  NOR2X1 G8970 (.A1(W2294), .A2(I1529), .ZN(W3360));
  NOR2X1 G8971 (.A1(W43017), .A2(W38014), .ZN(O16561));
  NOR2X1 G8972 (.A1(W4244), .A2(W23497), .ZN(W26508));
  NOR2X1 G8973 (.A1(W12439), .A2(W42296), .ZN(W47613));
  NOR2X1 G8974 (.A1(W22071), .A2(W16124), .ZN(O16568));
  NOR2X1 G8975 (.A1(W4444), .A2(W12774), .ZN(O16587));
  NOR2X1 G8976 (.A1(I1220), .A2(W7260), .ZN(W24234));
  NOR2X1 G8977 (.A1(W1366), .A2(W506), .ZN(W3351));
  NOR2X1 G8978 (.A1(W4263), .A2(W7222), .ZN(W26506));
  NOR2X1 G8979 (.A1(W1678), .A2(W2416), .ZN(W3349));
  NOR2X1 G8980 (.A1(W3167), .A2(I796), .ZN(W3348));
  NOR2X1 G8981 (.A1(W2071), .A2(W1038), .ZN(W3347));
  NOR2X1 G8982 (.A1(I66), .A2(W2558), .ZN(W3346));
  NOR2X1 G8983 (.A1(I1510), .A2(W28496), .ZN(O16610));
  NOR2X1 G8984 (.A1(W1508), .A2(I1348), .ZN(W3304));
  NOR2X1 G8985 (.A1(W3267), .A2(W34717), .ZN(O16604));
  NOR2X1 G8986 (.A1(I423), .A2(W298), .ZN(W3302));
  NOR2X1 G8987 (.A1(W835), .A2(I870), .ZN(W3301));
  NOR2X1 G8988 (.A1(I1262), .A2(W3064), .ZN(W3300));
  NOR2X1 G8989 (.A1(W23597), .A2(W14003), .ZN(O3017));
  NOR2X1 G8990 (.A1(W1258), .A2(I1626), .ZN(W3296));
  NOR2X1 G8991 (.A1(W12947), .A2(W2047), .ZN(O3018));
  NOR2X1 G8992 (.A1(W22505), .A2(W11866), .ZN(O16603));
  NOR2X1 G8993 (.A1(W11671), .A2(W6587), .ZN(W26487));
  NOR2X1 G8994 (.A1(I924), .A2(W2441), .ZN(W3290));
  NOR2X1 G8995 (.A1(W2867), .A2(W2268), .ZN(W3289));
  NOR2X1 G8996 (.A1(W7591), .A2(W43030), .ZN(O16615));
  NOR2X1 G8997 (.A1(W2860), .A2(W1965), .ZN(W3287));
  NOR2X1 G8998 (.A1(W32235), .A2(W8721), .ZN(O16616));
  NOR2X1 G8999 (.A1(W532), .A2(W1565), .ZN(W3285));
  NOR2X1 G9000 (.A1(I562), .A2(W23298), .ZN(W24254));
  NOR2X1 G9001 (.A1(W2643), .A2(W1192), .ZN(W3315));
  NOR2X1 G9002 (.A1(I1018), .A2(W21705), .ZN(W26499));
  NOR2X1 G9003 (.A1(W1699), .A2(W2975), .ZN(W3323));
  NOR2X1 G9004 (.A1(W39681), .A2(W10690), .ZN(O16591));
  NOR2X1 G9005 (.A1(W28814), .A2(W21828), .ZN(O16592));
  NOR2X1 G9006 (.A1(W538), .A2(W722), .ZN(W3319));
  NOR2X1 G9007 (.A1(W1682), .A2(W2747), .ZN(W3318));
  NOR2X1 G9008 (.A1(W2509), .A2(W1580), .ZN(W3317));
  NOR2X1 G9009 (.A1(W3339), .A2(W25260), .ZN(O16594));
  NOR2X1 G9010 (.A1(W528), .A2(W19890), .ZN(O3008));
  NOR2X1 G9011 (.A1(W44143), .A2(W5353), .ZN(O16595));
  NOR2X1 G9012 (.A1(W5900), .A2(W23340), .ZN(W24244));
  NOR2X1 G9013 (.A1(W20863), .A2(W13661), .ZN(O16597));
  NOR2X1 G9014 (.A1(W35584), .A2(W41645), .ZN(O16598));
  NOR2X1 G9015 (.A1(W1733), .A2(I433), .ZN(W3310));
  NOR2X1 G9016 (.A1(W13336), .A2(W45504), .ZN(O16600));
  NOR2X1 G9017 (.A1(W2586), .A2(W3122), .ZN(W3308));
  NOR2X1 G9018 (.A1(W14301), .A2(W14964), .ZN(W24216));
  NOR2X1 G9019 (.A1(W10761), .A2(W14584), .ZN(W26534));
  NOR2X1 G9020 (.A1(W124), .A2(W1403), .ZN(W3425));
  NOR2X1 G9021 (.A1(I1302), .A2(I44), .ZN(W3423));
  NOR2X1 G9022 (.A1(W2317), .A2(W431), .ZN(W3422));
  NOR2X1 G9023 (.A1(I1084), .A2(I741), .ZN(W3421));
  NOR2X1 G9024 (.A1(W2590), .A2(W1362), .ZN(W3418));
  NOR2X1 G9025 (.A1(W18093), .A2(W19777), .ZN(O16513));
  NOR2X1 G9026 (.A1(W1790), .A2(W332), .ZN(W3416));
  NOR2X1 G9027 (.A1(W664), .A2(W2335), .ZN(W3427));
  NOR2X1 G9028 (.A1(W1), .A2(W1118), .ZN(W3414));
  NOR2X1 G9029 (.A1(W37744), .A2(I1288), .ZN(W47557));
  NOR2X1 G9030 (.A1(W10829), .A2(W13003), .ZN(O16516));
  NOR2X1 G9031 (.A1(W27955), .A2(W38982), .ZN(W47559));
  NOR2X1 G9032 (.A1(W43110), .A2(W8889), .ZN(W47560));
  NOR2X1 G9033 (.A1(W2567), .A2(I1847), .ZN(W3409));
  NOR2X1 G9034 (.A1(W45699), .A2(W30787), .ZN(O16518));
  NOR2X1 G9035 (.A1(I878), .A2(W3194), .ZN(W3407));
  NOR2X1 G9036 (.A1(W34615), .A2(W33142), .ZN(O16502));
  NOR2X1 G9037 (.A1(W11952), .A2(W9097), .ZN(W47529));
  NOR2X1 G9038 (.A1(W19550), .A2(W5605), .ZN(O2999));
  NOR2X1 G9039 (.A1(W9617), .A2(W226), .ZN(W26538));
  NOR2X1 G9040 (.A1(W44882), .A2(W39382), .ZN(O16494));
  NOR2X1 G9041 (.A1(W1045), .A2(W255), .ZN(W3441));
  NOR2X1 G9042 (.A1(W9330), .A2(W13562), .ZN(O16495));
  NOR2X1 G9043 (.A1(W32263), .A2(W28149), .ZN(O16496));
  NOR2X1 G9044 (.A1(W4867), .A2(W18373), .ZN(O16501));
  NOR2X1 G9045 (.A1(W21697), .A2(W19315), .ZN(O16519));
  NOR2X1 G9046 (.A1(W3329), .A2(I1423), .ZN(W3435));
  NOR2X1 G9047 (.A1(I1919), .A2(W1084), .ZN(W3434));
  NOR2X1 G9048 (.A1(W1799), .A2(I332), .ZN(W3432));
  NOR2X1 G9049 (.A1(W768), .A2(W529), .ZN(W3431));
  NOR2X1 G9050 (.A1(W171), .A2(W2706), .ZN(W3430));
  NOR2X1 G9051 (.A1(W916), .A2(I1302), .ZN(W3429));
  NOR2X1 G9052 (.A1(W16054), .A2(W40171), .ZN(O16505));
  NOR2X1 G9053 (.A1(W1709), .A2(W535), .ZN(W3373));
  NOR2X1 G9054 (.A1(I1108), .A2(I164), .ZN(W3383));
  NOR2X1 G9055 (.A1(I1612), .A2(W24723), .ZN(O16540));
  NOR2X1 G9056 (.A1(W19047), .A2(W21937), .ZN(O3779));
  NOR2X1 G9057 (.A1(I1025), .A2(I1514), .ZN(W3379));
  NOR2X1 G9058 (.A1(W42918), .A2(W33352), .ZN(O16543));
  NOR2X1 G9059 (.A1(W16243), .A2(W7268), .ZN(W24227));
  NOR2X1 G9060 (.A1(W1711), .A2(W28219), .ZN(O16550));
  NOR2X1 G9061 (.A1(I1180), .A2(W2775), .ZN(W3374));
  NOR2X1 G9062 (.A1(W40216), .A2(W37393), .ZN(O16538));
  NOR2X1 G9063 (.A1(W2366), .A2(W388), .ZN(W3372));
  NOR2X1 G9064 (.A1(W10289), .A2(W9059), .ZN(W24229));
  NOR2X1 G9065 (.A1(W18731), .A2(W42805), .ZN(O16554));
  NOR2X1 G9066 (.A1(W1601), .A2(W510), .ZN(W3368));
  NOR2X1 G9067 (.A1(W2414), .A2(W230), .ZN(O34));
  NOR2X1 G9068 (.A1(I1078), .A2(I1970), .ZN(O33));
  NOR2X1 G9069 (.A1(W7400), .A2(W28397), .ZN(O16555));
  NOR2X1 G9070 (.A1(W1824), .A2(W1573), .ZN(W3393));
  NOR2X1 G9071 (.A1(W7101), .A2(W10213), .ZN(O16520));
  NOR2X1 G9072 (.A1(W10331), .A2(W16629), .ZN(O3784));
  NOR2X1 G9073 (.A1(W11062), .A2(W1766), .ZN(W26527));
  NOR2X1 G9074 (.A1(I224), .A2(W22), .ZN(O35));
  NOR2X1 G9075 (.A1(W20340), .A2(W10487), .ZN(O16524));
  NOR2X1 G9076 (.A1(I1675), .A2(W1121), .ZN(W3397));
  NOR2X1 G9077 (.A1(I1056), .A2(W44292), .ZN(O16527));
  NOR2X1 G9078 (.A1(W32374), .A2(W34230), .ZN(O16529));
  NOR2X1 G9079 (.A1(W37710), .A2(W38542), .ZN(O16619));
  NOR2X1 G9080 (.A1(W34583), .A2(W36435), .ZN(O16530));
  NOR2X1 G9081 (.A1(I1703), .A2(W2724), .ZN(W3391));
  NOR2X1 G9082 (.A1(W16205), .A2(W26408), .ZN(O16532));
  NOR2X1 G9083 (.A1(W3108), .A2(I1068), .ZN(W3389));
  NOR2X1 G9084 (.A1(W33528), .A2(W26358), .ZN(O16533));
  NOR2X1 G9085 (.A1(W2639), .A2(W3101), .ZN(W3387));
  NOR2X1 G9086 (.A1(W23292), .A2(W43492), .ZN(O16537));
  NOR2X1 G9087 (.A1(W34694), .A2(I830), .ZN(O16725));
  NOR2X1 G9088 (.A1(W24626), .A2(W15911), .ZN(W26457));
  NOR2X1 G9089 (.A1(I462), .A2(I1177), .ZN(W3185));
  NOR2X1 G9090 (.A1(I1034), .A2(I952), .ZN(W3184));
  NOR2X1 G9091 (.A1(I1048), .A2(I1452), .ZN(W3183));
  NOR2X1 G9092 (.A1(W24099), .A2(W17161), .ZN(W26455));
  NOR2X1 G9093 (.A1(W1690), .A2(W7877), .ZN(W24288));
  NOR2X1 G9094 (.A1(I263), .A2(W2850), .ZN(W3180));
  NOR2X1 G9095 (.A1(W2861), .A2(W10545), .ZN(W24289));
  NOR2X1 G9096 (.A1(I1816), .A2(W38818), .ZN(O16715));
  NOR2X1 G9097 (.A1(W15987), .A2(W32209), .ZN(O16728));
  NOR2X1 G9098 (.A1(W10233), .A2(W11410), .ZN(W24290));
  NOR2X1 G9099 (.A1(I235), .A2(W682), .ZN(W3175));
  NOR2X1 G9100 (.A1(W46852), .A2(W4845), .ZN(O16731));
  NOR2X1 G9101 (.A1(W23895), .A2(W4974), .ZN(W26454));
  NOR2X1 G9102 (.A1(W7014), .A2(W5002), .ZN(W24292));
  NOR2X1 G9103 (.A1(W1392), .A2(W3066), .ZN(W3170));
  NOR2X1 G9104 (.A1(I988), .A2(I431), .ZN(W3169));
  NOR2X1 G9105 (.A1(W11741), .A2(W4218), .ZN(W24284));
  NOR2X1 G9106 (.A1(W25416), .A2(W14582), .ZN(W26461));
  NOR2X1 G9107 (.A1(W25899), .A2(W4734), .ZN(O16702));
  NOR2X1 G9108 (.A1(W223), .A2(W40016), .ZN(O16704));
  NOR2X1 G9109 (.A1(W39574), .A2(W37575), .ZN(W47763));
  NOR2X1 G9110 (.A1(W35988), .A2(W35688), .ZN(O16705));
  NOR2X1 G9111 (.A1(W45845), .A2(W3847), .ZN(O16706));
  NOR2X1 G9112 (.A1(I1177), .A2(I776), .ZN(W3197));
  NOR2X1 G9113 (.A1(W6210), .A2(W27529), .ZN(O16708));
  NOR2X1 G9114 (.A1(W14387), .A2(W30291), .ZN(O16741));
  NOR2X1 G9115 (.A1(W19696), .A2(W27686), .ZN(O16709));
  NOR2X1 G9116 (.A1(W12905), .A2(W41371), .ZN(O16710));
  NOR2X1 G9117 (.A1(W38893), .A2(W3061), .ZN(O16712));
  NOR2X1 G9118 (.A1(W46606), .A2(W16082), .ZN(O16713));
  NOR2X1 G9119 (.A1(W938), .A2(I42), .ZN(W3190));
  NOR2X1 G9120 (.A1(W11978), .A2(I1041), .ZN(O3761));
  NOR2X1 G9121 (.A1(W7605), .A2(W14157), .ZN(W47775));
  NOR2X1 G9122 (.A1(I1988), .A2(W1125), .ZN(W3138));
  NOR2X1 G9123 (.A1(W1186), .A2(W1053), .ZN(W3147));
  NOR2X1 G9124 (.A1(W3399), .A2(W12070), .ZN(W24302));
  NOR2X1 G9125 (.A1(W2559), .A2(I1752), .ZN(W3145));
  NOR2X1 G9126 (.A1(W2495), .A2(I130), .ZN(W3144));
  NOR2X1 G9127 (.A1(W1970), .A2(I939), .ZN(W3143));
  NOR2X1 G9128 (.A1(W38822), .A2(W15547), .ZN(O16764));
  NOR2X1 G9129 (.A1(W22568), .A2(W20035), .ZN(O3039));
  NOR2X1 G9130 (.A1(I926), .A2(W2131), .ZN(W3139));
  NOR2X1 G9131 (.A1(W13569), .A2(W27996), .ZN(O16761));
  NOR2X1 G9132 (.A1(W7593), .A2(W25308), .ZN(O16771));
  NOR2X1 G9133 (.A1(I1364), .A2(W43459), .ZN(O16773));
  NOR2X1 G9134 (.A1(W2249), .A2(W39), .ZN(W3135));
  NOR2X1 G9135 (.A1(I376), .A2(W1346), .ZN(W3134));
  NOR2X1 G9136 (.A1(I708), .A2(W2164), .ZN(W3133));
  NOR2X1 G9137 (.A1(W14913), .A2(W17806), .ZN(W26438));
  NOR2X1 G9138 (.A1(I923), .A2(I421), .ZN(W3131));
  NOR2X1 G9139 (.A1(W27081), .A2(W24774), .ZN(O16754));
  NOR2X1 G9140 (.A1(W1219), .A2(I1501), .ZN(W3167));
  NOR2X1 G9141 (.A1(W12100), .A2(W18892), .ZN(W26451));
  NOR2X1 G9142 (.A1(I1938), .A2(W20052), .ZN(O16743));
  NOR2X1 G9143 (.A1(W2761), .A2(W18119), .ZN(W26450));
  NOR2X1 G9144 (.A1(W3245), .A2(W26980), .ZN(O16746));
  NOR2X1 G9145 (.A1(W32047), .A2(W7303), .ZN(W47815));
  NOR2X1 G9146 (.A1(W2100), .A2(W3139), .ZN(W3159));
  NOR2X1 G9147 (.A1(I777), .A2(W3157), .ZN(W3158));
  NOR2X1 G9148 (.A1(W1670), .A2(W3166), .ZN(W3204));
  NOR2X1 G9149 (.A1(W12895), .A2(W23579), .ZN(O3758));
  NOR2X1 G9150 (.A1(W27055), .A2(W11867), .ZN(O16758));
  NOR2X1 G9151 (.A1(W12582), .A2(W13691), .ZN(W47822));
  NOR2X1 G9152 (.A1(I958), .A2(I1976), .ZN(W3152));
  NOR2X1 G9153 (.A1(W10061), .A2(W586), .ZN(W24300));
  NOR2X1 G9154 (.A1(I818), .A2(W1860), .ZN(W3150));
  NOR2X1 G9155 (.A1(W14204), .A2(W8075), .ZN(O3037));
  NOR2X1 G9156 (.A1(W10300), .A2(W36295), .ZN(O16649));
  NOR2X1 G9157 (.A1(W36456), .A2(W31647), .ZN(O16637));
  NOR2X1 G9158 (.A1(W4542), .A2(W13373), .ZN(O3021));
  NOR2X1 G9159 (.A1(I280), .A2(W13304), .ZN(O16639));
  NOR2X1 G9160 (.A1(W2660), .A2(W18809), .ZN(O3022));
  NOR2X1 G9161 (.A1(W69), .A2(W43142), .ZN(O16643));
  NOR2X1 G9162 (.A1(W1440), .A2(W2455), .ZN(W3256));
  NOR2X1 G9163 (.A1(W8844), .A2(W23238), .ZN(O3023));
  NOR2X1 G9164 (.A1(W24790), .A2(W45728), .ZN(O16648));
  NOR2X1 G9165 (.A1(W363), .A2(W3032), .ZN(W3263));
  NOR2X1 G9166 (.A1(I686), .A2(W972), .ZN(W3251));
  NOR2X1 G9167 (.A1(W15035), .A2(W3385), .ZN(O16650));
  NOR2X1 G9168 (.A1(W1531), .A2(I121), .ZN(W3249));
  NOR2X1 G9169 (.A1(W3105), .A2(W1024), .ZN(W3248));
  NOR2X1 G9170 (.A1(W2269), .A2(I1488), .ZN(W3247));
  NOR2X1 G9171 (.A1(W2100), .A2(W2223), .ZN(W3246));
  NOR2X1 G9172 (.A1(W4746), .A2(W12844), .ZN(O16651));
  NOR2X1 G9173 (.A1(W19881), .A2(W25942), .ZN(O16653));
  NOR2X1 G9174 (.A1(I907), .A2(W43035), .ZN(O16633));
  NOR2X1 G9175 (.A1(W28965), .A2(W19177), .ZN(O16620));
  NOR2X1 G9176 (.A1(W23317), .A2(W18910), .ZN(W24256));
  NOR2X1 G9177 (.A1(W34610), .A2(W7348), .ZN(O16627));
  NOR2X1 G9178 (.A1(I809), .A2(W1256), .ZN(W3278));
  NOR2X1 G9179 (.A1(W11726), .A2(W20600), .ZN(W24257));
  NOR2X1 G9180 (.A1(W29101), .A2(W2645), .ZN(O16630));
  NOR2X1 G9181 (.A1(W17540), .A2(W8139), .ZN(W26480));
  NOR2X1 G9182 (.A1(W30665), .A2(W39674), .ZN(O16632));
  NOR2X1 G9183 (.A1(W34687), .A2(W28194), .ZN(O16654));
  NOR2X1 G9184 (.A1(W2424), .A2(W2559), .ZN(W3271));
  NOR2X1 G9185 (.A1(W137), .A2(W1519), .ZN(W3270));
  NOR2X1 G9186 (.A1(W3347), .A2(W16182), .ZN(O3769));
  NOR2X1 G9187 (.A1(W2552), .A2(I464), .ZN(W3268));
  NOR2X1 G9188 (.A1(W2639), .A2(I284), .ZN(W3267));
  NOR2X1 G9189 (.A1(W910), .A2(W2850), .ZN(W3266));
  NOR2X1 G9190 (.A1(W18589), .A2(W11945), .ZN(W24262));
  NOR2X1 G9191 (.A1(I282), .A2(W2032), .ZN(W3213));
  NOR2X1 G9192 (.A1(W8755), .A2(W7432), .ZN(W24276));
  NOR2X1 G9193 (.A1(W376), .A2(W8254), .ZN(W24277));
  NOR2X1 G9194 (.A1(I1802), .A2(W43), .ZN(W3219));
  NOR2X1 G9195 (.A1(W2676), .A2(W2402), .ZN(W3218));
  NOR2X1 G9196 (.A1(I1235), .A2(I916), .ZN(W3217));
  NOR2X1 G9197 (.A1(W1251), .A2(W36160), .ZN(O16678));
  NOR2X1 G9198 (.A1(W1938), .A2(W41293), .ZN(O16680));
  NOR2X1 G9199 (.A1(W4419), .A2(W9194), .ZN(O3030));
  NOR2X1 G9200 (.A1(W11827), .A2(W20894), .ZN(O3029));
  NOR2X1 G9201 (.A1(W7992), .A2(W14123), .ZN(W24279));
  NOR2X1 G9202 (.A1(W27695), .A2(W17391), .ZN(O16686));
  NOR2X1 G9203 (.A1(W3080), .A2(W2344), .ZN(W3210));
  NOR2X1 G9204 (.A1(W20852), .A2(W11913), .ZN(O3031));
  NOR2X1 G9205 (.A1(W2798), .A2(W4862), .ZN(W24281));
  NOR2X1 G9206 (.A1(W20752), .A2(W9351), .ZN(O16692));
  NOR2X1 G9207 (.A1(W30908), .A2(W18818), .ZN(W47751));
  NOR2X1 G9208 (.A1(W2214), .A2(W33991), .ZN(O16667));
  NOR2X1 G9209 (.A1(W23284), .A2(W6289), .ZN(W26468));
  NOR2X1 G9210 (.A1(W26325), .A2(W7015), .ZN(W26467));
  NOR2X1 G9211 (.A1(W17992), .A2(W23097), .ZN(O3025));
  NOR2X1 G9212 (.A1(W35727), .A2(W17296), .ZN(O16662));
  NOR2X1 G9213 (.A1(I520), .A2(W1375), .ZN(W3237));
  NOR2X1 G9214 (.A1(W203), .A2(I521), .ZN(W3236));
  NOR2X1 G9215 (.A1(W32804), .A2(W4718), .ZN(O16665));
  NOR2X1 G9216 (.A1(W39507), .A2(W41666), .ZN(O16666));
  NOR2X1 G9217 (.A1(W21658), .A2(W4216), .ZN(O16491));
  NOR2X1 G9218 (.A1(W1828), .A2(W1877), .ZN(W3231));
  NOR2X1 G9219 (.A1(W763), .A2(I1985), .ZN(W3228));
  NOR2X1 G9220 (.A1(W2371), .A2(W1584), .ZN(W3227));
  NOR2X1 G9221 (.A1(W2068), .A2(W337), .ZN(W3226));
  NOR2X1 G9222 (.A1(I566), .A2(I827), .ZN(W3225));
  NOR2X1 G9223 (.A1(W19949), .A2(W7459), .ZN(O16672));
  NOR2X1 G9224 (.A1(W956), .A2(W2012), .ZN(W3223));
  NOR2X1 G9225 (.A1(I938), .A2(W2148), .ZN(W3647));
  NOR2X1 G9226 (.A1(W9028), .A2(W2599), .ZN(O16304));
  NOR2X1 G9227 (.A1(W1429), .A2(W232), .ZN(W3654));
  NOR2X1 G9228 (.A1(W2323), .A2(W852), .ZN(W3653));
  NOR2X1 G9229 (.A1(W1562), .A2(W2380), .ZN(W3652));
  NOR2X1 G9230 (.A1(I862), .A2(I1859), .ZN(W3651));
  NOR2X1 G9231 (.A1(W9513), .A2(W10233), .ZN(O16308));
  NOR2X1 G9232 (.A1(W19481), .A2(W1140), .ZN(W26596));
  NOR2X1 G9233 (.A1(W1412), .A2(W6759), .ZN(O2983));
  NOR2X1 G9234 (.A1(W5210), .A2(W5277), .ZN(W26597));
  NOR2X1 G9235 (.A1(W1003), .A2(I608), .ZN(W3646));
  NOR2X1 G9236 (.A1(W11269), .A2(W15062), .ZN(O2984));
  NOR2X1 G9237 (.A1(W919), .A2(I999), .ZN(W3644));
  NOR2X1 G9238 (.A1(W3428), .A2(I1577), .ZN(W3643));
  NOR2X1 G9239 (.A1(W10307), .A2(W23313), .ZN(O2985));
  NOR2X1 G9240 (.A1(W42145), .A2(W10295), .ZN(O16318));
  NOR2X1 G9241 (.A1(W63), .A2(W4), .ZN(W3640));
  NOR2X1 G9242 (.A1(I1145), .A2(I1234), .ZN(W3639));
  NOR2X1 G9243 (.A1(W12337), .A2(W23003), .ZN(O16299));
  NOR2X1 G9244 (.A1(W11509), .A2(W36215), .ZN(O16290));
  NOR2X1 G9245 (.A1(W6561), .A2(W23674), .ZN(O16291));
  NOR2X1 G9246 (.A1(W1810), .A2(I839), .ZN(W3671));
  NOR2X1 G9247 (.A1(W5338), .A2(W6765), .ZN(W24142));
  NOR2X1 G9248 (.A1(W17502), .A2(W5599), .ZN(O16293));
  NOR2X1 G9249 (.A1(W6332), .A2(W11830), .ZN(O2981));
  NOR2X1 G9250 (.A1(W16055), .A2(W24643), .ZN(O16296));
  NOR2X1 G9251 (.A1(W33300), .A2(W24441), .ZN(O16297));
  NOR2X1 G9252 (.A1(W3218), .A2(I505), .ZN(W3638));
  NOR2X1 G9253 (.A1(W46974), .A2(W35958), .ZN(O16300));
  NOR2X1 G9254 (.A1(I656), .A2(W2145), .ZN(W3663));
  NOR2X1 G9255 (.A1(W2627), .A2(I1372), .ZN(W3661));
  NOR2X1 G9256 (.A1(I518), .A2(W2532), .ZN(W3660));
  NOR2X1 G9257 (.A1(I1654), .A2(W1757), .ZN(W3659));
  NOR2X1 G9258 (.A1(W6867), .A2(W42594), .ZN(W47319));
  NOR2X1 G9259 (.A1(W17224), .A2(W42783), .ZN(O16302));
  NOR2X1 G9260 (.A1(W15638), .A2(W15490), .ZN(O16344));
  NOR2X1 G9261 (.A1(W27712), .A2(W10627), .ZN(O16336));
  NOR2X1 G9262 (.A1(W16091), .A2(W23996), .ZN(O2986));
  NOR2X1 G9263 (.A1(W2928), .A2(W2887), .ZN(W3617));
  NOR2X1 G9264 (.A1(W1964), .A2(I813), .ZN(W3616));
  NOR2X1 G9265 (.A1(W202), .A2(I1252), .ZN(W3615));
  NOR2X1 G9266 (.A1(W2317), .A2(W14669), .ZN(O3804));
  NOR2X1 G9267 (.A1(W3226), .A2(W15900), .ZN(O16341));
  NOR2X1 G9268 (.A1(W11329), .A2(W3468), .ZN(W24154));
  NOR2X1 G9269 (.A1(W38199), .A2(W45237), .ZN(O16335));
  NOR2X1 G9270 (.A1(W279), .A2(W3112), .ZN(W3610));
  NOR2X1 G9271 (.A1(W3191), .A2(W12056), .ZN(O16346));
  NOR2X1 G9272 (.A1(W2344), .A2(I316), .ZN(W3608));
  NOR2X1 G9273 (.A1(W19594), .A2(I462), .ZN(W26592));
  NOR2X1 G9274 (.A1(W1437), .A2(W1575), .ZN(W3605));
  NOR2X1 G9275 (.A1(W7777), .A2(W18499), .ZN(W47372));
  NOR2X1 G9276 (.A1(I198), .A2(W8808), .ZN(W24158));
  NOR2X1 G9277 (.A1(W10264), .A2(W8870), .ZN(O16325));
  NOR2X1 G9278 (.A1(W6420), .A2(W13789), .ZN(W47338));
  NOR2X1 G9279 (.A1(W39089), .A2(W21401), .ZN(O16323));
  NOR2X1 G9280 (.A1(I1419), .A2(W2482), .ZN(W3635));
  NOR2X1 G9281 (.A1(W1970), .A2(W3416), .ZN(W3634));
  NOR2X1 G9282 (.A1(I1346), .A2(W1676), .ZN(W3633));
  NOR2X1 G9283 (.A1(W1687), .A2(W1353), .ZN(W3632));
  NOR2X1 G9284 (.A1(W13494), .A2(W18721), .ZN(O16324));
  NOR2X1 G9285 (.A1(W539), .A2(I1881), .ZN(W3630));
  NOR2X1 G9286 (.A1(W20564), .A2(W23082), .ZN(W24141));
  NOR2X1 G9287 (.A1(W11404), .A2(W22300), .ZN(O16326));
  NOR2X1 G9288 (.A1(W19846), .A2(W8997), .ZN(W24150));
  NOR2X1 G9289 (.A1(W27717), .A2(W35585), .ZN(O16330));
  NOR2X1 G9290 (.A1(W2819), .A2(I455), .ZN(W3625));
  NOR2X1 G9291 (.A1(W21911), .A2(W20256), .ZN(O16331));
  NOR2X1 G9292 (.A1(I478), .A2(W1091), .ZN(W3623));
  NOR2X1 G9293 (.A1(I413), .A2(I853), .ZN(W3621));
  NOR2X1 G9294 (.A1(W5812), .A2(W6310), .ZN(O16238));
  NOR2X1 G9295 (.A1(W10745), .A2(W1799), .ZN(O3810));
  NOR2X1 G9296 (.A1(W5542), .A2(W44071), .ZN(O16231));
  NOR2X1 G9297 (.A1(W8237), .A2(W15685), .ZN(W47239));
  NOR2X1 G9298 (.A1(W14257), .A2(W5471), .ZN(O16233));
  NOR2X1 G9299 (.A1(W18407), .A2(W21157), .ZN(O16234));
  NOR2X1 G9300 (.A1(I1786), .A2(W2994), .ZN(W3731));
  NOR2X1 G9301 (.A1(W21443), .A2(W12109), .ZN(W24119));
  NOR2X1 G9302 (.A1(W11400), .A2(W7721), .ZN(W24120));
  NOR2X1 G9303 (.A1(W6277), .A2(W10469), .ZN(W24116));
  NOR2X1 G9304 (.A1(W665), .A2(W2446), .ZN(W3727));
  NOR2X1 G9305 (.A1(W32028), .A2(W16339), .ZN(O16242));
  NOR2X1 G9306 (.A1(W2035), .A2(W3323), .ZN(W3725));
  NOR2X1 G9307 (.A1(W3066), .A2(W2000), .ZN(W3724));
  NOR2X1 G9308 (.A1(W2357), .A2(I1217), .ZN(W26618));
  NOR2X1 G9309 (.A1(I1331), .A2(I1114), .ZN(W3721));
  NOR2X1 G9310 (.A1(W14135), .A2(W19306), .ZN(W24123));
  NOR2X1 G9311 (.A1(W22283), .A2(W14283), .ZN(W24124));
  NOR2X1 G9312 (.A1(W13091), .A2(W5489), .ZN(W26629));
  NOR2X1 G9313 (.A1(W54), .A2(W3193), .ZN(W3756));
  NOR2X1 G9314 (.A1(W36133), .A2(W15628), .ZN(O16212));
  NOR2X1 G9315 (.A1(W15078), .A2(W28780), .ZN(O16214));
  NOR2X1 G9316 (.A1(W3471), .A2(W1540), .ZN(O3813));
  NOR2X1 G9317 (.A1(I1510), .A2(W2545), .ZN(W3752));
  NOR2X1 G9318 (.A1(W12925), .A2(W35807), .ZN(O16216));
  NOR2X1 G9319 (.A1(W5923), .A2(W38054), .ZN(O16219));
  NOR2X1 G9320 (.A1(W7047), .A2(W44348), .ZN(O16220));
  NOR2X1 G9321 (.A1(W5174), .A2(W24117), .ZN(O16249));
  NOR2X1 G9322 (.A1(I912), .A2(W13995), .ZN(W24114));
  NOR2X1 G9323 (.A1(W35277), .A2(W3978), .ZN(O16223));
  NOR2X1 G9324 (.A1(W12490), .A2(W41469), .ZN(O16224));
  NOR2X1 G9325 (.A1(W1646), .A2(W3158), .ZN(W3743));
  NOR2X1 G9326 (.A1(I1565), .A2(I1003), .ZN(W3742));
  NOR2X1 G9327 (.A1(W148), .A2(W537), .ZN(W3741));
  NOR2X1 G9328 (.A1(W31259), .A2(W11209), .ZN(O16225));
  NOR2X1 G9329 (.A1(W43942), .A2(W43947), .ZN(O16274));
  NOR2X1 G9330 (.A1(W9822), .A2(W14493), .ZN(O16266));
  NOR2X1 G9331 (.A1(W2915), .A2(I21), .ZN(W3696));
  NOR2X1 G9332 (.A1(W3039), .A2(W13580), .ZN(W26609));
  NOR2X1 G9333 (.A1(W26484), .A2(W21946), .ZN(W47278));
  NOR2X1 G9334 (.A1(W5529), .A2(W21049), .ZN(W24132));
  NOR2X1 G9335 (.A1(W27070), .A2(W20089), .ZN(O16272));
  NOR2X1 G9336 (.A1(W37917), .A2(W41647), .ZN(W47285));
  NOR2X1 G9337 (.A1(W250), .A2(W3562), .ZN(W3688));
  NOR2X1 G9338 (.A1(W12821), .A2(W16055), .ZN(W26610));
  NOR2X1 G9339 (.A1(W2378), .A2(I1184), .ZN(W3686));
  NOR2X1 G9340 (.A1(W11784), .A2(W37797), .ZN(O16275));
  NOR2X1 G9341 (.A1(I782), .A2(I1913), .ZN(W3684));
  NOR2X1 G9342 (.A1(W28804), .A2(W30455), .ZN(O16277));
  NOR2X1 G9343 (.A1(W5830), .A2(W47041), .ZN(O16279));
  NOR2X1 G9344 (.A1(W1743), .A2(W20219), .ZN(O3806));
  NOR2X1 G9345 (.A1(W36757), .A2(W33644), .ZN(W47299));
  NOR2X1 G9346 (.A1(I708), .A2(W2361), .ZN(W3708));
  NOR2X1 G9347 (.A1(W1352), .A2(I169), .ZN(W3717));
  NOR2X1 G9348 (.A1(W1615), .A2(W2521), .ZN(W3716));
  NOR2X1 G9349 (.A1(I1834), .A2(I995), .ZN(W3715));
  NOR2X1 G9350 (.A1(W46242), .A2(W43981), .ZN(O16251));
  NOR2X1 G9351 (.A1(W187), .A2(W44), .ZN(W3712));
  NOR2X1 G9352 (.A1(W13005), .A2(W520), .ZN(W24126));
  NOR2X1 G9353 (.A1(W1026), .A2(W180), .ZN(W3710));
  NOR2X1 G9354 (.A1(I1714), .A2(W1064), .ZN(W3709));
  NOR2X1 G9355 (.A1(W25797), .A2(W32220), .ZN(O16353));
  NOR2X1 G9356 (.A1(W506), .A2(W3219), .ZN(W3707));
  NOR2X1 G9357 (.A1(W4325), .A2(W17618), .ZN(W47266));
  NOR2X1 G9358 (.A1(W3293), .A2(W3062), .ZN(W3704));
  NOR2X1 G9359 (.A1(W4053), .A2(W7492), .ZN(O16261));
  NOR2X1 G9360 (.A1(W10455), .A2(W20913), .ZN(W26611));
  NOR2X1 G9361 (.A1(I1712), .A2(W3598), .ZN(W3700));
  NOR2X1 G9362 (.A1(W20135), .A2(W44406), .ZN(O16264));
  NOR2X1 G9363 (.A1(W118), .A2(I912), .ZN(W3492));
  NOR2X1 G9364 (.A1(W14764), .A2(W8706), .ZN(W26558));
  NOR2X1 G9365 (.A1(W13119), .A2(W10406), .ZN(W24193));
  NOR2X1 G9366 (.A1(W3186), .A2(W19133), .ZN(W24194));
  NOR2X1 G9367 (.A1(W17494), .A2(W17873), .ZN(O2998));
  NOR2X1 G9368 (.A1(W1319), .A2(W1483), .ZN(W3496));
  NOR2X1 G9369 (.A1(W38973), .A2(W271), .ZN(O16448));
  NOR2X1 G9370 (.A1(W12073), .A2(W12775), .ZN(W24196));
  NOR2X1 G9371 (.A1(W170), .A2(I1938), .ZN(W3493));
  NOR2X1 G9372 (.A1(W12241), .A2(W8779), .ZN(W24191));
  NOR2X1 G9373 (.A1(W25), .A2(W3033), .ZN(W3491));
  NOR2X1 G9374 (.A1(W3166), .A2(W1659), .ZN(W3490));
  NOR2X1 G9375 (.A1(W33407), .A2(W9665), .ZN(O16452));
  NOR2X1 G9376 (.A1(I777), .A2(I668), .ZN(W3488));
  NOR2X1 G9377 (.A1(W8911), .A2(W1998), .ZN(W24197));
  NOR2X1 G9378 (.A1(W3452), .A2(W3144), .ZN(W3486));
  NOR2X1 G9379 (.A1(W1223), .A2(W2566), .ZN(W3485));
  NOR2X1 G9380 (.A1(W14244), .A2(W13496), .ZN(W24198));
  NOR2X1 G9381 (.A1(W8772), .A2(W29923), .ZN(O16427));
  NOR2X1 G9382 (.A1(W20968), .A2(W19917), .ZN(O16420));
  NOR2X1 G9383 (.A1(W5920), .A2(W36827), .ZN(O16421));
  NOR2X1 G9384 (.A1(W10178), .A2(W12484), .ZN(W26563));
  NOR2X1 G9385 (.A1(W3509), .A2(W16855), .ZN(O2994));
  NOR2X1 G9386 (.A1(I710), .A2(I1754), .ZN(W3515));
  NOR2X1 G9387 (.A1(W2051), .A2(W18325), .ZN(O2995));
  NOR2X1 G9388 (.A1(W1702), .A2(I1943), .ZN(W3513));
  NOR2X1 G9389 (.A1(W8958), .A2(W21655), .ZN(O16426));
  NOR2X1 G9390 (.A1(I233), .A2(W2383), .ZN(W3483));
  NOR2X1 G9391 (.A1(W11028), .A2(W19673), .ZN(W24186));
  NOR2X1 G9392 (.A1(W2287), .A2(W20096), .ZN(W24187));
  NOR2X1 G9393 (.A1(W45639), .A2(W9042), .ZN(O16431));
  NOR2X1 G9394 (.A1(W44766), .A2(W39098), .ZN(O16433));
  NOR2X1 G9395 (.A1(W1108), .A2(W2958), .ZN(W3505));
  NOR2X1 G9396 (.A1(W31819), .A2(W38622), .ZN(O16437));
  NOR2X1 G9397 (.A1(W11511), .A2(W7711), .ZN(W24190));
  NOR2X1 G9398 (.A1(W19918), .A2(W29299), .ZN(O16482));
  NOR2X1 G9399 (.A1(W3185), .A2(W3453), .ZN(W3463));
  NOR2X1 G9400 (.A1(W30261), .A2(W38770), .ZN(O16479));
  NOR2X1 G9401 (.A1(W7392), .A2(W16157), .ZN(W24205));
  NOR2X1 G9402 (.A1(W38148), .A2(W27484), .ZN(O16480));
  NOR2X1 G9403 (.A1(I1445), .A2(W2022), .ZN(W3459));
  NOR2X1 G9404 (.A1(W44976), .A2(W27803), .ZN(W47516));
  NOR2X1 G9405 (.A1(W903), .A2(W30617), .ZN(O16481));
  NOR2X1 G9406 (.A1(W825), .A2(I32), .ZN(W3456));
  NOR2X1 G9407 (.A1(W12710), .A2(W2296), .ZN(O16477));
  NOR2X1 G9408 (.A1(W19949), .A2(W40608), .ZN(O16483));
  NOR2X1 G9409 (.A1(W3381), .A2(W32450), .ZN(O16484));
  NOR2X1 G9410 (.A1(W214), .A2(W5248), .ZN(O16486));
  NOR2X1 G9411 (.A1(W1120), .A2(W1610), .ZN(W3450));
  NOR2X1 G9412 (.A1(W5342), .A2(W6186), .ZN(W26542));
  NOR2X1 G9413 (.A1(W100), .A2(W472), .ZN(W3448));
  NOR2X1 G9414 (.A1(W34753), .A2(W12434), .ZN(O16490));
  NOR2X1 G9415 (.A1(W3471), .A2(W2383), .ZN(W3472));
  NOR2X1 G9416 (.A1(W35877), .A2(W549), .ZN(O16459));
  NOR2X1 G9417 (.A1(W1692), .A2(W1741), .ZN(W3481));
  NOR2X1 G9418 (.A1(W3704), .A2(W17904), .ZN(W26556));
  NOR2X1 G9419 (.A1(W8031), .A2(W5353), .ZN(O16465));
  NOR2X1 G9420 (.A1(W8927), .A2(I1497), .ZN(O16466));
  NOR2X1 G9421 (.A1(W3454), .A2(W43117), .ZN(O16467));
  NOR2X1 G9422 (.A1(W1163), .A2(W259), .ZN(W3476));
  NOR2X1 G9423 (.A1(W1763), .A2(W474), .ZN(W26555));
  NOR2X1 G9424 (.A1(I1689), .A2(W19601), .ZN(W24182));
  NOR2X1 G9425 (.A1(W46915), .A2(W5086), .ZN(O16471));
  NOR2X1 G9426 (.A1(W15270), .A2(W2247), .ZN(O16473));
  NOR2X1 G9427 (.A1(W4605), .A2(W8215), .ZN(O3792));
  NOR2X1 G9428 (.A1(W16037), .A2(W1143), .ZN(O16475));
  NOR2X1 G9429 (.A1(W1147), .A2(W19998), .ZN(W26545));
  NOR2X1 G9430 (.A1(W3152), .A2(I1773), .ZN(W3466));
  NOR2X1 G9431 (.A1(W158), .A2(W893), .ZN(W3465));
  NOR2X1 G9432 (.A1(W38600), .A2(W6344), .ZN(O16382));
  NOR2X1 G9433 (.A1(W1992), .A2(W2046), .ZN(W3581));
  NOR2X1 G9434 (.A1(W46648), .A2(W24926), .ZN(O16370));
  NOR2X1 G9435 (.A1(W580), .A2(W2248), .ZN(W3578));
  NOR2X1 G9436 (.A1(W1554), .A2(W227), .ZN(W3576));
  NOR2X1 G9437 (.A1(I1671), .A2(W3396), .ZN(W3575));
  NOR2X1 G9438 (.A1(W3432), .A2(W1759), .ZN(W3574));
  NOR2X1 G9439 (.A1(W8187), .A2(W12848), .ZN(W26579));
  NOR2X1 G9440 (.A1(W11700), .A2(W41722), .ZN(O16379));
  NOR2X1 G9441 (.A1(I1375), .A2(W1552), .ZN(W3582));
  NOR2X1 G9442 (.A1(I684), .A2(I1146), .ZN(W3569));
  NOR2X1 G9443 (.A1(I521), .A2(W378), .ZN(W3568));
  NOR2X1 G9444 (.A1(W19998), .A2(W18669), .ZN(W26575));
  NOR2X1 G9445 (.A1(W36397), .A2(W45595), .ZN(O16384));
  NOR2X1 G9446 (.A1(W1469), .A2(W2396), .ZN(W3565));
  NOR2X1 G9447 (.A1(W13278), .A2(W16613), .ZN(O2989));
  NOR2X1 G9448 (.A1(W15291), .A2(W8173), .ZN(W24172));
  NOR2X1 G9449 (.A1(W24531), .A2(W7849), .ZN(O16394));
  NOR2X1 G9450 (.A1(W13020), .A2(W46074), .ZN(W47386));
  NOR2X1 G9451 (.A1(I446), .A2(I289), .ZN(W3600));
  NOR2X1 G9452 (.A1(W5793), .A2(I1760), .ZN(W26588));
  NOR2X1 G9453 (.A1(W7679), .A2(W17167), .ZN(W26585));
  NOR2X1 G9454 (.A1(W23483), .A2(W45999), .ZN(O16355));
  NOR2X1 G9455 (.A1(W1352), .A2(W96), .ZN(W3596));
  NOR2X1 G9456 (.A1(W27232), .A2(W15476), .ZN(O16356));
  NOR2X1 G9457 (.A1(W20365), .A2(W45732), .ZN(O16360));
  NOR2X1 G9458 (.A1(I791), .A2(W1738), .ZN(W3592));
  NOR2X1 G9459 (.A1(W2269), .A2(I1254), .ZN(W3558));
  NOR2X1 G9460 (.A1(W2652), .A2(W2245), .ZN(O40));
  NOR2X1 G9461 (.A1(W2310), .A2(W2228), .ZN(W3589));
  NOR2X1 G9462 (.A1(I748), .A2(W3420), .ZN(W3588));
  NOR2X1 G9463 (.A1(W46753), .A2(W45161), .ZN(O16361));
  NOR2X1 G9464 (.A1(W15568), .A2(W13661), .ZN(W26583));
  NOR2X1 G9465 (.A1(W2225), .A2(W2938), .ZN(W3585));
  NOR2X1 G9466 (.A1(W19163), .A2(I1754), .ZN(O16367));
  NOR2X1 G9467 (.A1(W18402), .A2(W15559), .ZN(W24180));
  NOR2X1 G9468 (.A1(W9047), .A2(W6954), .ZN(O16406));
  NOR2X1 G9469 (.A1(W24776), .A2(W10129), .ZN(W26568));
  NOR2X1 G9470 (.A1(W22244), .A2(W12119), .ZN(O16408));
  NOR2X1 G9471 (.A1(W2666), .A2(I168), .ZN(W3536));
  NOR2X1 G9472 (.A1(W6823), .A2(W31642), .ZN(O16409));
  NOR2X1 G9473 (.A1(W20161), .A2(W15222), .ZN(O16410));
  NOR2X1 G9474 (.A1(W1399), .A2(W355), .ZN(W3532));
  NOR2X1 G9475 (.A1(W3222), .A2(W2619), .ZN(W3530));
  NOR2X1 G9476 (.A1(W15894), .A2(W9011), .ZN(O16405));
  NOR2X1 G9477 (.A1(W24791), .A2(W9941), .ZN(O16415));
  NOR2X1 G9478 (.A1(W47117), .A2(W30582), .ZN(O16417));
  NOR2X1 G9479 (.A1(W761), .A2(W1136), .ZN(W3525));
  NOR2X1 G9480 (.A1(I285), .A2(W18488), .ZN(O16418));
  NOR2X1 G9481 (.A1(W21985), .A2(W20375), .ZN(W47448));
  NOR2X1 G9482 (.A1(W982), .A2(W2030), .ZN(W3522));
  NOR2X1 G9483 (.A1(W2882), .A2(W1353), .ZN(W3521));
  NOR2X1 G9484 (.A1(W21349), .A2(W43672), .ZN(O16400));
  NOR2X1 G9485 (.A1(W2189), .A2(W2117), .ZN(W3556));
  NOR2X1 G9486 (.A1(W24299), .A2(W15725), .ZN(O16396));
  NOR2X1 G9487 (.A1(W26666), .A2(W47010), .ZN(O16397));
  NOR2X1 G9488 (.A1(W8713), .A2(W9728), .ZN(W24175));
  NOR2X1 G9489 (.A1(W1648), .A2(W2119), .ZN(W3552));
  NOR2X1 G9490 (.A1(W3346), .A2(I1502), .ZN(W24176));
  NOR2X1 G9491 (.A1(W1812), .A2(W3503), .ZN(W3550));
  NOR2X1 G9492 (.A1(W293), .A2(W2151), .ZN(W3549));
  NOR2X1 G9493 (.A1(W10555), .A2(W12543), .ZN(O16775));
  NOR2X1 G9494 (.A1(W1425), .A2(W2682), .ZN(W3547));
  NOR2X1 G9495 (.A1(W47), .A2(W778), .ZN(W3546));
  NOR2X1 G9496 (.A1(W28358), .A2(W19348), .ZN(O16401));
  NOR2X1 G9497 (.A1(I100), .A2(W3483), .ZN(W3544));
  NOR2X1 G9498 (.A1(W25584), .A2(W17030), .ZN(O16402));
  NOR2X1 G9499 (.A1(W39644), .A2(W4311), .ZN(O16404));
  NOR2X1 G9500 (.A1(W2444), .A2(I991), .ZN(W3541));
  NOR2X1 G9501 (.A1(W630), .A2(W2563), .ZN(W2712));
  NOR2X1 G9502 (.A1(W2177), .A2(W1673), .ZN(W2721));
  NOR2X1 G9503 (.A1(W57), .A2(W708), .ZN(W2720));
  NOR2X1 G9504 (.A1(W414), .A2(W2407), .ZN(W2718));
  NOR2X1 G9505 (.A1(W2426), .A2(I1122), .ZN(W2717));
  NOR2X1 G9506 (.A1(W12924), .A2(W20667), .ZN(W26300));
  NOR2X1 G9507 (.A1(W2426), .A2(I7), .ZN(W2715));
  NOR2X1 G9508 (.A1(W2393), .A2(I0), .ZN(W2714));
  NOR2X1 G9509 (.A1(W23631), .A2(W19184), .ZN(W26299));
  NOR2X1 G9510 (.A1(W17587), .A2(W24381), .ZN(W24444));
  NOR2X1 G9511 (.A1(W16947), .A2(W30855), .ZN(O17166));
  NOR2X1 G9512 (.A1(W1226), .A2(I1465), .ZN(W2710));
  NOR2X1 G9513 (.A1(W149), .A2(W5022), .ZN(O17167));
  NOR2X1 G9514 (.A1(W13724), .A2(W12762), .ZN(O17168));
  NOR2X1 G9515 (.A1(W30276), .A2(W17101), .ZN(O17169));
  NOR2X1 G9516 (.A1(W20129), .A2(W17103), .ZN(W48274));
  NOR2X1 G9517 (.A1(W2539), .A2(I880), .ZN(W2705));
  NOR2X1 G9518 (.A1(W13548), .A2(W15332), .ZN(W26298));
  NOR2X1 G9519 (.A1(W20916), .A2(W5243), .ZN(O17150));
  NOR2X1 G9520 (.A1(W43142), .A2(W28560), .ZN(O17136));
  NOR2X1 G9521 (.A1(W23427), .A2(W15060), .ZN(W24440));
  NOR2X1 G9522 (.A1(W127), .A2(W24380), .ZN(W24441));
  NOR2X1 G9523 (.A1(I1367), .A2(W2646), .ZN(W2735));
  NOR2X1 G9524 (.A1(W11518), .A2(W43352), .ZN(O17142));
  NOR2X1 G9525 (.A1(W922), .A2(W3473), .ZN(W24442));
  NOR2X1 G9526 (.A1(I1300), .A2(W720), .ZN(W2732));
  NOR2X1 G9527 (.A1(W1178), .A2(W35077), .ZN(O17144));
  NOR2X1 G9528 (.A1(W347), .A2(W1004), .ZN(W2702));
  NOR2X1 G9529 (.A1(W42788), .A2(W1139), .ZN(W48254));
  NOR2X1 G9530 (.A1(W17213), .A2(I787), .ZN(O3084));
  NOR2X1 G9531 (.A1(W20313), .A2(W37557), .ZN(W48256));
  NOR2X1 G9532 (.A1(W40047), .A2(W10418), .ZN(O17156));
  NOR2X1 G9533 (.A1(W4583), .A2(W12449), .ZN(O17157));
  NOR2X1 G9534 (.A1(I409), .A2(W2411), .ZN(W2724));
  NOR2X1 G9535 (.A1(W1435), .A2(W42796), .ZN(O17161));
  NOR2X1 G9536 (.A1(W965), .A2(I1382), .ZN(W2674));
  NOR2X1 G9537 (.A1(W2315), .A2(W769), .ZN(W2682));
  NOR2X1 G9538 (.A1(W862), .A2(I1490), .ZN(W2681));
  NOR2X1 G9539 (.A1(W15388), .A2(W11134), .ZN(O17194));
  NOR2X1 G9540 (.A1(I452), .A2(W1363), .ZN(W2679));
  NOR2X1 G9541 (.A1(W1667), .A2(W2583), .ZN(W2678));
  NOR2X1 G9542 (.A1(W848), .A2(W751), .ZN(W2677));
  NOR2X1 G9543 (.A1(W46661), .A2(W19583), .ZN(O17196));
  NOR2X1 G9544 (.A1(W23891), .A2(W4337), .ZN(O3706));
  NOR2X1 G9545 (.A1(W41861), .A2(W31395), .ZN(O17193));
  NOR2X1 G9546 (.A1(W23600), .A2(W22656), .ZN(W26289));
  NOR2X1 G9547 (.A1(W3103), .A2(W16146), .ZN(O17202));
  NOR2X1 G9548 (.A1(W319), .A2(W2105), .ZN(W2671));
  NOR2X1 G9549 (.A1(W7144), .A2(I1260), .ZN(O3089));
  NOR2X1 G9550 (.A1(W42404), .A2(W30525), .ZN(O17205));
  NOR2X1 G9551 (.A1(W30020), .A2(W24109), .ZN(O17207));
  NOR2X1 G9552 (.A1(W9843), .A2(W36444), .ZN(O17208));
  NOR2X1 G9553 (.A1(W9812), .A2(W18479), .ZN(W26287));
  NOR2X1 G9554 (.A1(W1887), .A2(I1738), .ZN(W2691));
  NOR2X1 G9555 (.A1(W266), .A2(I863), .ZN(W2701));
  NOR2X1 G9556 (.A1(W2116), .A2(W12217), .ZN(O17177));
  NOR2X1 G9557 (.A1(W14028), .A2(W18329), .ZN(W26295));
  NOR2X1 G9558 (.A1(W36079), .A2(W28198), .ZN(W48283));
  NOR2X1 G9559 (.A1(I200), .A2(W29487), .ZN(O17180));
  NOR2X1 G9560 (.A1(W33836), .A2(W25121), .ZN(O17182));
  NOR2X1 G9561 (.A1(I1382), .A2(W1803), .ZN(W2694));
  NOR2X1 G9562 (.A1(W2100), .A2(W1658), .ZN(W2693));
  NOR2X1 G9563 (.A1(W9201), .A2(W23040), .ZN(W24439));
  NOR2X1 G9564 (.A1(W1151), .A2(W2284), .ZN(W2690));
  NOR2X1 G9565 (.A1(W37685), .A2(W13506), .ZN(O17185));
  NOR2X1 G9566 (.A1(I1459), .A2(W2636), .ZN(W2688));
  NOR2X1 G9567 (.A1(W10554), .A2(W22992), .ZN(W24453));
  NOR2X1 G9568 (.A1(W8376), .A2(W2422), .ZN(W24454));
  NOR2X1 G9569 (.A1(W15106), .A2(W30316), .ZN(O17191));
  NOR2X1 G9570 (.A1(W24178), .A2(W15515), .ZN(O17192));
  NOR2X1 G9571 (.A1(W14991), .A2(W24175), .ZN(O3078));
  NOR2X1 G9572 (.A1(W225), .A2(W758), .ZN(W2798));
  NOR2X1 G9573 (.A1(W18822), .A2(W1914), .ZN(O17078));
  NOR2X1 G9574 (.A1(W19282), .A2(W39420), .ZN(O17080));
  NOR2X1 G9575 (.A1(W44567), .A2(W20702), .ZN(O17081));
  NOR2X1 G9576 (.A1(W2767), .A2(I355), .ZN(W2794));
  NOR2X1 G9577 (.A1(W1855), .A2(W6341), .ZN(O3719));
  NOR2X1 G9578 (.A1(W18637), .A2(W9397), .ZN(O17084));
  NOR2X1 G9579 (.A1(W44812), .A2(W42344), .ZN(O17085));
  NOR2X1 G9580 (.A1(W17809), .A2(W7394), .ZN(W24415));
  NOR2X1 G9581 (.A1(W7903), .A2(W1951), .ZN(O17087));
  NOR2X1 G9582 (.A1(W46888), .A2(W36667), .ZN(O17088));
  NOR2X1 G9583 (.A1(W943), .A2(I1013), .ZN(W2786));
  NOR2X1 G9584 (.A1(W2512), .A2(W2903), .ZN(W26325));
  NOR2X1 G9585 (.A1(W1053), .A2(W16677), .ZN(O17091));
  NOR2X1 G9586 (.A1(W46122), .A2(W28158), .ZN(O17092));
  NOR2X1 G9587 (.A1(I1522), .A2(W10126), .ZN(O3715));
  NOR2X1 G9588 (.A1(W37130), .A2(W39456), .ZN(O17095));
  NOR2X1 G9589 (.A1(W42236), .A2(W26990), .ZN(O17071));
  NOR2X1 G9590 (.A1(W743), .A2(W559), .ZN(W2816));
  NOR2X1 G9591 (.A1(W33169), .A2(W11250), .ZN(O17063));
  NOR2X1 G9592 (.A1(W13575), .A2(W17162), .ZN(W26332));
  NOR2X1 G9593 (.A1(W83), .A2(W632), .ZN(W2813));
  NOR2X1 G9594 (.A1(W25460), .A2(W44161), .ZN(O17065));
  NOR2X1 G9595 (.A1(I962), .A2(W41117), .ZN(W48160));
  NOR2X1 G9596 (.A1(W1456), .A2(W2427), .ZN(W2810));
  NOR2X1 G9597 (.A1(W8816), .A2(W21208), .ZN(O17069));
  NOR2X1 G9598 (.A1(W26284), .A2(W46968), .ZN(O17096));
  NOR2X1 G9599 (.A1(W3309), .A2(W2384), .ZN(O17072));
  NOR2X1 G9600 (.A1(W10033), .A2(W46867), .ZN(W48165));
  NOR2X1 G9601 (.A1(W18099), .A2(W21132), .ZN(O3720));
  NOR2X1 G9602 (.A1(W384), .A2(W2790), .ZN(W2804));
  NOR2X1 G9603 (.A1(W873), .A2(I136), .ZN(W2803));
  NOR2X1 G9604 (.A1(W36332), .A2(W1306), .ZN(O17075));
  NOR2X1 G9605 (.A1(I207), .A2(I1914), .ZN(W2800));
  NOR2X1 G9606 (.A1(W8500), .A2(W9119), .ZN(W24435));
  NOR2X1 G9607 (.A1(W2579), .A2(W1682), .ZN(W2758));
  NOR2X1 G9608 (.A1(I1100), .A2(W426), .ZN(W2757));
  NOR2X1 G9609 (.A1(W18572), .A2(W6645), .ZN(O17125));
  NOR2X1 G9610 (.A1(W1837), .A2(W1434), .ZN(W2754));
  NOR2X1 G9611 (.A1(I1597), .A2(I1558), .ZN(W2752));
  NOR2X1 G9612 (.A1(W1824), .A2(W903), .ZN(W2751));
  NOR2X1 G9613 (.A1(W0), .A2(W2455), .ZN(W2750));
  NOR2X1 G9614 (.A1(I262), .A2(W2517), .ZN(W2749));
  NOR2X1 G9615 (.A1(W16483), .A2(W5042), .ZN(W26310));
  NOR2X1 G9616 (.A1(W2174), .A2(W12926), .ZN(O3083));
  NOR2X1 G9617 (.A1(W8244), .A2(W8820), .ZN(W24437));
  NOR2X1 G9618 (.A1(I228), .A2(W448), .ZN(W2745));
  NOR2X1 G9619 (.A1(W20112), .A2(W25328), .ZN(O17130));
  NOR2X1 G9620 (.A1(W21416), .A2(W28217), .ZN(O17134));
  NOR2X1 G9621 (.A1(W618), .A2(W1862), .ZN(W2741));
  NOR2X1 G9622 (.A1(I1792), .A2(W39666), .ZN(O17135));
  NOR2X1 G9623 (.A1(W15670), .A2(W43062), .ZN(O17108));
  NOR2X1 G9624 (.A1(W20463), .A2(W12311), .ZN(O3714));
  NOR2X1 G9625 (.A1(I1150), .A2(I1689), .ZN(W2777));
  NOR2X1 G9626 (.A1(W6337), .A2(W5411), .ZN(O17101));
  NOR2X1 G9627 (.A1(W3447), .A2(I118), .ZN(W24423));
  NOR2X1 G9628 (.A1(I1739), .A2(W10543), .ZN(W24424));
  NOR2X1 G9629 (.A1(W45951), .A2(W20959), .ZN(O17105));
  NOR2X1 G9630 (.A1(W28653), .A2(W26861), .ZN(O17106));
  NOR2X1 G9631 (.A1(W1189), .A2(I705), .ZN(W2771));
  NOR2X1 G9632 (.A1(W2221), .A2(W994), .ZN(W2665));
  NOR2X1 G9633 (.A1(W19417), .A2(W5559), .ZN(O3711));
  NOR2X1 G9634 (.A1(W13290), .A2(W10761), .ZN(O3710));
  NOR2X1 G9635 (.A1(W2253), .A2(W1634), .ZN(W2765));
  NOR2X1 G9636 (.A1(W13914), .A2(W8408), .ZN(W26312));
  NOR2X1 G9637 (.A1(W22134), .A2(W19643), .ZN(W26311));
  NOR2X1 G9638 (.A1(W952), .A2(I815), .ZN(W2762));
  NOR2X1 G9639 (.A1(I1881), .A2(W138), .ZN(W2761));
  NOR2X1 G9640 (.A1(W7441), .A2(W10092), .ZN(O17297));
  NOR2X1 G9641 (.A1(W33555), .A2(W3386), .ZN(O17287));
  NOR2X1 G9642 (.A1(W19294), .A2(W9355), .ZN(W26252));
  NOR2X1 G9643 (.A1(I722), .A2(I9), .ZN(W2570));
  NOR2X1 G9644 (.A1(W30203), .A2(W44545), .ZN(O17292));
  NOR2X1 G9645 (.A1(W1079), .A2(W2373), .ZN(W2568));
  NOR2X1 G9646 (.A1(W18793), .A2(W42891), .ZN(O17293));
  NOR2X1 G9647 (.A1(W31360), .A2(W37515), .ZN(O17294));
  NOR2X1 G9648 (.A1(W5647), .A2(W6956), .ZN(W26250));
  NOR2X1 G9649 (.A1(W14380), .A2(W8230), .ZN(O3096));
  NOR2X1 G9650 (.A1(I1386), .A2(W106), .ZN(W2563));
  NOR2X1 G9651 (.A1(W17326), .A2(W47751), .ZN(O17299));
  NOR2X1 G9652 (.A1(W4465), .A2(W37037), .ZN(O17300));
  NOR2X1 G9653 (.A1(W4977), .A2(W3118), .ZN(W24490));
  NOR2X1 G9654 (.A1(W27719), .A2(I1566), .ZN(O17307));
  NOR2X1 G9655 (.A1(I113), .A2(I1695), .ZN(W2557));
  NOR2X1 G9656 (.A1(I975), .A2(W1854), .ZN(W2556));
  NOR2X1 G9657 (.A1(I723), .A2(W136), .ZN(W2555));
  NOR2X1 G9658 (.A1(W38613), .A2(W30794), .ZN(O17280));
  NOR2X1 G9659 (.A1(I410), .A2(W2388), .ZN(W2590));
  NOR2X1 G9660 (.A1(W8429), .A2(W11528), .ZN(W26261));
  NOR2X1 G9661 (.A1(W6674), .A2(W13175), .ZN(O17274));
  NOR2X1 G9662 (.A1(W17102), .A2(W3662), .ZN(O3696));
  NOR2X1 G9663 (.A1(W22458), .A2(W12429), .ZN(W24481));
  NOR2X1 G9664 (.A1(W17444), .A2(W554), .ZN(O3695));
  NOR2X1 G9665 (.A1(W30718), .A2(W37609), .ZN(O17278));
  NOR2X1 G9666 (.A1(W4203), .A2(W11789), .ZN(O17279));
  NOR2X1 G9667 (.A1(W15229), .A2(W4959), .ZN(W24491));
  NOR2X1 G9668 (.A1(W99), .A2(W2040), .ZN(W2581));
  NOR2X1 G9669 (.A1(W22098), .A2(W33497), .ZN(O17281));
  NOR2X1 G9670 (.A1(W39536), .A2(W48325), .ZN(O17282));
  NOR2X1 G9671 (.A1(W35879), .A2(W45490), .ZN(O17283));
  NOR2X1 G9672 (.A1(W9128), .A2(W9534), .ZN(O17285));
  NOR2X1 G9673 (.A1(I1554), .A2(I1722), .ZN(W26255));
  NOR2X1 G9674 (.A1(W11837), .A2(W15139), .ZN(W26254));
  NOR2X1 G9675 (.A1(W18035), .A2(W8259), .ZN(O17341));
  NOR2X1 G9676 (.A1(W20658), .A2(I1773), .ZN(W26233));
  NOR2X1 G9677 (.A1(W13672), .A2(W9393), .ZN(O3686));
  NOR2X1 G9678 (.A1(W22525), .A2(W45211), .ZN(O17337));
  NOR2X1 G9679 (.A1(W124), .A2(W250), .ZN(W2530));
  NOR2X1 G9680 (.A1(W1918), .A2(W1628), .ZN(W2529));
  NOR2X1 G9681 (.A1(I1124), .A2(W35224), .ZN(O17339));
  NOR2X1 G9682 (.A1(W852), .A2(W2319), .ZN(W2527));
  NOR2X1 G9683 (.A1(W6747), .A2(W10761), .ZN(W24503));
  NOR2X1 G9684 (.A1(W37998), .A2(W6600), .ZN(O17333));
  NOR2X1 G9685 (.A1(W20206), .A2(W11503), .ZN(W24505));
  NOR2X1 G9686 (.A1(I906), .A2(W1038), .ZN(W2522));
  NOR2X1 G9687 (.A1(I1535), .A2(I524), .ZN(W2521));
  NOR2X1 G9688 (.A1(W24469), .A2(W13017), .ZN(O17345));
  NOR2X1 G9689 (.A1(W3675), .A2(W10731), .ZN(W48459));
  NOR2X1 G9690 (.A1(W2021), .A2(W1722), .ZN(W2517));
  NOR2X1 G9691 (.A1(W20582), .A2(W23125), .ZN(W24507));
  NOR2X1 G9692 (.A1(W8844), .A2(W24015), .ZN(W26238));
  NOR2X1 G9693 (.A1(I1189), .A2(W955), .ZN(W2553));
  NOR2X1 G9694 (.A1(W14732), .A2(W5814), .ZN(O3693));
  NOR2X1 G9695 (.A1(I862), .A2(I1786), .ZN(W2551));
  NOR2X1 G9696 (.A1(I1296), .A2(I1286), .ZN(W2550));
  NOR2X1 G9697 (.A1(W15041), .A2(W24620), .ZN(W26244));
  NOR2X1 G9698 (.A1(W2534), .A2(W18877), .ZN(W24495));
  NOR2X1 G9699 (.A1(W2284), .A2(I36), .ZN(W2546));
  NOR2X1 G9700 (.A1(W18226), .A2(W46754), .ZN(O17315));
  NOR2X1 G9701 (.A1(W2110), .A2(W21892), .ZN(O17270));
  NOR2X1 G9702 (.A1(W586), .A2(I297), .ZN(W2543));
  NOR2X1 G9703 (.A1(W3759), .A2(I291), .ZN(O17319));
  NOR2X1 G9704 (.A1(W30612), .A2(W27983), .ZN(O17320));
  NOR2X1 G9705 (.A1(W18328), .A2(W24642), .ZN(W26236));
  NOR2X1 G9706 (.A1(W36191), .A2(W20576), .ZN(O17324));
  NOR2X1 G9707 (.A1(W32740), .A2(W6604), .ZN(O17328));
  NOR2X1 G9708 (.A1(W4018), .A2(W9241), .ZN(O3687));
  NOR2X1 G9709 (.A1(W14557), .A2(W47319), .ZN(O17230));
  NOR2X1 G9710 (.A1(W1942), .A2(W251), .ZN(W2647));
  NOR2X1 G9711 (.A1(W799), .A2(I870), .ZN(W2646));
  NOR2X1 G9712 (.A1(W826), .A2(W2519), .ZN(W2645));
  NOR2X1 G9713 (.A1(W2462), .A2(I429), .ZN(W2644));
  NOR2X1 G9714 (.A1(W4043), .A2(W4448), .ZN(W26283));
  NOR2X1 G9715 (.A1(W2172), .A2(I1991), .ZN(W2642));
  NOR2X1 G9716 (.A1(W1541), .A2(W1564), .ZN(O17228));
  NOR2X1 G9717 (.A1(W16725), .A2(I1832), .ZN(W26282));
  NOR2X1 G9718 (.A1(W22328), .A2(W42791), .ZN(O17225));
  NOR2X1 G9719 (.A1(I1117), .A2(W255), .ZN(W2636));
  NOR2X1 G9720 (.A1(W23912), .A2(W5625), .ZN(O17233));
  NOR2X1 G9721 (.A1(W44473), .A2(W370), .ZN(O17234));
  NOR2X1 G9722 (.A1(W16424), .A2(W13050), .ZN(O17237));
  NOR2X1 G9723 (.A1(W38664), .A2(W34944), .ZN(O17238));
  NOR2X1 G9724 (.A1(W6904), .A2(W14597), .ZN(O3701));
  NOR2X1 G9725 (.A1(W8098), .A2(W13204), .ZN(W24468));
  NOR2X1 G9726 (.A1(W34674), .A2(W27184), .ZN(O17243));
  NOR2X1 G9727 (.A1(W3216), .A2(W22783), .ZN(W48325));
  NOR2X1 G9728 (.A1(W30844), .A2(W29676), .ZN(O17211));
  NOR2X1 G9729 (.A1(W12982), .A2(W16262), .ZN(O17212));
  NOR2X1 G9730 (.A1(W22668), .A2(W23707), .ZN(W26286));
  NOR2X1 G9731 (.A1(I1815), .A2(I916), .ZN(W2661));
  NOR2X1 G9732 (.A1(W8102), .A2(W14486), .ZN(W24460));
  NOR2X1 G9733 (.A1(W15888), .A2(W8514), .ZN(W26284));
  NOR2X1 G9734 (.A1(W28841), .A2(W21212), .ZN(O17219));
  NOR2X1 G9735 (.A1(W2437), .A2(W1205), .ZN(W2657));
  NOR2X1 G9736 (.A1(W6720), .A2(W29971), .ZN(W48350));
  NOR2X1 G9737 (.A1(W39), .A2(I1005), .ZN(W2655));
  NOR2X1 G9738 (.A1(W1023), .A2(I1486), .ZN(W2654));
  NOR2X1 G9739 (.A1(W35331), .A2(W33074), .ZN(O17220));
  NOR2X1 G9740 (.A1(W639), .A2(W565), .ZN(W2652));
  NOR2X1 G9741 (.A1(I1722), .A2(W930), .ZN(W2651));
  NOR2X1 G9742 (.A1(W34), .A2(W22095), .ZN(O3091));
  NOR2X1 G9743 (.A1(W40957), .A2(W12110), .ZN(O17224));
  NOR2X1 G9744 (.A1(W25646), .A2(W9898), .ZN(O17263));
  NOR2X1 G9745 (.A1(W1555), .A2(I1436), .ZN(W2609));
  NOR2X1 G9746 (.A1(W2330), .A2(W23), .ZN(W2608));
  NOR2X1 G9747 (.A1(W2484), .A2(W1278), .ZN(W2607));
  NOR2X1 G9748 (.A1(W207), .A2(W1740), .ZN(W26265));
  NOR2X1 G9749 (.A1(W2128), .A2(W1225), .ZN(W2605));
  NOR2X1 G9750 (.A1(I1754), .A2(W2473), .ZN(W2604));
  NOR2X1 G9751 (.A1(I24), .A2(W1221), .ZN(W2603));
  NOR2X1 G9752 (.A1(W5723), .A2(W21696), .ZN(O3094));
  NOR2X1 G9753 (.A1(W667), .A2(W673), .ZN(W2610));
  NOR2X1 G9754 (.A1(W892), .A2(W1600), .ZN(W2600));
  NOR2X1 G9755 (.A1(W47897), .A2(W9166), .ZN(O17265));
  NOR2X1 G9756 (.A1(W38563), .A2(W15473), .ZN(O17266));
  NOR2X1 G9757 (.A1(W19287), .A2(W19224), .ZN(W26262));
  NOR2X1 G9758 (.A1(W1619), .A2(I1522), .ZN(W2594));
  NOR2X1 G9759 (.A1(W5507), .A2(W46052), .ZN(O17269));
  NOR2X1 G9760 (.A1(I603), .A2(W2580), .ZN(W2592));
  NOR2X1 G9761 (.A1(W735), .A2(W3526), .ZN(O17252));
  NOR2X1 G9762 (.A1(W1528), .A2(W2622), .ZN(W2627));
  NOR2X1 G9763 (.A1(W339), .A2(W509), .ZN(W2626));
  NOR2X1 G9764 (.A1(W3185), .A2(W41024), .ZN(O17244));
  NOR2X1 G9765 (.A1(I1818), .A2(I708), .ZN(W2624));
  NOR2X1 G9766 (.A1(W9929), .A2(W7492), .ZN(O3700));
  NOR2X1 G9767 (.A1(W46754), .A2(W35466), .ZN(O17246));
  NOR2X1 G9768 (.A1(W1351), .A2(W831), .ZN(W2621));
  NOR2X1 G9769 (.A1(W30361), .A2(W18939), .ZN(O17249));
  NOR2X1 G9770 (.A1(W46517), .A2(W47504), .ZN(O17061));
  NOR2X1 G9771 (.A1(W4266), .A2(W13461), .ZN(O3699));
  NOR2X1 G9772 (.A1(W25838), .A2(W31155), .ZN(O17254));
  NOR2X1 G9773 (.A1(W28855), .A2(W36351), .ZN(O17255));
  NOR2X1 G9774 (.A1(W16035), .A2(W16581), .ZN(O3093));
  NOR2X1 G9775 (.A1(W9875), .A2(W5567), .ZN(W26267));
  NOR2X1 G9776 (.A1(W27369), .A2(W10987), .ZN(O17259));
  NOR2X1 G9777 (.A1(W26252), .A2(W15418), .ZN(O17260));
  NOR2X1 G9778 (.A1(I1736), .A2(W2550), .ZN(W3025));
  NOR2X1 G9779 (.A1(W17409), .A2(W19949), .ZN(W24337));
  NOR2X1 G9780 (.A1(I1794), .A2(W11429), .ZN(O16869));
  NOR2X1 G9781 (.A1(I1861), .A2(I1358), .ZN(W3031));
  NOR2X1 G9782 (.A1(W587), .A2(W3734), .ZN(W26407));
  NOR2X1 G9783 (.A1(W2605), .A2(W2264), .ZN(W3029));
  NOR2X1 G9784 (.A1(W1908), .A2(W1978), .ZN(W3028));
  NOR2X1 G9785 (.A1(W2323), .A2(W1881), .ZN(W3027));
  NOR2X1 G9786 (.A1(W775), .A2(W1112), .ZN(W3026));
  NOR2X1 G9787 (.A1(W22765), .A2(W5076), .ZN(W24336));
  NOR2X1 G9788 (.A1(W33612), .A2(W39415), .ZN(O16871));
  NOR2X1 G9789 (.A1(W1182), .A2(W666), .ZN(W3022));
  NOR2X1 G9790 (.A1(W40431), .A2(W27865), .ZN(O16876));
  NOR2X1 G9791 (.A1(W1432), .A2(W2188), .ZN(W3020));
  NOR2X1 G9792 (.A1(W19437), .A2(W19058), .ZN(W47952));
  NOR2X1 G9793 (.A1(W14184), .A2(W22810), .ZN(O16877));
  NOR2X1 G9794 (.A1(W7779), .A2(W9918), .ZN(O16878));
  NOR2X1 G9795 (.A1(W44902), .A2(W9939), .ZN(O16879));
  NOR2X1 G9796 (.A1(W31226), .A2(W16605), .ZN(O16860));
  NOR2X1 G9797 (.A1(W22799), .A2(W28734), .ZN(O16854));
  NOR2X1 G9798 (.A1(W36388), .A2(W26380), .ZN(O16855));
  NOR2X1 G9799 (.A1(W21642), .A2(W20472), .ZN(W26409));
  NOR2X1 G9800 (.A1(I967), .A2(W1065), .ZN(W3047));
  NOR2X1 G9801 (.A1(W4504), .A2(W419), .ZN(W24333));
  NOR2X1 G9802 (.A1(W17783), .A2(W15007), .ZN(W24334));
  NOR2X1 G9803 (.A1(W21013), .A2(W42522), .ZN(O16859));
  NOR2X1 G9804 (.A1(I270), .A2(I1533), .ZN(W3043));
  NOR2X1 G9805 (.A1(W41091), .A2(W28215), .ZN(W47957));
  NOR2X1 G9806 (.A1(I874), .A2(I490), .ZN(O27));
  NOR2X1 G9807 (.A1(W425), .A2(I1820), .ZN(W3040));
  NOR2X1 G9808 (.A1(W1611), .A2(I444), .ZN(W3039));
  NOR2X1 G9809 (.A1(W4283), .A2(I1224), .ZN(W26408));
  NOR2X1 G9810 (.A1(W26779), .A2(W11713), .ZN(O16862));
  NOR2X1 G9811 (.A1(W1499), .A2(W2160), .ZN(W3036));
  NOR2X1 G9812 (.A1(W267), .A2(W2015), .ZN(W3035));
  NOR2X1 G9813 (.A1(I38), .A2(I92), .ZN(W2985));
  NOR2X1 G9814 (.A1(W21207), .A2(W14697), .ZN(O16896));
  NOR2X1 G9815 (.A1(W15141), .A2(W345), .ZN(W26399));
  NOR2X1 G9816 (.A1(W1452), .A2(W19349), .ZN(W26398));
  NOR2X1 G9817 (.A1(W40614), .A2(I1646), .ZN(O16899));
  NOR2X1 G9818 (.A1(W2627), .A2(W11503), .ZN(W26397));
  NOR2X1 G9819 (.A1(W30011), .A2(W26793), .ZN(O16901));
  NOR2X1 G9820 (.A1(W14704), .A2(W42616), .ZN(O16903));
  NOR2X1 G9821 (.A1(W2176), .A2(W1401), .ZN(W2986));
  NOR2X1 G9822 (.A1(W22464), .A2(W15343), .ZN(W24345));
  NOR2X1 G9823 (.A1(W669), .A2(W133), .ZN(W2984));
  NOR2X1 G9824 (.A1(I956), .A2(W1529), .ZN(W2983));
  NOR2X1 G9825 (.A1(I1491), .A2(W45108), .ZN(O16904));
  NOR2X1 G9826 (.A1(I1361), .A2(W1309), .ZN(W2981));
  NOR2X1 G9827 (.A1(W796), .A2(W2511), .ZN(W2980));
  NOR2X1 G9828 (.A1(W17778), .A2(W23497), .ZN(O16905));
  NOR2X1 G9829 (.A1(W23426), .A2(W4861), .ZN(W24350));
  NOR2X1 G9830 (.A1(W9980), .A2(W6157), .ZN(O16888));
  NOR2X1 G9831 (.A1(W159), .A2(W2525), .ZN(W3014));
  NOR2X1 G9832 (.A1(W560), .A2(I818), .ZN(W3013));
  NOR2X1 G9833 (.A1(W6423), .A2(W10907), .ZN(W26404));
  NOR2X1 G9834 (.A1(I1704), .A2(I954), .ZN(W3011));
  NOR2X1 G9835 (.A1(W389), .A2(W625), .ZN(W3009));
  NOR2X1 G9836 (.A1(W25788), .A2(W12044), .ZN(O16885));
  NOR2X1 G9837 (.A1(I1231), .A2(W2645), .ZN(W3007));
  NOR2X1 G9838 (.A1(W9409), .A2(W4634), .ZN(W24342));
  NOR2X1 G9839 (.A1(W9296), .A2(W3185), .ZN(W24331));
  NOR2X1 G9840 (.A1(I1976), .A2(W1066), .ZN(W3004));
  NOR2X1 G9841 (.A1(W2907), .A2(W2444), .ZN(W3003));
  NOR2X1 G9842 (.A1(W2637), .A2(W108), .ZN(W3000));
  NOR2X1 G9843 (.A1(W1389), .A2(W1886), .ZN(W2999));
  NOR2X1 G9844 (.A1(W36467), .A2(W36177), .ZN(O16892));
  NOR2X1 G9845 (.A1(W2407), .A2(W1265), .ZN(W2997));
  NOR2X1 G9846 (.A1(W6992), .A2(W18521), .ZN(O16893));
  NOR2X1 G9847 (.A1(W1793), .A2(W3099), .ZN(W3102));
  NOR2X1 G9848 (.A1(W15881), .A2(W31962), .ZN(O16794));
  NOR2X1 G9849 (.A1(W11854), .A2(W7868), .ZN(O16797));
  NOR2X1 G9850 (.A1(W24240), .A2(W18383), .ZN(O3754));
  NOR2X1 G9851 (.A1(W11871), .A2(I1843), .ZN(W26431));
  NOR2X1 G9852 (.A1(W1322), .A2(I303), .ZN(W3108));
  NOR2X1 G9853 (.A1(W1917), .A2(I1712), .ZN(W3107));
  NOR2X1 G9854 (.A1(I1298), .A2(W795), .ZN(W3106));
  NOR2X1 G9855 (.A1(I223), .A2(I514), .ZN(W3104));
  NOR2X1 G9856 (.A1(W33372), .A2(W33560), .ZN(O16793));
  NOR2X1 G9857 (.A1(W44814), .A2(W28571), .ZN(O16805));
  NOR2X1 G9858 (.A1(W9800), .A2(W17717), .ZN(W24315));
  NOR2X1 G9859 (.A1(W20564), .A2(W1224), .ZN(W24316));
  NOR2X1 G9860 (.A1(W25864), .A2(W3213), .ZN(W47877));
  NOR2X1 G9861 (.A1(W20), .A2(W139), .ZN(W3097));
  NOR2X1 G9862 (.A1(W11360), .A2(W41700), .ZN(O16810));
  NOR2X1 G9863 (.A1(W23510), .A2(W645), .ZN(O3752));
  NOR2X1 G9864 (.A1(W19145), .A2(W19708), .ZN(W26425));
  NOR2X1 G9865 (.A1(W23689), .A2(W19257), .ZN(W26436));
  NOR2X1 G9866 (.A1(W2207), .A2(W30320), .ZN(O16778));
  NOR2X1 G9867 (.A1(W3579), .A2(W6037), .ZN(O16784));
  NOR2X1 G9868 (.A1(W24732), .A2(W29474), .ZN(O16787));
  NOR2X1 G9869 (.A1(W1141), .A2(W5326), .ZN(W24306));
  NOR2X1 G9870 (.A1(I1222), .A2(W602), .ZN(W3125));
  NOR2X1 G9871 (.A1(W2704), .A2(W415), .ZN(W3124));
  NOR2X1 G9872 (.A1(W717), .A2(I1326), .ZN(W3123));
  NOR2X1 G9873 (.A1(I1221), .A2(I697), .ZN(W3122));
  NOR2X1 G9874 (.A1(W15567), .A2(W44383), .ZN(O16814));
  NOR2X1 G9875 (.A1(W20259), .A2(W15768), .ZN(W24308));
  NOR2X1 G9876 (.A1(W1627), .A2(W2868), .ZN(W3119));
  NOR2X1 G9877 (.A1(W2770), .A2(W1170), .ZN(W3118));
  NOR2X1 G9878 (.A1(W25458), .A2(W4840), .ZN(O3755));
  NOR2X1 G9879 (.A1(W29611), .A2(W9029), .ZN(O16792));
  NOR2X1 G9880 (.A1(W6139), .A2(W11395), .ZN(O3041));
  NOR2X1 G9881 (.A1(I1204), .A2(W920), .ZN(W3114));
  NOR2X1 G9882 (.A1(I337), .A2(I1495), .ZN(W3060));
  NOR2X1 G9883 (.A1(W2583), .A2(I206), .ZN(W3072));
  NOR2X1 G9884 (.A1(I303), .A2(W2748), .ZN(W3069));
  NOR2X1 G9885 (.A1(W28028), .A2(W7290), .ZN(O16837));
  NOR2X1 G9886 (.A1(W2691), .A2(W1005), .ZN(W3066));
  NOR2X1 G9887 (.A1(W16119), .A2(W28327), .ZN(O16839));
  NOR2X1 G9888 (.A1(W13981), .A2(W40461), .ZN(O16841));
  NOR2X1 G9889 (.A1(W45371), .A2(W19186), .ZN(O16842));
  NOR2X1 G9890 (.A1(I904), .A2(W40317), .ZN(O16844));
  NOR2X1 G9891 (.A1(W7136), .A2(W3197), .ZN(O3748));
  NOR2X1 G9892 (.A1(W1302), .A2(I1629), .ZN(W3059));
  NOR2X1 G9893 (.A1(W21941), .A2(W10905), .ZN(W26411));
  NOR2X1 G9894 (.A1(W2735), .A2(W1555), .ZN(W3057));
  NOR2X1 G9895 (.A1(W628), .A2(I1392), .ZN(W3056));
  NOR2X1 G9896 (.A1(W1880), .A2(W2647), .ZN(W3054));
  NOR2X1 G9897 (.A1(W2027), .A2(I1240), .ZN(W3053));
  NOR2X1 G9898 (.A1(W37679), .A2(W14062), .ZN(O16849));
  NOR2X1 G9899 (.A1(I316), .A2(I1927), .ZN(W3081));
  NOR2X1 G9900 (.A1(I687), .A2(W5592), .ZN(O16816));
  NOR2X1 G9901 (.A1(W6793), .A2(W29771), .ZN(O16817));
  NOR2X1 G9902 (.A1(W43535), .A2(W41757), .ZN(O16818));
  NOR2X1 G9903 (.A1(W32888), .A2(W46511), .ZN(W47892));
  NOR2X1 G9904 (.A1(W1873), .A2(I1758), .ZN(W3086));
  NOR2X1 G9905 (.A1(W6476), .A2(W6602), .ZN(O16821));
  NOR2X1 G9906 (.A1(W22637), .A2(W22688), .ZN(O16822));
  NOR2X1 G9907 (.A1(I1748), .A2(W6708), .ZN(O3043));
  NOR2X1 G9908 (.A1(W21434), .A2(W5657), .ZN(O16907));
  NOR2X1 G9909 (.A1(I1425), .A2(W406), .ZN(W3080));
  NOR2X1 G9910 (.A1(W2703), .A2(W147), .ZN(W3079));
  NOR2X1 G9911 (.A1(W11441), .A2(W44581), .ZN(O16826));
  NOR2X1 G9912 (.A1(W5630), .A2(W23674), .ZN(W26422));
  NOR2X1 G9913 (.A1(W369), .A2(I469), .ZN(W3076));
  NOR2X1 G9914 (.A1(W277), .A2(W519), .ZN(W3075));
  NOR2X1 G9915 (.A1(W28091), .A2(W32295), .ZN(O16828));
  NOR2X1 G9916 (.A1(W2406), .A2(I772), .ZN(W2866));
  NOR2X1 G9917 (.A1(W5688), .A2(W34603), .ZN(O17009));
  NOR2X1 G9918 (.A1(I1502), .A2(I827), .ZN(W2874));
  NOR2X1 G9919 (.A1(W47375), .A2(W42928), .ZN(O17010));
  NOR2X1 G9920 (.A1(W24649), .A2(W4292), .ZN(W26355));
  NOR2X1 G9921 (.A1(W1197), .A2(W34335), .ZN(O17016));
  NOR2X1 G9922 (.A1(W2634), .A2(W229), .ZN(W2870));
  NOR2X1 G9923 (.A1(W30755), .A2(W12108), .ZN(O17018));
  NOR2X1 G9924 (.A1(I208), .A2(I1274), .ZN(W2868));
  NOR2X1 G9925 (.A1(I626), .A2(I1141), .ZN(W2876));
  NOR2X1 G9926 (.A1(I1189), .A2(W1643), .ZN(W2864));
  NOR2X1 G9927 (.A1(W40194), .A2(W7176), .ZN(O17023));
  NOR2X1 G9928 (.A1(W38348), .A2(W5738), .ZN(O17024));
  NOR2X1 G9929 (.A1(W1480), .A2(W27024), .ZN(O17025));
  NOR2X1 G9930 (.A1(W3305), .A2(W40000), .ZN(O17026));
  NOR2X1 G9931 (.A1(W20829), .A2(W11500), .ZN(W26351));
  NOR2X1 G9932 (.A1(W15705), .A2(W15417), .ZN(W24396));
  NOR2X1 G9933 (.A1(W596), .A2(W528), .ZN(W2857));
  NOR2X1 G9934 (.A1(W953), .A2(I285), .ZN(W2884));
  NOR2X1 G9935 (.A1(W2616), .A2(I552), .ZN(W2894));
  NOR2X1 G9936 (.A1(W46987), .A2(W37722), .ZN(W48074));
  NOR2X1 G9937 (.A1(W8312), .A2(W9583), .ZN(O16991));
  NOR2X1 G9938 (.A1(W45766), .A2(W37411), .ZN(O16992));
  NOR2X1 G9939 (.A1(W8095), .A2(W9455), .ZN(W24385));
  NOR2X1 G9940 (.A1(W6127), .A2(W17816), .ZN(O3068));
  NOR2X1 G9941 (.A1(I194), .A2(I1301), .ZN(W2888));
  NOR2X1 G9942 (.A1(W23548), .A2(W20767), .ZN(O16998));
  NOR2X1 G9943 (.A1(W6540), .A2(W18454), .ZN(W24397));
  NOR2X1 G9944 (.A1(W1193), .A2(W13327), .ZN(O3729));
  NOR2X1 G9945 (.A1(W8918), .A2(W18561), .ZN(W48087));
  NOR2X1 G9946 (.A1(W5090), .A2(W1332), .ZN(W26358));
  NOR2X1 G9947 (.A1(W165), .A2(I432), .ZN(W2880));
  NOR2X1 G9948 (.A1(W11517), .A2(W15187), .ZN(W24391));
  NOR2X1 G9949 (.A1(I310), .A2(W2584), .ZN(W2878));
  NOR2X1 G9950 (.A1(W28771), .A2(W27625), .ZN(O17008));
  NOR2X1 G9951 (.A1(W46345), .A2(W32995), .ZN(W48145));
  NOR2X1 G9952 (.A1(W11335), .A2(W11570), .ZN(W26342));
  NOR2X1 G9953 (.A1(W21764), .A2(W9074), .ZN(O3725));
  NOR2X1 G9954 (.A1(W8497), .A2(W20211), .ZN(W24407));
  NOR2X1 G9955 (.A1(I702), .A2(W134), .ZN(W2832));
  NOR2X1 G9956 (.A1(W19082), .A2(W6743), .ZN(W26337));
  NOR2X1 G9957 (.A1(W29880), .A2(W3558), .ZN(O17052));
  NOR2X1 G9958 (.A1(I1289), .A2(W2404), .ZN(W2829));
  NOR2X1 G9959 (.A1(W5221), .A2(W4197), .ZN(W24409));
  NOR2X1 G9960 (.A1(W7754), .A2(W9756), .ZN(W26343));
  NOR2X1 G9961 (.A1(W18942), .A2(W1224), .ZN(O17057));
  NOR2X1 G9962 (.A1(I6), .A2(W2532), .ZN(W2825));
  NOR2X1 G9963 (.A1(W24069), .A2(I1021), .ZN(W48147));
  NOR2X1 G9964 (.A1(W5838), .A2(W11817), .ZN(W48148));
  NOR2X1 G9965 (.A1(W1225), .A2(W1699), .ZN(W2821));
  NOR2X1 G9966 (.A1(W913), .A2(W2811), .ZN(W2820));
  NOR2X1 G9967 (.A1(W5190), .A2(W8547), .ZN(O17059));
  NOR2X1 G9968 (.A1(I1908), .A2(W2101), .ZN(W2847));
  NOR2X1 G9969 (.A1(I792), .A2(W257), .ZN(W2855));
  NOR2X1 G9970 (.A1(W20265), .A2(W9837), .ZN(W24398));
  NOR2X1 G9971 (.A1(W2646), .A2(W2283), .ZN(W2853));
  NOR2X1 G9972 (.A1(W21199), .A2(W19523), .ZN(W26350));
  NOR2X1 G9973 (.A1(W502), .A2(I496), .ZN(W2851));
  NOR2X1 G9974 (.A1(W17504), .A2(W18849), .ZN(O17036));
  NOR2X1 G9975 (.A1(W2275), .A2(W19192), .ZN(W24400));
  NOR2X1 G9976 (.A1(I1858), .A2(I491), .ZN(W2848));
  NOR2X1 G9977 (.A1(W6869), .A2(W3800), .ZN(W26364));
  NOR2X1 G9978 (.A1(I1054), .A2(W1007), .ZN(W2845));
  NOR2X1 G9979 (.A1(W866), .A2(W612), .ZN(W2844));
  NOR2X1 G9980 (.A1(I706), .A2(W182), .ZN(W2843));
  NOR2X1 G9981 (.A1(I493), .A2(I1296), .ZN(W2842));
  NOR2X1 G9982 (.A1(I5), .A2(W163), .ZN(W2841));
  NOR2X1 G9983 (.A1(W557), .A2(W1451), .ZN(W2839));
  NOR2X1 G9984 (.A1(W7776), .A2(W13419), .ZN(O17041));
  NOR2X1 G9985 (.A1(W35457), .A2(W7489), .ZN(O16941));
  NOR2X1 G9986 (.A1(W23097), .A2(W14502), .ZN(W26384));
  NOR2X1 G9987 (.A1(W44504), .A2(W18137), .ZN(O16933));
  NOR2X1 G9988 (.A1(W12195), .A2(W6534), .ZN(O3057));
  NOR2X1 G9989 (.A1(W36099), .A2(W9273), .ZN(O16935));
  NOR2X1 G9990 (.A1(W429), .A2(W633), .ZN(W2950));
  NOR2X1 G9991 (.A1(I156), .A2(W1490), .ZN(W2949));
  NOR2X1 G9992 (.A1(W552), .A2(W18106), .ZN(O16936));
  NOR2X1 G9993 (.A1(W15989), .A2(W22227), .ZN(O3058));
  NOR2X1 G9994 (.A1(I1669), .A2(W1000), .ZN(W2955));
  NOR2X1 G9995 (.A1(W19452), .A2(W9537), .ZN(O3734));
  NOR2X1 G9996 (.A1(W1445), .A2(I1712), .ZN(W2943));
  NOR2X1 G9997 (.A1(W11204), .A2(W24424), .ZN(O16943));
  NOR2X1 G9998 (.A1(W2643), .A2(W282), .ZN(W2941));
  NOR2X1 G9999 (.A1(W573), .A2(W2515), .ZN(W2939));
  NOR2X1 G10000 (.A1(I1509), .A2(W971), .ZN(W2938));
  NOR2X1 G10001 (.A1(W38505), .A2(W3893), .ZN(O16945));
  NOR2X1 G10002 (.A1(W2340), .A2(W457), .ZN(W2935));
  NOR2X1 G10003 (.A1(W2815), .A2(W1843), .ZN(W2966));
  NOR2X1 G10004 (.A1(W2572), .A2(W2176), .ZN(W2976));
  NOR2X1 G10005 (.A1(I1890), .A2(W1571), .ZN(W2974));
  NOR2X1 G10006 (.A1(W1587), .A2(W21859), .ZN(W26393));
  NOR2X1 G10007 (.A1(W11163), .A2(W8431), .ZN(O16912));
  NOR2X1 G10008 (.A1(W13008), .A2(W5176), .ZN(O3742));
  NOR2X1 G10009 (.A1(W5301), .A2(W16729), .ZN(W26390));
  NOR2X1 G10010 (.A1(W15511), .A2(W1670), .ZN(O3741));
  NOR2X1 G10011 (.A1(W8805), .A2(W22220), .ZN(O3740));
  NOR2X1 G10012 (.A1(W1988), .A2(I1308), .ZN(W2934));
  NOR2X1 G10013 (.A1(I1516), .A2(W2746), .ZN(W2964));
  NOR2X1 G10014 (.A1(W3201), .A2(W24295), .ZN(O3055));
  NOR2X1 G10015 (.A1(W1320), .A2(W53), .ZN(W2961));
  NOR2X1 G10016 (.A1(W2684), .A2(I448), .ZN(W2960));
  NOR2X1 G10017 (.A1(W38678), .A2(W13718), .ZN(O16925));
  NOR2X1 G10018 (.A1(W10752), .A2(W2435), .ZN(O16926));
  NOR2X1 G10019 (.A1(W2266), .A2(W3836), .ZN(W24362));
  NOR2X1 G10020 (.A1(W74), .A2(W323), .ZN(W2903));
  NOR2X1 G10021 (.A1(I1540), .A2(W1234), .ZN(W2913));
  NOR2X1 G10022 (.A1(I731), .A2(W1309), .ZN(W2912));
  NOR2X1 G10023 (.A1(W5545), .A2(W904), .ZN(W24378));
  NOR2X1 G10024 (.A1(W650), .A2(W88), .ZN(W2910));
  NOR2X1 G10025 (.A1(W1243), .A2(W959), .ZN(W2908));
  NOR2X1 G10026 (.A1(W11977), .A2(W2643), .ZN(O16979));
  NOR2X1 G10027 (.A1(W1923), .A2(I1953), .ZN(O26));
  NOR2X1 G10028 (.A1(W4448), .A2(W21114), .ZN(W48063));
  NOR2X1 G10029 (.A1(W25789), .A2(W17794), .ZN(O16972));
  NOR2X1 G10030 (.A1(W5948), .A2(W16856), .ZN(W26365));
  NOR2X1 G10031 (.A1(W1691), .A2(I1416), .ZN(W2901));
  NOR2X1 G10032 (.A1(W6324), .A2(W8687), .ZN(O3067));
  NOR2X1 G10033 (.A1(W46036), .A2(W19433), .ZN(O16986));
  NOR2X1 G10034 (.A1(I772), .A2(W792), .ZN(W2898));
  NOR2X1 G10035 (.A1(W25184), .A2(I1544), .ZN(O16988));
  NOR2X1 G10036 (.A1(W21039), .A2(W16004), .ZN(W24383));
  NOR2X1 G10037 (.A1(W5725), .A2(W37973), .ZN(O16961));
  NOR2X1 G10038 (.A1(W22515), .A2(W34346), .ZN(O16950));
  NOR2X1 G10039 (.A1(W18194), .A2(W22833), .ZN(O3732));
  NOR2X1 G10040 (.A1(W33938), .A2(W30827), .ZN(O16952));
  NOR2X1 G10041 (.A1(W1734), .A2(W1140), .ZN(W2928));
  NOR2X1 G10042 (.A1(W976), .A2(W966), .ZN(W2927));
  NOR2X1 G10043 (.A1(W2578), .A2(I536), .ZN(W2925));
  NOR2X1 G10044 (.A1(W14362), .A2(W2363), .ZN(W24374));
  NOR2X1 G10045 (.A1(W17094), .A2(W5525), .ZN(W26369));
  NOR2X1 G10046 (.A1(W45988), .A2(W5382), .ZN(W47214));
  NOR2X1 G10047 (.A1(W28534), .A2(W2584), .ZN(O16962));
  NOR2X1 G10048 (.A1(I245), .A2(W1627), .ZN(W2920));
  NOR2X1 G10049 (.A1(W3240), .A2(W13723), .ZN(W24376));
  NOR2X1 G10050 (.A1(W1261), .A2(W383), .ZN(W24377));
  NOR2X1 G10051 (.A1(W11683), .A2(W43453), .ZN(O16968));
  NOR2X1 G10052 (.A1(W36716), .A2(W39271), .ZN(O16969));
  NOR2X1 G10053 (.A1(W35282), .A2(W28490), .ZN(O16971));
  NOR2X1 G10054 (.A1(W2413), .A2(W27986), .ZN(O15553));
  NOR2X1 G10055 (.A1(W3456), .A2(W4273), .ZN(W4590));
  NOR2X1 G10056 (.A1(W46229), .A2(W30409), .ZN(O15547));
  NOR2X1 G10057 (.A1(W2438), .A2(I614), .ZN(W4588));
  NOR2X1 G10058 (.A1(W14113), .A2(W14832), .ZN(O15548));
  NOR2X1 G10059 (.A1(I1770), .A2(I1090), .ZN(W4585));
  NOR2X1 G10060 (.A1(W19042), .A2(W12009), .ZN(W23836));
  NOR2X1 G10061 (.A1(I1495), .A2(I1399), .ZN(W4583));
  NOR2X1 G10062 (.A1(W22840), .A2(I1139), .ZN(W26878));
  NOR2X1 G10063 (.A1(W9956), .A2(W15971), .ZN(W23834));
  NOR2X1 G10064 (.A1(W1146), .A2(W725), .ZN(W4580));
  NOR2X1 G10065 (.A1(W689), .A2(W2375), .ZN(W4579));
  NOR2X1 G10066 (.A1(W18426), .A2(W20556), .ZN(W23838));
  NOR2X1 G10067 (.A1(W4253), .A2(I285), .ZN(W4577));
  NOR2X1 G10068 (.A1(W33893), .A2(W14052), .ZN(O15555));
  NOR2X1 G10069 (.A1(I1401), .A2(W3573), .ZN(W4575));
  NOR2X1 G10070 (.A1(W34254), .A2(W13283), .ZN(O15561));
  NOR2X1 G10071 (.A1(W42908), .A2(W21198), .ZN(O15562));
  NOR2X1 G10072 (.A1(W4044), .A2(W1238), .ZN(W4599));
  NOR2X1 G10073 (.A1(I1708), .A2(W2031), .ZN(W4608));
  NOR2X1 G10074 (.A1(W1649), .A2(W2731), .ZN(W4607));
  NOR2X1 G10075 (.A1(W19011), .A2(W4926), .ZN(O3907));
  NOR2X1 G10076 (.A1(W4078), .A2(W3864), .ZN(W4605));
  NOR2X1 G10077 (.A1(W1531), .A2(I1024), .ZN(W4604));
  NOR2X1 G10078 (.A1(W2132), .A2(W3020), .ZN(W4603));
  NOR2X1 G10079 (.A1(I1979), .A2(W4110), .ZN(W4602));
  NOR2X1 G10080 (.A1(W16790), .A2(W10166), .ZN(O3906));
  NOR2X1 G10081 (.A1(W3987), .A2(W709), .ZN(W4569));
  NOR2X1 G10082 (.A1(W16739), .A2(W8220), .ZN(O15538));
  NOR2X1 G10083 (.A1(W15142), .A2(W22807), .ZN(O3903));
  NOR2X1 G10084 (.A1(W26444), .A2(W24423), .ZN(W26882));
  NOR2X1 G10085 (.A1(W645), .A2(W29040), .ZN(W46432));
  NOR2X1 G10086 (.A1(W34121), .A2(W36602), .ZN(O15542));
  NOR2X1 G10087 (.A1(W32568), .A2(W29705), .ZN(O15543));
  NOR2X1 G10088 (.A1(W20527), .A2(W11609), .ZN(W23833));
  NOR2X1 G10089 (.A1(W3219), .A2(I652), .ZN(W4541));
  NOR2X1 G10090 (.A1(W23612), .A2(W2485), .ZN(W26870));
  NOR2X1 G10091 (.A1(W488), .A2(W24765), .ZN(W46473));
  NOR2X1 G10092 (.A1(W279), .A2(W1292), .ZN(W4547));
  NOR2X1 G10093 (.A1(W34930), .A2(W25013), .ZN(O15581));
  NOR2X1 G10094 (.A1(W35238), .A2(W42431), .ZN(O15583));
  NOR2X1 G10095 (.A1(W3806), .A2(W2007), .ZN(W4544));
  NOR2X1 G10096 (.A1(W35111), .A2(W4865), .ZN(O15584));
  NOR2X1 G10097 (.A1(I604), .A2(W2963), .ZN(W4542));
  NOR2X1 G10098 (.A1(W1998), .A2(W4340), .ZN(W4551));
  NOR2X1 G10099 (.A1(W2545), .A2(W23399), .ZN(O15586));
  NOR2X1 G10100 (.A1(W42927), .A2(W37650), .ZN(W46486));
  NOR2X1 G10101 (.A1(W7306), .A2(W38137), .ZN(O15591));
  NOR2X1 G10102 (.A1(W42030), .A2(W2233), .ZN(O15593));
  NOR2X1 G10103 (.A1(W39469), .A2(W33384), .ZN(O15594));
  NOR2X1 G10104 (.A1(W35529), .A2(W3349), .ZN(O15595));
  NOR2X1 G10105 (.A1(W635), .A2(I1565), .ZN(W4533));
  NOR2X1 G10106 (.A1(W4521), .A2(W22159), .ZN(W23849));
  NOR2X1 G10107 (.A1(W16215), .A2(W45564), .ZN(O15571));
  NOR2X1 G10108 (.A1(W8892), .A2(W5800), .ZN(O2896));
  NOR2X1 G10109 (.A1(W37373), .A2(W5885), .ZN(O15565));
  NOR2X1 G10110 (.A1(W7576), .A2(W5698), .ZN(O15567));
  NOR2X1 G10111 (.A1(W744), .A2(W583), .ZN(W4565));
  NOR2X1 G10112 (.A1(W9265), .A2(W14947), .ZN(O15568));
  NOR2X1 G10113 (.A1(W412), .A2(W2454), .ZN(W4563));
  NOR2X1 G10114 (.A1(W8231), .A2(W39988), .ZN(O15569));
  NOR2X1 G10115 (.A1(W4441), .A2(W33799), .ZN(O15570));
  NOR2X1 G10116 (.A1(W385), .A2(W3400), .ZN(W4609));
  NOR2X1 G10117 (.A1(W3110), .A2(W8672), .ZN(O2897));
  NOR2X1 G10118 (.A1(W5305), .A2(W6309), .ZN(O15575));
  NOR2X1 G10119 (.A1(W13269), .A2(W18605), .ZN(O2898));
  NOR2X1 G10120 (.A1(W1248), .A2(I1606), .ZN(W4555));
  NOR2X1 G10121 (.A1(W956), .A2(I315), .ZN(W4554));
  NOR2X1 G10122 (.A1(W20405), .A2(W24164), .ZN(O15577));
  NOR2X1 G10123 (.A1(I1856), .A2(W1824), .ZN(W4552));
  NOR2X1 G10124 (.A1(W1055), .A2(I1959), .ZN(W4659));
  NOR2X1 G10125 (.A1(W10180), .A2(W19652), .ZN(O3917));
  NOR2X1 G10126 (.A1(W3255), .A2(W2186), .ZN(W4667));
  NOR2X1 G10127 (.A1(W15333), .A2(W19114), .ZN(W23802));
  NOR2X1 G10128 (.A1(W3355), .A2(W1214), .ZN(W4665));
  NOR2X1 G10129 (.A1(W17794), .A2(W30085), .ZN(O15489));
  NOR2X1 G10130 (.A1(W22353), .A2(W24634), .ZN(W26911));
  NOR2X1 G10131 (.A1(W1558), .A2(W11250), .ZN(W26909));
  NOR2X1 G10132 (.A1(W2805), .A2(W1924), .ZN(W4661));
  NOR2X1 G10133 (.A1(W4313), .A2(W3266), .ZN(W4669));
  NOR2X1 G10134 (.A1(W19043), .A2(W26514), .ZN(O15492));
  NOR2X1 G10135 (.A1(I1416), .A2(W593), .ZN(W26906));
  NOR2X1 G10136 (.A1(W11656), .A2(W154), .ZN(O2886));
  NOR2X1 G10137 (.A1(W6096), .A2(W1912), .ZN(O15499));
  NOR2X1 G10138 (.A1(W25239), .A2(W16406), .ZN(W26904));
  NOR2X1 G10139 (.A1(I112), .A2(W2377), .ZN(W4652));
  NOR2X1 G10140 (.A1(W10762), .A2(W19983), .ZN(W23810));
  NOR2X1 G10141 (.A1(W39973), .A2(W20749), .ZN(O15502));
  NOR2X1 G10142 (.A1(W17290), .A2(W14419), .ZN(O2884));
  NOR2X1 G10143 (.A1(I1194), .A2(W1565), .ZN(W4688));
  NOR2X1 G10144 (.A1(W42926), .A2(W45225), .ZN(O15474));
  NOR2X1 G10145 (.A1(W734), .A2(W4274), .ZN(W4685));
  NOR2X1 G10146 (.A1(W35204), .A2(W35687), .ZN(O15475));
  NOR2X1 G10147 (.A1(W6348), .A2(W23814), .ZN(O15480));
  NOR2X1 G10148 (.A1(W2242), .A2(W1047), .ZN(W4680));
  NOR2X1 G10149 (.A1(W44158), .A2(W10524), .ZN(W46360));
  NOR2X1 G10150 (.A1(W1782), .A2(W42273), .ZN(W46361));
  NOR2X1 G10151 (.A1(W23982), .A2(W3350), .ZN(O15503));
  NOR2X1 G10152 (.A1(W1275), .A2(W526), .ZN(W4676));
  NOR2X1 G10153 (.A1(W2768), .A2(W3223), .ZN(W4675));
  NOR2X1 G10154 (.A1(W1595), .A2(W2135), .ZN(W4674));
  NOR2X1 G10155 (.A1(W37439), .A2(W19984), .ZN(O15483));
  NOR2X1 G10156 (.A1(W385), .A2(W1804), .ZN(W4672));
  NOR2X1 G10157 (.A1(W1922), .A2(W748), .ZN(W4671));
  NOR2X1 G10158 (.A1(W1591), .A2(W3802), .ZN(W23800));
  NOR2X1 G10159 (.A1(I1386), .A2(I613), .ZN(W4618));
  NOR2X1 G10160 (.A1(I454), .A2(I120), .ZN(W4628));
  NOR2X1 G10161 (.A1(W45919), .A2(W1711), .ZN(O15522));
  NOR2X1 G10162 (.A1(W647), .A2(W1207), .ZN(W4626));
  NOR2X1 G10163 (.A1(W1749), .A2(W3462), .ZN(W4624));
  NOR2X1 G10164 (.A1(W3815), .A2(W6274), .ZN(W26894));
  NOR2X1 G10165 (.A1(W2064), .A2(W3528), .ZN(W4622));
  NOR2X1 G10166 (.A1(W2682), .A2(W2906), .ZN(W4621));
  NOR2X1 G10167 (.A1(W16325), .A2(W22263), .ZN(W46415));
  NOR2X1 G10168 (.A1(W35719), .A2(W29879), .ZN(O15521));
  NOR2X1 G10169 (.A1(W53), .A2(W11116), .ZN(O15528));
  NOR2X1 G10170 (.A1(W3231), .A2(W1456), .ZN(W4616));
  NOR2X1 G10171 (.A1(W7822), .A2(W231), .ZN(W26891));
  NOR2X1 G10172 (.A1(W22135), .A2(W44474), .ZN(O15531));
  NOR2X1 G10173 (.A1(W4907), .A2(W14562), .ZN(W23826));
  NOR2X1 G10174 (.A1(W13770), .A2(W29061), .ZN(W46422));
  NOR2X1 G10175 (.A1(W1148), .A2(W601), .ZN(W4610));
  NOR2X1 G10176 (.A1(W29633), .A2(W29052), .ZN(O15511));
  NOR2X1 G10177 (.A1(W7700), .A2(W15856), .ZN(W23812));
  NOR2X1 G10178 (.A1(W4814), .A2(W25204), .ZN(W26902));
  NOR2X1 G10179 (.A1(W113), .A2(I468), .ZN(W4645));
  NOR2X1 G10180 (.A1(W3507), .A2(W1521), .ZN(W4644));
  NOR2X1 G10181 (.A1(W21668), .A2(W22828), .ZN(W23814));
  NOR2X1 G10182 (.A1(W2968), .A2(I226), .ZN(W4642));
  NOR2X1 G10183 (.A1(W6680), .A2(W4657), .ZN(W23815));
  NOR2X1 G10184 (.A1(I866), .A2(I1928), .ZN(W4640));
  NOR2X1 G10185 (.A1(W40905), .A2(W18843), .ZN(O15597));
  NOR2X1 G10186 (.A1(W592), .A2(I603), .ZN(W4637));
  NOR2X1 G10187 (.A1(W12524), .A2(W15053), .ZN(O2888));
  NOR2X1 G10188 (.A1(W2919), .A2(W4472), .ZN(W4635));
  NOR2X1 G10189 (.A1(W2419), .A2(W3995), .ZN(O2889));
  NOR2X1 G10190 (.A1(W16869), .A2(W15449), .ZN(O3913));
  NOR2X1 G10191 (.A1(W320), .A2(I370), .ZN(W4632));
  NOR2X1 G10192 (.A1(W14107), .A2(W2497), .ZN(W23821));
  NOR2X1 G10193 (.A1(W1713), .A2(W28792), .ZN(W46587));
  NOR2X1 G10194 (.A1(W24555), .A2(W7073), .ZN(O3886));
  NOR2X1 G10195 (.A1(W7153), .A2(W24444), .ZN(O15668));
  NOR2X1 G10196 (.A1(W19484), .A2(W19897), .ZN(O2915));
  NOR2X1 G10197 (.A1(W464), .A2(W1763), .ZN(W4428));
  NOR2X1 G10198 (.A1(W10210), .A2(W13620), .ZN(O15670));
  NOR2X1 G10199 (.A1(W32348), .A2(W7310), .ZN(O15671));
  NOR2X1 G10200 (.A1(I644), .A2(I768), .ZN(O3885));
  NOR2X1 G10201 (.A1(W2634), .A2(I14), .ZN(W4423));
  NOR2X1 G10202 (.A1(W3442), .A2(W2894), .ZN(W4432));
  NOR2X1 G10203 (.A1(W14617), .A2(W20402), .ZN(O15675));
  NOR2X1 G10204 (.A1(W38717), .A2(W16936), .ZN(O15677));
  NOR2X1 G10205 (.A1(W4214), .A2(W3294), .ZN(O15678));
  NOR2X1 G10206 (.A1(W39181), .A2(W21477), .ZN(W46595));
  NOR2X1 G10207 (.A1(W3399), .A2(W3332), .ZN(W4414));
  NOR2X1 G10208 (.A1(W143), .A2(W4332), .ZN(W4413));
  NOR2X1 G10209 (.A1(W2724), .A2(W4205), .ZN(W4412));
  NOR2X1 G10210 (.A1(W767), .A2(W2888), .ZN(W4410));
  NOR2X1 G10211 (.A1(W752), .A2(I779), .ZN(W4441));
  NOR2X1 G10212 (.A1(W2290), .A2(I1392), .ZN(W4452));
  NOR2X1 G10213 (.A1(W13357), .A2(W26467), .ZN(O11981));
  NOR2X1 G10214 (.A1(W26632), .A2(W24907), .ZN(W26835));
  NOR2X1 G10215 (.A1(I679), .A2(W15579), .ZN(W23880));
  NOR2X1 G10216 (.A1(W2388), .A2(W2784), .ZN(W4448));
  NOR2X1 G10217 (.A1(W24678), .A2(I914), .ZN(O3887));
  NOR2X1 G10218 (.A1(W1350), .A2(W415), .ZN(W4443));
  NOR2X1 G10219 (.A1(I50), .A2(W991), .ZN(W4442));
  NOR2X1 G10220 (.A1(W1733), .A2(I582), .ZN(W4409));
  NOR2X1 G10221 (.A1(W5036), .A2(I60), .ZN(O15660));
  NOR2X1 G10222 (.A1(I299), .A2(W1743), .ZN(W4439));
  NOR2X1 G10223 (.A1(W36517), .A2(W6830), .ZN(O15661));
  NOR2X1 G10224 (.A1(W23467), .A2(I1460), .ZN(W23885));
  NOR2X1 G10225 (.A1(W19447), .A2(W7573), .ZN(W46573));
  NOR2X1 G10226 (.A1(W10632), .A2(W39023), .ZN(O15663));
  NOR2X1 G10227 (.A1(I1053), .A2(W787), .ZN(W4433));
  NOR2X1 G10228 (.A1(I398), .A2(I1102), .ZN(W4382));
  NOR2X1 G10229 (.A1(W3861), .A2(W847), .ZN(W4390));
  NOR2X1 G10230 (.A1(W34230), .A2(W35600), .ZN(O15700));
  NOR2X1 G10231 (.A1(W12626), .A2(I1484), .ZN(W26819));
  NOR2X1 G10232 (.A1(W6437), .A2(W21479), .ZN(W23899));
  NOR2X1 G10233 (.A1(W3350), .A2(W3906), .ZN(W4386));
  NOR2X1 G10234 (.A1(W15236), .A2(W17821), .ZN(O2917));
  NOR2X1 G10235 (.A1(W3525), .A2(W2967), .ZN(W4384));
  NOR2X1 G10236 (.A1(W651), .A2(I828), .ZN(W4383));
  NOR2X1 G10237 (.A1(W726), .A2(W2783), .ZN(W4391));
  NOR2X1 G10238 (.A1(W1525), .A2(W2889), .ZN(W4381));
  NOR2X1 G10239 (.A1(W274), .A2(W22886), .ZN(O3883));
  NOR2X1 G10240 (.A1(W689), .A2(W4158), .ZN(W4379));
  NOR2X1 G10241 (.A1(W21046), .A2(W982), .ZN(O15704));
  NOR2X1 G10242 (.A1(I1358), .A2(W2248), .ZN(W4377));
  NOR2X1 G10243 (.A1(W45977), .A2(W33140), .ZN(O15706));
  NOR2X1 G10244 (.A1(W22562), .A2(W14098), .ZN(O15707));
  NOR2X1 G10245 (.A1(W27869), .A2(W43205), .ZN(O15693));
  NOR2X1 G10246 (.A1(W5270), .A2(W7486), .ZN(O15686));
  NOR2X1 G10247 (.A1(W867), .A2(W2067), .ZN(W23895));
  NOR2X1 G10248 (.A1(W20875), .A2(W7299), .ZN(O15689));
  NOR2X1 G10249 (.A1(I62), .A2(W4542), .ZN(W46605));
  NOR2X1 G10250 (.A1(W6070), .A2(W13586), .ZN(W46606));
  NOR2X1 G10251 (.A1(W2798), .A2(I1516), .ZN(W4403));
  NOR2X1 G10252 (.A1(W4224), .A2(W28004), .ZN(O15691));
  NOR2X1 G10253 (.A1(W20734), .A2(W12806), .ZN(W23897));
  NOR2X1 G10254 (.A1(W3058), .A2(W2015), .ZN(W4453));
  NOR2X1 G10255 (.A1(W45714), .A2(W27746), .ZN(O15694));
  NOR2X1 G10256 (.A1(W46212), .A2(W42521), .ZN(O15695));
  NOR2X1 G10257 (.A1(W15463), .A2(W21182), .ZN(O15697));
  NOR2X1 G10258 (.A1(W30147), .A2(W34195), .ZN(W46615));
  NOR2X1 G10259 (.A1(W233), .A2(W2005), .ZN(W4394));
  NOR2X1 G10260 (.A1(W36978), .A2(W23715), .ZN(O15699));
  NOR2X1 G10261 (.A1(W1996), .A2(I95), .ZN(W4392));
  NOR2X1 G10262 (.A1(W2689), .A2(W1836), .ZN(W4502));
  NOR2X1 G10263 (.A1(W13738), .A2(W24691), .ZN(W46511));
  NOR2X1 G10264 (.A1(W2337), .A2(W924), .ZN(W4509));
  NOR2X1 G10265 (.A1(W20700), .A2(W24363), .ZN(W26861));
  NOR2X1 G10266 (.A1(W18283), .A2(W7471), .ZN(W26860));
  NOR2X1 G10267 (.A1(W2822), .A2(W3819), .ZN(W4506));
  NOR2X1 G10268 (.A1(W284), .A2(W1262), .ZN(W4505));
  NOR2X1 G10269 (.A1(W14219), .A2(W8942), .ZN(O2904));
  NOR2X1 G10270 (.A1(I1694), .A2(I1415), .ZN(W4503));
  NOR2X1 G10271 (.A1(W10064), .A2(W34482), .ZN(O15611));
  NOR2X1 G10272 (.A1(W38729), .A2(W27814), .ZN(O15615));
  NOR2X1 G10273 (.A1(W21217), .A2(W8574), .ZN(W26859));
  NOR2X1 G10274 (.A1(W3448), .A2(W13570), .ZN(O3894));
  NOR2X1 G10275 (.A1(W23490), .A2(W6543), .ZN(O3893));
  NOR2X1 G10276 (.A1(I1477), .A2(W3400), .ZN(W4497));
  NOR2X1 G10277 (.A1(W24514), .A2(W17192), .ZN(W26853));
  NOR2X1 G10278 (.A1(W38087), .A2(W5522), .ZN(O15623));
  NOR2X1 G10279 (.A1(W531), .A2(I400), .ZN(W4494));
  NOR2X1 G10280 (.A1(W3217), .A2(I542), .ZN(W4520));
  NOR2X1 G10281 (.A1(W23072), .A2(W25901), .ZN(O3896));
  NOR2X1 G10282 (.A1(W25943), .A2(W5507), .ZN(O15599));
  NOR2X1 G10283 (.A1(W386), .A2(W11285), .ZN(O2900));
  NOR2X1 G10284 (.A1(I626), .A2(W4070), .ZN(W4527));
  NOR2X1 G10285 (.A1(W35731), .A2(W38436), .ZN(O15602));
  NOR2X1 G10286 (.A1(W29452), .A2(W35182), .ZN(O15603));
  NOR2X1 G10287 (.A1(W17449), .A2(W18511), .ZN(W23853));
  NOR2X1 G10288 (.A1(W4233), .A2(W321), .ZN(W4522));
  NOR2X1 G10289 (.A1(W21763), .A2(W16301), .ZN(W26852));
  NOR2X1 G10290 (.A1(W13920), .A2(W23894), .ZN(W26862));
  NOR2X1 G10291 (.A1(W829), .A2(W4243), .ZN(W4517));
  NOR2X1 G10292 (.A1(W15604), .A2(W24114), .ZN(O15608));
  NOR2X1 G10293 (.A1(W1227), .A2(I1131), .ZN(W4515));
  NOR2X1 G10294 (.A1(W259), .A2(W584), .ZN(W4514));
  NOR2X1 G10295 (.A1(W2101), .A2(W2121), .ZN(W4513));
  NOR2X1 G10296 (.A1(W27219), .A2(W36470), .ZN(O15610));
  NOR2X1 G10297 (.A1(W42864), .A2(W40319), .ZN(O15645));
  NOR2X1 G10298 (.A1(W3408), .A2(W3974), .ZN(W4471));
  NOR2X1 G10299 (.A1(W118), .A2(I389), .ZN(W4470));
  NOR2X1 G10300 (.A1(W2103), .A2(I1660), .ZN(W4469));
  NOR2X1 G10301 (.A1(W5450), .A2(W4021), .ZN(W23873));
  NOR2X1 G10302 (.A1(W14841), .A2(W11978), .ZN(W26838));
  NOR2X1 G10303 (.A1(W1772), .A2(W969), .ZN(W4466));
  NOR2X1 G10304 (.A1(W1739), .A2(W2393), .ZN(W4464));
  NOR2X1 G10305 (.A1(W35), .A2(W25994), .ZN(O15644));
  NOR2X1 G10306 (.A1(W1022), .A2(W1905), .ZN(W4472));
  NOR2X1 G10307 (.A1(W2404), .A2(I1542), .ZN(W4461));
  NOR2X1 G10308 (.A1(W31967), .A2(W17025), .ZN(O15646));
  NOR2X1 G10309 (.A1(W34828), .A2(W27199), .ZN(O15647));
  NOR2X1 G10310 (.A1(W3136), .A2(W144), .ZN(W4458));
  NOR2X1 G10311 (.A1(W6671), .A2(W3586), .ZN(W23876));
  NOR2X1 G10312 (.A1(W19040), .A2(W7662), .ZN(W23877));
  NOR2X1 G10313 (.A1(W324), .A2(W3534), .ZN(W4454));
  NOR2X1 G10314 (.A1(W1710), .A2(W1128), .ZN(W4481));
  NOR2X1 G10315 (.A1(W1291), .A2(W571), .ZN(W4492));
  NOR2X1 G10316 (.A1(W15378), .A2(W8980), .ZN(W26848));
  NOR2X1 G10317 (.A1(W43462), .A2(W32530), .ZN(W46533));
  NOR2X1 G10318 (.A1(W24950), .A2(W4611), .ZN(W26847));
  NOR2X1 G10319 (.A1(W3223), .A2(W36965), .ZN(O15632));
  NOR2X1 G10320 (.A1(W2944), .A2(W1726), .ZN(W4484));
  NOR2X1 G10321 (.A1(W24136), .A2(W28689), .ZN(O15634));
  NOR2X1 G10322 (.A1(W2595), .A2(W1696), .ZN(W4482));
  NOR2X1 G10323 (.A1(W2485), .A2(W2565), .ZN(O2882));
  NOR2X1 G10324 (.A1(W17443), .A2(W17680), .ZN(O15637));
  NOR2X1 G10325 (.A1(W497), .A2(W157), .ZN(W4479));
  NOR2X1 G10326 (.A1(W13383), .A2(W16514), .ZN(O3890));
  NOR2X1 G10327 (.A1(W356), .A2(W20743), .ZN(O2912));
  NOR2X1 G10328 (.A1(W2250), .A2(I224), .ZN(W4475));
  NOR2X1 G10329 (.A1(W24578), .A2(W2711), .ZN(O15640));
  NOR2X1 G10330 (.A1(I1968), .A2(W2665), .ZN(W4473));
  NOR2X1 G10331 (.A1(W25316), .A2(W39053), .ZN(W46100));
  NOR2X1 G10332 (.A1(W22589), .A2(W20222), .ZN(O3956));
  NOR2X1 G10333 (.A1(W14300), .A2(W11810), .ZN(O15253));
  NOR2X1 G10334 (.A1(W6141), .A2(W13383), .ZN(W23720));
  NOR2X1 G10335 (.A1(W5597), .A2(W23439), .ZN(W23721));
  NOR2X1 G10336 (.A1(W977), .A2(W18728), .ZN(W46094));
  NOR2X1 G10337 (.A1(W3866), .A2(W421), .ZN(W4897));
  NOR2X1 G10338 (.A1(W25143), .A2(I1389), .ZN(O15256));
  NOR2X1 G10339 (.A1(W23453), .A2(W1796), .ZN(W26999));
  NOR2X1 G10340 (.A1(W3715), .A2(W20548), .ZN(W23718));
  NOR2X1 G10341 (.A1(W7828), .A2(W30202), .ZN(O15261));
  NOR2X1 G10342 (.A1(W1754), .A2(I71), .ZN(W4892));
  NOR2X1 G10343 (.A1(W9463), .A2(W45590), .ZN(W46102));
  NOR2X1 G10344 (.A1(W6004), .A2(W4995), .ZN(W23723));
  NOR2X1 G10345 (.A1(W1468), .A2(I934), .ZN(W4889));
  NOR2X1 G10346 (.A1(W35683), .A2(W36936), .ZN(W46107));
  NOR2X1 G10347 (.A1(W17830), .A2(W15199), .ZN(W23724));
  NOR2X1 G10348 (.A1(W6377), .A2(W5046), .ZN(O15267));
  NOR2X1 G10349 (.A1(I1124), .A2(W725), .ZN(W4911));
  NOR2X1 G10350 (.A1(W3660), .A2(I255), .ZN(W27012));
  NOR2X1 G10351 (.A1(I1564), .A2(W3249), .ZN(W4919));
  NOR2X1 G10352 (.A1(W23390), .A2(W7228), .ZN(O2856));
  NOR2X1 G10353 (.A1(W10794), .A2(W11629), .ZN(W27010));
  NOR2X1 G10354 (.A1(W15364), .A2(W4998), .ZN(O15238));
  NOR2X1 G10355 (.A1(W38050), .A2(W25130), .ZN(O15240));
  NOR2X1 G10356 (.A1(W5312), .A2(W39724), .ZN(W46074));
  NOR2X1 G10357 (.A1(W41190), .A2(W16284), .ZN(O15241));
  NOR2X1 G10358 (.A1(W25444), .A2(W18632), .ZN(O3955));
  NOR2X1 G10359 (.A1(W921), .A2(I1377), .ZN(W4910));
  NOR2X1 G10360 (.A1(W1931), .A2(I1473), .ZN(O3958));
  NOR2X1 G10361 (.A1(W8054), .A2(W10560), .ZN(W27005));
  NOR2X1 G10362 (.A1(W5691), .A2(W25546), .ZN(W27004));
  NOR2X1 G10363 (.A1(W17440), .A2(W35528), .ZN(W46082));
  NOR2X1 G10364 (.A1(W11662), .A2(W2950), .ZN(W23717));
  NOR2X1 G10365 (.A1(W943), .A2(W2725), .ZN(W4904));
  NOR2X1 G10366 (.A1(W2708), .A2(W1483), .ZN(W4859));
  NOR2X1 G10367 (.A1(W45953), .A2(W24055), .ZN(O15282));
  NOR2X1 G10368 (.A1(W19391), .A2(W22041), .ZN(W26994));
  NOR2X1 G10369 (.A1(W15160), .A2(I566), .ZN(W26993));
  NOR2X1 G10370 (.A1(W4121), .A2(W5024), .ZN(O15287));
  NOR2X1 G10371 (.A1(W1535), .A2(W3588), .ZN(W4863));
  NOR2X1 G10372 (.A1(W12614), .A2(W15175), .ZN(W23732));
  NOR2X1 G10373 (.A1(W30627), .A2(W24535), .ZN(O15289));
  NOR2X1 G10374 (.A1(W21965), .A2(W455), .ZN(O15290));
  NOR2X1 G10375 (.A1(W22069), .A2(W42752), .ZN(O15281));
  NOR2X1 G10376 (.A1(I444), .A2(I1764), .ZN(W4858));
  NOR2X1 G10377 (.A1(W16631), .A2(W18792), .ZN(W23733));
  NOR2X1 G10378 (.A1(W159), .A2(W18217), .ZN(O15292));
  NOR2X1 G10379 (.A1(W6065), .A2(W19030), .ZN(W26992));
  NOR2X1 G10380 (.A1(W15750), .A2(W45587), .ZN(O15294));
  NOR2X1 G10381 (.A1(W34428), .A2(W32686), .ZN(O15295));
  NOR2X1 G10382 (.A1(I923), .A2(W4392), .ZN(W4852));
  NOR2X1 G10383 (.A1(W4010), .A2(W487), .ZN(W4876));
  NOR2X1 G10384 (.A1(W27984), .A2(W10603), .ZN(O15269));
  NOR2X1 G10385 (.A1(W3368), .A2(W2171), .ZN(W4883));
  NOR2X1 G10386 (.A1(W8457), .A2(W3681), .ZN(W23726));
  NOR2X1 G10387 (.A1(W25696), .A2(W14), .ZN(O15271));
  NOR2X1 G10388 (.A1(W2208), .A2(I1455), .ZN(W4880));
  NOR2X1 G10389 (.A1(I1166), .A2(W878), .ZN(O15272));
  NOR2X1 G10390 (.A1(W36593), .A2(W38338), .ZN(O15273));
  NOR2X1 G10391 (.A1(W3862), .A2(I486), .ZN(W4877));
  NOR2X1 G10392 (.A1(W8054), .A2(W32081), .ZN(W46059));
  NOR2X1 G10393 (.A1(W19045), .A2(W23133), .ZN(O2860));
  NOR2X1 G10394 (.A1(W2461), .A2(W3946), .ZN(W4874));
  NOR2X1 G10395 (.A1(W904), .A2(W3622), .ZN(W4873));
  NOR2X1 G10396 (.A1(W10528), .A2(W16084), .ZN(O3953));
  NOR2X1 G10397 (.A1(W2204), .A2(W1611), .ZN(W4871));
  NOR2X1 G10398 (.A1(I1957), .A2(W78), .ZN(W4870));
  NOR2X1 G10399 (.A1(W10565), .A2(W22402), .ZN(W23729));
  NOR2X1 G10400 (.A1(W22287), .A2(W4875), .ZN(W45993));
  NOR2X1 G10401 (.A1(I615), .A2(W3146), .ZN(W4982));
  NOR2X1 G10402 (.A1(W20111), .A2(W9153), .ZN(W27036));
  NOR2X1 G10403 (.A1(I1881), .A2(W4420), .ZN(W4980));
  NOR2X1 G10404 (.A1(W21811), .A2(W18635), .ZN(O15165));
  NOR2X1 G10405 (.A1(W7725), .A2(W17046), .ZN(W23685));
  NOR2X1 G10406 (.A1(I750), .A2(I661), .ZN(W4977));
  NOR2X1 G10407 (.A1(I1609), .A2(W35090), .ZN(O15168));
  NOR2X1 G10408 (.A1(I1432), .A2(W21797), .ZN(O15170));
  NOR2X1 G10409 (.A1(W3466), .A2(W6137), .ZN(W27037));
  NOR2X1 G10410 (.A1(W8387), .A2(W16681), .ZN(W23687));
  NOR2X1 G10411 (.A1(W958), .A2(W14518), .ZN(W27034));
  NOR2X1 G10412 (.A1(W44864), .A2(W33916), .ZN(O15174));
  NOR2X1 G10413 (.A1(W3437), .A2(W328), .ZN(W23689));
  NOR2X1 G10414 (.A1(W35230), .A2(W5190), .ZN(O15178));
  NOR2X1 G10415 (.A1(W42790), .A2(W20091), .ZN(O15179));
  NOR2X1 G10416 (.A1(W19394), .A2(W31634), .ZN(O15182));
  NOR2X1 G10417 (.A1(W1350), .A2(W21171), .ZN(O3963));
  NOR2X1 G10418 (.A1(I1176), .A2(I1856), .ZN(O3966));
  NOR2X1 G10419 (.A1(W11214), .A2(W4746), .ZN(W45967));
  NOR2X1 G10420 (.A1(W2845), .A2(W2635), .ZN(W5001));
  NOR2X1 G10421 (.A1(W36754), .A2(W16223), .ZN(O15151));
  NOR2X1 G10422 (.A1(W34653), .A2(W43568), .ZN(W45971));
  NOR2X1 G10423 (.A1(I1523), .A2(W1487), .ZN(W4998));
  NOR2X1 G10424 (.A1(W42414), .A2(W40860), .ZN(O15154));
  NOR2X1 G10425 (.A1(W13518), .A2(W19534), .ZN(W27047));
  NOR2X1 G10426 (.A1(I684), .A2(W2049), .ZN(W4995));
  NOR2X1 G10427 (.A1(W14435), .A2(W19324), .ZN(O3962));
  NOR2X1 G10428 (.A1(W40582), .A2(W33686), .ZN(O15159));
  NOR2X1 G10429 (.A1(I903), .A2(I1445), .ZN(W4990));
  NOR2X1 G10430 (.A1(I86), .A2(W1492), .ZN(W4989));
  NOR2X1 G10431 (.A1(W3173), .A2(W1625), .ZN(W4988));
  NOR2X1 G10432 (.A1(W4775), .A2(W2174), .ZN(W4987));
  NOR2X1 G10433 (.A1(W8506), .A2(W31281), .ZN(O15160));
  NOR2X1 G10434 (.A1(W45470), .A2(W15118), .ZN(W45980));
  NOR2X1 G10435 (.A1(I456), .A2(W2163), .ZN(W4930));
  NOR2X1 G10436 (.A1(W11089), .A2(W6297), .ZN(O2853));
  NOR2X1 G10437 (.A1(W4458), .A2(W4020), .ZN(W4940));
  NOR2X1 G10438 (.A1(W13077), .A2(W8489), .ZN(W27020));
  NOR2X1 G10439 (.A1(W968), .A2(W31), .ZN(W4937));
  NOR2X1 G10440 (.A1(W2586), .A2(I1640), .ZN(W4934));
  NOR2X1 G10441 (.A1(I896), .A2(W1528), .ZN(W4933));
  NOR2X1 G10442 (.A1(W21857), .A2(W23551), .ZN(W27016));
  NOR2X1 G10443 (.A1(W10322), .A2(W14654), .ZN(W23707));
  NOR2X1 G10444 (.A1(W16845), .A2(W1775), .ZN(W23700));
  NOR2X1 G10445 (.A1(W4312), .A2(W2389), .ZN(W4929));
  NOR2X1 G10446 (.A1(I1732), .A2(W2764), .ZN(W4928));
  NOR2X1 G10447 (.A1(W32694), .A2(W18193), .ZN(W46052));
  NOR2X1 G10448 (.A1(W1174), .A2(I753), .ZN(W4926));
  NOR2X1 G10449 (.A1(W22241), .A2(W19028), .ZN(W27014));
  NOR2X1 G10450 (.A1(W6359), .A2(W11992), .ZN(O15224));
  NOR2X1 G10451 (.A1(W35835), .A2(W41938), .ZN(O15225));
  NOR2X1 G10452 (.A1(W2521), .A2(W15605), .ZN(W27023));
  NOR2X1 G10453 (.A1(W36413), .A2(W23114), .ZN(O15187));
  NOR2X1 G10454 (.A1(W14542), .A2(W31394), .ZN(O15190));
  NOR2X1 G10455 (.A1(W32929), .A2(W19187), .ZN(O15192));
  NOR2X1 G10456 (.A1(W19942), .A2(W13629), .ZN(W23696));
  NOR2X1 G10457 (.A1(W70), .A2(W5), .ZN(W4955));
  NOR2X1 G10458 (.A1(W38382), .A2(W27954), .ZN(O15200));
  NOR2X1 G10459 (.A1(W14176), .A2(W1239), .ZN(W23697));
  NOR2X1 G10460 (.A1(I1632), .A2(W11234), .ZN(O15202));
  NOR2X1 G10461 (.A1(W19873), .A2(I1497), .ZN(W23735));
  NOR2X1 G10462 (.A1(W3126), .A2(W2488), .ZN(W4949));
  NOR2X1 G10463 (.A1(W5287), .A2(W19855), .ZN(O15206));
  NOR2X1 G10464 (.A1(W25184), .A2(W20035), .ZN(W46037));
  NOR2X1 G10465 (.A1(I1113), .A2(I290), .ZN(W4946));
  NOR2X1 G10466 (.A1(W16139), .A2(W45236), .ZN(O15208));
  NOR2X1 G10467 (.A1(W10717), .A2(W8221), .ZN(O15209));
  NOR2X1 G10468 (.A1(W3085), .A2(W25815), .ZN(O15210));
  NOR2X1 G10469 (.A1(W3397), .A2(W2489), .ZN(W4736));
  NOR2X1 G10470 (.A1(W3596), .A2(I1859), .ZN(W4744));
  NOR2X1 G10471 (.A1(W22465), .A2(W14779), .ZN(O15413));
  NOR2X1 G10472 (.A1(W3327), .A2(W849), .ZN(W4742));
  NOR2X1 G10473 (.A1(W12398), .A2(W18547), .ZN(O15415));
  NOR2X1 G10474 (.A1(W8894), .A2(W11987), .ZN(O3933));
  NOR2X1 G10475 (.A1(W19189), .A2(W31513), .ZN(O15418));
  NOR2X1 G10476 (.A1(W2890), .A2(W4373), .ZN(W4738));
  NOR2X1 G10477 (.A1(W12751), .A2(W22600), .ZN(W23779));
  NOR2X1 G10478 (.A1(W27619), .A2(W23128), .ZN(O15412));
  NOR2X1 G10479 (.A1(W9718), .A2(W26921), .ZN(O15420));
  NOR2X1 G10480 (.A1(I1398), .A2(W26138), .ZN(O3932));
  NOR2X1 G10481 (.A1(W10184), .A2(W22620), .ZN(O3931));
  NOR2X1 G10482 (.A1(W1543), .A2(W505), .ZN(W4732));
  NOR2X1 G10483 (.A1(W12680), .A2(W29378), .ZN(O15424));
  NOR2X1 G10484 (.A1(W32445), .A2(W5298), .ZN(O15425));
  NOR2X1 G10485 (.A1(W110), .A2(W3148), .ZN(O3930));
  NOR2X1 G10486 (.A1(I988), .A2(W3750), .ZN(W4728));
  NOR2X1 G10487 (.A1(W12775), .A2(W4019), .ZN(W26944));
  NOR2X1 G10488 (.A1(W4543), .A2(W38474), .ZN(O15391));
  NOR2X1 G10489 (.A1(W38519), .A2(W35452), .ZN(O15392));
  NOR2X1 G10490 (.A1(W2246), .A2(W1651), .ZN(W4762));
  NOR2X1 G10491 (.A1(W10781), .A2(W31987), .ZN(O15393));
  NOR2X1 G10492 (.A1(W3855), .A2(W9380), .ZN(O3938));
  NOR2X1 G10493 (.A1(W2739), .A2(W1944), .ZN(W4759));
  NOR2X1 G10494 (.A1(W26469), .A2(W1595), .ZN(O15397));
  NOR2X1 G10495 (.A1(W4974), .A2(W8298), .ZN(W26947));
  NOR2X1 G10496 (.A1(W4903), .A2(W12846), .ZN(W23783));
  NOR2X1 G10497 (.A1(W4745), .A2(I506), .ZN(O2875));
  NOR2X1 G10498 (.A1(W1515), .A2(W3851), .ZN(W4752));
  NOR2X1 G10499 (.A1(W10078), .A2(W23497), .ZN(O3935));
  NOR2X1 G10500 (.A1(W14154), .A2(W16785), .ZN(O2876));
  NOR2X1 G10501 (.A1(W17510), .A2(I7), .ZN(O15410));
  NOR2X1 G10502 (.A1(W2866), .A2(I340), .ZN(O63));
  NOR2X1 G10503 (.A1(W4182), .A2(I686), .ZN(W4746));
  NOR2X1 G10504 (.A1(W1721), .A2(I586), .ZN(W4697));
  NOR2X1 G10505 (.A1(W26616), .A2(W8840), .ZN(O3922));
  NOR2X1 G10506 (.A1(W20215), .A2(W41219), .ZN(O15459));
  NOR2X1 G10507 (.A1(W21530), .A2(W18541), .ZN(O15460));
  NOR2X1 G10508 (.A1(I1981), .A2(W616), .ZN(W4703));
  NOR2X1 G10509 (.A1(W10574), .A2(W11485), .ZN(O3921));
  NOR2X1 G10510 (.A1(W188), .A2(W3192), .ZN(W4700));
  NOR2X1 G10511 (.A1(W454), .A2(I1633), .ZN(W4699));
  NOR2X1 G10512 (.A1(W4089), .A2(I1977), .ZN(W4698));
  NOR2X1 G10513 (.A1(I1794), .A2(W1218), .ZN(W4707));
  NOR2X1 G10514 (.A1(W27744), .A2(W35285), .ZN(O15463));
  NOR2X1 G10515 (.A1(W14030), .A2(W44384), .ZN(O15464));
  NOR2X1 G10516 (.A1(W27911), .A2(W44231), .ZN(O15465));
  NOR2X1 G10517 (.A1(W483), .A2(W17518), .ZN(O3920));
  NOR2X1 G10518 (.A1(W11875), .A2(W293), .ZN(O3919));
  NOR2X1 G10519 (.A1(W44590), .A2(W3615), .ZN(W46345));
  NOR2X1 G10520 (.A1(W37011), .A2(I162), .ZN(O15471));
  NOR2X1 G10521 (.A1(W3117), .A2(W2435), .ZN(W4716));
  NOR2X1 G10522 (.A1(W11503), .A2(W9881), .ZN(O3927));
  NOR2X1 G10523 (.A1(W23986), .A2(W13061), .ZN(O15437));
  NOR2X1 G10524 (.A1(W46124), .A2(W4235), .ZN(O15438));
  NOR2X1 G10525 (.A1(W388), .A2(W4102), .ZN(O62));
  NOR2X1 G10526 (.A1(W3135), .A2(W3745), .ZN(W4720));
  NOR2X1 G10527 (.A1(W10306), .A2(W7053), .ZN(O15440));
  NOR2X1 G10528 (.A1(W16411), .A2(W1634), .ZN(O15441));
  NOR2X1 G10529 (.A1(W40305), .A2(W9190), .ZN(O15443));
  NOR2X1 G10530 (.A1(I225), .A2(I137), .ZN(W4765));
  NOR2X1 G10531 (.A1(W29318), .A2(W27364), .ZN(O15448));
  NOR2X1 G10532 (.A1(W4961), .A2(W17635), .ZN(W26930));
  NOR2X1 G10533 (.A1(I960), .A2(W3598), .ZN(W4713));
  NOR2X1 G10534 (.A1(W577), .A2(W41683), .ZN(O15452));
  NOR2X1 G10535 (.A1(W4293), .A2(W14102), .ZN(W26929));
  NOR2X1 G10536 (.A1(W629), .A2(W16234), .ZN(W46329));
  NOR2X1 G10537 (.A1(W16256), .A2(W7785), .ZN(O15456));
  NOR2X1 G10538 (.A1(W28997), .A2(W4554), .ZN(O15343));
  NOR2X1 G10539 (.A1(W1564), .A2(W17480), .ZN(O15325));
  NOR2X1 G10540 (.A1(W1327), .A2(W24277), .ZN(W26977));
  NOR2X1 G10541 (.A1(W3385), .A2(W18846), .ZN(O15332));
  NOR2X1 G10542 (.A1(W1023), .A2(I1572), .ZN(W4825));
  NOR2X1 G10543 (.A1(W12376), .A2(I790), .ZN(W23746));
  NOR2X1 G10544 (.A1(W7418), .A2(W11558), .ZN(O2867));
  NOR2X1 G10545 (.A1(I1963), .A2(W3003), .ZN(W4819));
  NOR2X1 G10546 (.A1(W15846), .A2(W24657), .ZN(O15342));
  NOR2X1 G10547 (.A1(W5335), .A2(W1750), .ZN(O15322));
  NOR2X1 G10548 (.A1(W40913), .A2(W40256), .ZN(O15344));
  NOR2X1 G10549 (.A1(W9820), .A2(W44414), .ZN(O15346));
  NOR2X1 G10550 (.A1(W22835), .A2(W3227), .ZN(W26971));
  NOR2X1 G10551 (.A1(W39271), .A2(W38614), .ZN(O15349));
  NOR2X1 G10552 (.A1(W19463), .A2(W26933), .ZN(W26970));
  NOR2X1 G10553 (.A1(W1310), .A2(W2563), .ZN(W4810));
  NOR2X1 G10554 (.A1(I1894), .A2(W4477), .ZN(W4809));
  NOR2X1 G10555 (.A1(W3682), .A2(W3905), .ZN(W4807));
  NOR2X1 G10556 (.A1(W14878), .A2(W34142), .ZN(O15310));
  NOR2X1 G10557 (.A1(W25725), .A2(W39889), .ZN(O15298));
  NOR2X1 G10558 (.A1(W13917), .A2(W3569), .ZN(O15299));
  NOR2X1 G10559 (.A1(W1416), .A2(W4107), .ZN(W4846));
  NOR2X1 G10560 (.A1(W1215), .A2(W18482), .ZN(O15302));
  NOR2X1 G10561 (.A1(W21037), .A2(W5334), .ZN(W23738));
  NOR2X1 G10562 (.A1(W16572), .A2(W17434), .ZN(O3950));
  NOR2X1 G10563 (.A1(W3521), .A2(W3341), .ZN(W4841));
  NOR2X1 G10564 (.A1(W10632), .A2(W17863), .ZN(O15309));
  NOR2X1 G10565 (.A1(W1904), .A2(W2681), .ZN(W4806));
  NOR2X1 G10566 (.A1(W4206), .A2(I842), .ZN(W4838));
  NOR2X1 G10567 (.A1(W22138), .A2(W19873), .ZN(O2864));
  NOR2X1 G10568 (.A1(W532), .A2(W89), .ZN(W4835));
  NOR2X1 G10569 (.A1(W4190), .A2(W1539), .ZN(W4834));
  NOR2X1 G10570 (.A1(W36255), .A2(W18027), .ZN(O15315));
  NOR2X1 G10571 (.A1(W4759), .A2(W520), .ZN(W4832));
  NOR2X1 G10572 (.A1(W26898), .A2(W7925), .ZN(W26980));
  NOR2X1 G10573 (.A1(W4310), .A2(W1003), .ZN(W4773));
  NOR2X1 G10574 (.A1(W1117), .A2(W3741), .ZN(O15373));
  NOR2X1 G10575 (.A1(W324), .A2(W1128), .ZN(W4784));
  NOR2X1 G10576 (.A1(W12171), .A2(W1107), .ZN(W23762));
  NOR2X1 G10577 (.A1(W3696), .A2(W42382), .ZN(O15375));
  NOR2X1 G10578 (.A1(W32406), .A2(W7839), .ZN(W46242));
  NOR2X1 G10579 (.A1(W28721), .A2(W8845), .ZN(O15377));
  NOR2X1 G10580 (.A1(W18697), .A2(W72), .ZN(O15379));
  NOR2X1 G10581 (.A1(W5864), .A2(W4954), .ZN(O15382));
  NOR2X1 G10582 (.A1(W3471), .A2(W2621), .ZN(W4786));
  NOR2X1 G10583 (.A1(W21567), .A2(W16291), .ZN(W26952));
  NOR2X1 G10584 (.A1(W254), .A2(I417), .ZN(W4771));
  NOR2X1 G10585 (.A1(I481), .A2(W653), .ZN(W4770));
  NOR2X1 G10586 (.A1(W5199), .A2(W44185), .ZN(O15384));
  NOR2X1 G10587 (.A1(W20999), .A2(W16327), .ZN(O3939));
  NOR2X1 G10588 (.A1(W11458), .A2(W12245), .ZN(O15388));
  NOR2X1 G10589 (.A1(W14049), .A2(W26068), .ZN(O15389));
  NOR2X1 G10590 (.A1(W25526), .A2(W28810), .ZN(W46227));
  NOR2X1 G10591 (.A1(W10653), .A2(W23959), .ZN(W46210));
  NOR2X1 G10592 (.A1(W14402), .A2(W38748), .ZN(W46212));
  NOR2X1 G10593 (.A1(W21512), .A2(W13583), .ZN(O3945));
  NOR2X1 G10594 (.A1(W42976), .A2(I641), .ZN(O15357));
  NOR2X1 G10595 (.A1(W17397), .A2(W4924), .ZN(W23756));
  NOR2X1 G10596 (.A1(I1096), .A2(W6802), .ZN(O2868));
  NOR2X1 G10597 (.A1(W13123), .A2(W3614), .ZN(W46219));
  NOR2X1 G10598 (.A1(W24949), .A2(W10583), .ZN(W26964));
  NOR2X1 G10599 (.A1(W43732), .A2(W10640), .ZN(O15708));
  NOR2X1 G10600 (.A1(W4725), .A2(W450), .ZN(W4794));
  NOR2X1 G10601 (.A1(W28868), .A2(W39767), .ZN(O15366));
  NOR2X1 G10602 (.A1(W3009), .A2(I1860), .ZN(W4792));
  NOR2X1 G10603 (.A1(W7340), .A2(W29814), .ZN(W46229));
  NOR2X1 G10604 (.A1(W7337), .A2(W40577), .ZN(O15367));
  NOR2X1 G10605 (.A1(W16364), .A2(W24006), .ZN(O15368));
  NOR2X1 G10606 (.A1(W3617), .A2(W101), .ZN(W4788));
  NOR2X1 G10607 (.A1(W8328), .A2(W14489), .ZN(W24052));
  NOR2X1 G10608 (.A1(W21288), .A2(W24803), .ZN(O3834));
  NOR2X1 G10609 (.A1(W876), .A2(W3065), .ZN(W3965));
  NOR2X1 G10610 (.A1(W3141), .A2(W27002), .ZN(O16025));
  NOR2X1 G10611 (.A1(W30495), .A2(W3890), .ZN(W47007));
  NOR2X1 G10612 (.A1(W20603), .A2(W6435), .ZN(O3833));
  NOR2X1 G10613 (.A1(W34642), .A2(W15942), .ZN(O16029));
  NOR2X1 G10614 (.A1(I1296), .A2(W577), .ZN(W3960));
  NOR2X1 G10615 (.A1(W16709), .A2(W9156), .ZN(W24051));
  NOR2X1 G10616 (.A1(W2558), .A2(W9108), .ZN(W26686));
  NOR2X1 G10617 (.A1(W2312), .A2(W884), .ZN(W3957));
  NOR2X1 G10618 (.A1(W20694), .A2(W19232), .ZN(W24053));
  NOR2X1 G10619 (.A1(W27558), .A2(W25473), .ZN(O16037));
  NOR2X1 G10620 (.A1(I54), .A2(I86), .ZN(W3954));
  NOR2X1 G10621 (.A1(W29370), .A2(W44375), .ZN(O16038));
  NOR2X1 G10622 (.A1(W512), .A2(W1320), .ZN(W3951));
  NOR2X1 G10623 (.A1(W2020), .A2(W3433), .ZN(W3949));
  NOR2X1 G10624 (.A1(W2050), .A2(W1749), .ZN(W3948));
  NOR2X1 G10625 (.A1(W29500), .A2(W12806), .ZN(O16018));
  NOR2X1 G10626 (.A1(W24315), .A2(W17860), .ZN(W26693));
  NOR2X1 G10627 (.A1(W14666), .A2(W22149), .ZN(W26691));
  NOR2X1 G10628 (.A1(W20175), .A2(W23222), .ZN(O2957));
  NOR2X1 G10629 (.A1(W1218), .A2(I1960), .ZN(W3981));
  NOR2X1 G10630 (.A1(W30742), .A2(W34687), .ZN(O16013));
  NOR2X1 G10631 (.A1(W32481), .A2(W22397), .ZN(O16014));
  NOR2X1 G10632 (.A1(W41190), .A2(W24742), .ZN(O16015));
  NOR2X1 G10633 (.A1(I521), .A2(I948), .ZN(W3977));
  NOR2X1 G10634 (.A1(W10170), .A2(W20704), .ZN(O2961));
  NOR2X1 G10635 (.A1(W25506), .A2(W5657), .ZN(O16019));
  NOR2X1 G10636 (.A1(W44751), .A2(W46817), .ZN(W46999));
  NOR2X1 G10637 (.A1(W10122), .A2(W2529), .ZN(W24045));
  NOR2X1 G10638 (.A1(W20159), .A2(W9685), .ZN(W26687));
  NOR2X1 G10639 (.A1(W14150), .A2(W42846), .ZN(O16023));
  NOR2X1 G10640 (.A1(I1659), .A2(I668), .ZN(W3969));
  NOR2X1 G10641 (.A1(I1128), .A2(W2055), .ZN(W3968));
  NOR2X1 G10642 (.A1(I11), .A2(W765), .ZN(W3920));
  NOR2X1 G10643 (.A1(I1679), .A2(W1842), .ZN(W3928));
  NOR2X1 G10644 (.A1(W1132), .A2(W2164), .ZN(W3927));
  NOR2X1 G10645 (.A1(W2653), .A2(W2872), .ZN(W3926));
  NOR2X1 G10646 (.A1(W14330), .A2(W15197), .ZN(O16055));
  NOR2X1 G10647 (.A1(I1104), .A2(I1597), .ZN(W3924));
  NOR2X1 G10648 (.A1(W3986), .A2(W16315), .ZN(W26675));
  NOR2X1 G10649 (.A1(W28369), .A2(W15301), .ZN(O16057));
  NOR2X1 G10650 (.A1(W32318), .A2(W26065), .ZN(O16058));
  NOR2X1 G10651 (.A1(W13081), .A2(W18554), .ZN(W24061));
  NOR2X1 G10652 (.A1(W23020), .A2(W21187), .ZN(W24063));
  NOR2X1 G10653 (.A1(W25775), .A2(W39719), .ZN(O16061));
  NOR2X1 G10654 (.A1(W3657), .A2(W1686), .ZN(W3917));
  NOR2X1 G10655 (.A1(W46102), .A2(W35330), .ZN(O16063));
  NOR2X1 G10656 (.A1(W2232), .A2(W2654), .ZN(W3914));
  NOR2X1 G10657 (.A1(W26629), .A2(W6316), .ZN(O16067));
  NOR2X1 G10658 (.A1(W65), .A2(I422), .ZN(W3912));
  NOR2X1 G10659 (.A1(W46894), .A2(W3670), .ZN(O16070));
  NOR2X1 G10660 (.A1(W11944), .A2(W23191), .ZN(W24058));
  NOR2X1 G10661 (.A1(W421), .A2(I1776), .ZN(W3946));
  NOR2X1 G10662 (.A1(I697), .A2(W172), .ZN(W3945));
  NOR2X1 G10663 (.A1(W9076), .A2(I1909), .ZN(O16044));
  NOR2X1 G10664 (.A1(W24598), .A2(W30955), .ZN(O16045));
  NOR2X1 G10665 (.A1(W19213), .A2(I716), .ZN(O2962));
  NOR2X1 G10666 (.A1(W16756), .A2(W20620), .ZN(O16047));
  NOR2X1 G10667 (.A1(W37472), .A2(W38276), .ZN(O16048));
  NOR2X1 G10668 (.A1(I44), .A2(W883), .ZN(W3939));
  NOR2X1 G10669 (.A1(W13785), .A2(W3017), .ZN(W24038));
  NOR2X1 G10670 (.A1(I1954), .A2(W682), .ZN(W3937));
  NOR2X1 G10671 (.A1(W3250), .A2(W3281), .ZN(W3936));
  NOR2X1 G10672 (.A1(W2449), .A2(W21855), .ZN(O3830));
  NOR2X1 G10673 (.A1(I1377), .A2(W505), .ZN(W3934));
  NOR2X1 G10674 (.A1(W32781), .A2(W12756), .ZN(O16051));
  NOR2X1 G10675 (.A1(W29058), .A2(W24174), .ZN(O16052));
  NOR2X1 G10676 (.A1(W409), .A2(W1839), .ZN(W3930));
  NOR2X1 G10677 (.A1(W11482), .A2(W14863), .ZN(O15962));
  NOR2X1 G10678 (.A1(W38341), .A2(W36886), .ZN(O15955));
  NOR2X1 G10679 (.A1(W3181), .A2(W666), .ZN(W4044));
  NOR2X1 G10680 (.A1(I818), .A2(W6332), .ZN(O3845));
  NOR2X1 G10681 (.A1(W2914), .A2(W1793), .ZN(W4042));
  NOR2X1 G10682 (.A1(W33529), .A2(W44656), .ZN(W46928));
  NOR2X1 G10683 (.A1(W10835), .A2(W550), .ZN(W24020));
  NOR2X1 G10684 (.A1(W23320), .A2(W18910), .ZN(O2949));
  NOR2X1 G10685 (.A1(W43683), .A2(W21793), .ZN(W46931));
  NOR2X1 G10686 (.A1(W12955), .A2(W9912), .ZN(W24016));
  NOR2X1 G10687 (.A1(W3968), .A2(W2373), .ZN(W4035));
  NOR2X1 G10688 (.A1(W2211), .A2(W2855), .ZN(W4034));
  NOR2X1 G10689 (.A1(W3988), .A2(W37487), .ZN(O15963));
  NOR2X1 G10690 (.A1(W8125), .A2(W2972), .ZN(O15964));
  NOR2X1 G10691 (.A1(W374), .A2(W139), .ZN(W4031));
  NOR2X1 G10692 (.A1(W8906), .A2(W18723), .ZN(O2950));
  NOR2X1 G10693 (.A1(W35146), .A2(W25892), .ZN(O15967));
  NOR2X1 G10694 (.A1(W25113), .A2(W22470), .ZN(W26716));
  NOR2X1 G10695 (.A1(W3899), .A2(W3126), .ZN(W4057));
  NOR2X1 G10696 (.A1(W1639), .A2(W2016), .ZN(W4065));
  NOR2X1 G10697 (.A1(W42786), .A2(W34114), .ZN(O15940));
  NOR2X1 G10698 (.A1(I19), .A2(W3636), .ZN(O51));
  NOR2X1 G10699 (.A1(W6666), .A2(W22101), .ZN(W24008));
  NOR2X1 G10700 (.A1(W25156), .A2(W724), .ZN(O15942));
  NOR2X1 G10701 (.A1(W12582), .A2(W1020), .ZN(W24009));
  NOR2X1 G10702 (.A1(W8142), .A2(W2529), .ZN(O15944));
  NOR2X1 G10703 (.A1(W41196), .A2(W28074), .ZN(W46915));
  NOR2X1 G10704 (.A1(W4049), .A2(W20639), .ZN(W26713));
  NOR2X1 G10705 (.A1(W2945), .A2(W602), .ZN(W4056));
  NOR2X1 G10706 (.A1(W3035), .A2(I1265), .ZN(W4055));
  NOR2X1 G10707 (.A1(W23208), .A2(W14030), .ZN(W24011));
  NOR2X1 G10708 (.A1(W19636), .A2(W13740), .ZN(W24012));
  NOR2X1 G10709 (.A1(W4229), .A2(W8983), .ZN(O2948));
  NOR2X1 G10710 (.A1(W17138), .A2(W3390), .ZN(W24014));
  NOR2X1 G10711 (.A1(I198), .A2(W2091), .ZN(W4048));
  NOR2X1 G10712 (.A1(W878), .A2(W3146), .ZN(W3997));
  NOR2X1 G10713 (.A1(W9639), .A2(W21152), .ZN(O15991));
  NOR2X1 G10714 (.A1(W24722), .A2(W19292), .ZN(W26702));
  NOR2X1 G10715 (.A1(W12685), .A2(W9137), .ZN(W46969));
  NOR2X1 G10716 (.A1(W1771), .A2(I1068), .ZN(W4003));
  NOR2X1 G10717 (.A1(W6048), .A2(W23733), .ZN(W24033));
  NOR2X1 G10718 (.A1(W33868), .A2(W41374), .ZN(W46974));
  NOR2X1 G10719 (.A1(W2139), .A2(W3787), .ZN(W3999));
  NOR2X1 G10720 (.A1(W22160), .A2(W19042), .ZN(W26699));
  NOR2X1 G10721 (.A1(W12139), .A2(W19336), .ZN(W26705));
  NOR2X1 G10722 (.A1(W4533), .A2(W14114), .ZN(W24035));
  NOR2X1 G10723 (.A1(W10223), .A2(W40693), .ZN(O16001));
  NOR2X1 G10724 (.A1(W3836), .A2(W1781), .ZN(W3994));
  NOR2X1 G10725 (.A1(W811), .A2(W1769), .ZN(W3992));
  NOR2X1 G10726 (.A1(W461), .A2(W2818), .ZN(W26696));
  NOR2X1 G10727 (.A1(I1236), .A2(W1715), .ZN(W3990));
  NOR2X1 G10728 (.A1(W1835), .A2(I520), .ZN(W3989));
  NOR2X1 G10729 (.A1(W6476), .A2(W29881), .ZN(O15978));
  NOR2X1 G10730 (.A1(W1682), .A2(W546), .ZN(W4025));
  NOR2X1 G10731 (.A1(W34145), .A2(W32903), .ZN(O15973));
  NOR2X1 G10732 (.A1(W2800), .A2(W2713), .ZN(W4023));
  NOR2X1 G10733 (.A1(W860), .A2(W6133), .ZN(O3843));
  NOR2X1 G10734 (.A1(W2745), .A2(W35146), .ZN(O15976));
  NOR2X1 G10735 (.A1(I498), .A2(W32171), .ZN(W46948));
  NOR2X1 G10736 (.A1(W40114), .A2(W17550), .ZN(O15977));
  NOR2X1 G10737 (.A1(W3183), .A2(W972), .ZN(W4018));
  NOR2X1 G10738 (.A1(W9766), .A2(W14258), .ZN(W24066));
  NOR2X1 G10739 (.A1(I416), .A2(W2498), .ZN(W4016));
  NOR2X1 G10740 (.A1(W34625), .A2(W45387), .ZN(W46951));
  NOR2X1 G10741 (.A1(I1984), .A2(W243), .ZN(W4014));
  NOR2X1 G10742 (.A1(W24215), .A2(W6057), .ZN(O3842));
  NOR2X1 G10743 (.A1(W27621), .A2(W24183), .ZN(O15984));
  NOR2X1 G10744 (.A1(W1817), .A2(W23375), .ZN(O15986));
  NOR2X1 G10745 (.A1(I1619), .A2(W681), .ZN(W4008));
  NOR2X1 G10746 (.A1(W15427), .A2(W14872), .ZN(W24097));
  NOR2X1 G10747 (.A1(W35227), .A2(W31933), .ZN(W47158));
  NOR2X1 G10748 (.A1(W23948), .A2(W5466), .ZN(O16161));
  NOR2X1 G10749 (.A1(W25212), .A2(W11427), .ZN(O16162));
  NOR2X1 G10750 (.A1(W4860), .A2(W36572), .ZN(O16163));
  NOR2X1 G10751 (.A1(W2373), .A2(W2113), .ZN(W3811));
  NOR2X1 G10752 (.A1(W11195), .A2(W22415), .ZN(O16167));
  NOR2X1 G10753 (.A1(W197), .A2(I1687), .ZN(W3806));
  NOR2X1 G10754 (.A1(W8487), .A2(W37960), .ZN(O16169));
  NOR2X1 G10755 (.A1(W1529), .A2(I1847), .ZN(W3816));
  NOR2X1 G10756 (.A1(I146), .A2(W10521), .ZN(O16171));
  NOR2X1 G10757 (.A1(W16029), .A2(W35867), .ZN(O16174));
  NOR2X1 G10758 (.A1(W2363), .A2(W142), .ZN(W3800));
  NOR2X1 G10759 (.A1(W30), .A2(W1275), .ZN(W3798));
  NOR2X1 G10760 (.A1(W1411), .A2(I1381), .ZN(W3797));
  NOR2X1 G10761 (.A1(I1526), .A2(W3129), .ZN(W3796));
  NOR2X1 G10762 (.A1(W4941), .A2(W3737), .ZN(O2970));
  NOR2X1 G10763 (.A1(W32179), .A2(W10375), .ZN(O16177));
  NOR2X1 G10764 (.A1(W3220), .A2(I1336), .ZN(W3826));
  NOR2X1 G10765 (.A1(W2403), .A2(I1410), .ZN(W3834));
  NOR2X1 G10766 (.A1(W23108), .A2(W9830), .ZN(W24087));
  NOR2X1 G10767 (.A1(W20976), .A2(W39514), .ZN(O16136));
  NOR2X1 G10768 (.A1(W12838), .A2(I56), .ZN(O3818));
  NOR2X1 G10769 (.A1(W39144), .A2(W18069), .ZN(O16142));
  NOR2X1 G10770 (.A1(W34885), .A2(W18478), .ZN(O16146));
  NOR2X1 G10771 (.A1(W864), .A2(W3490), .ZN(W3828));
  NOR2X1 G10772 (.A1(W24587), .A2(W19760), .ZN(O16148));
  NOR2X1 G10773 (.A1(W2386), .A2(W236), .ZN(W3793));
  NOR2X1 G10774 (.A1(W31132), .A2(W18441), .ZN(O16150));
  NOR2X1 G10775 (.A1(W26563), .A2(W8095), .ZN(W26648));
  NOR2X1 G10776 (.A1(W1938), .A2(I24), .ZN(W3823));
  NOR2X1 G10777 (.A1(W9408), .A2(W23993), .ZN(W24090));
  NOR2X1 G10778 (.A1(W1636), .A2(W2301), .ZN(W3821));
  NOR2X1 G10779 (.A1(W21266), .A2(W13666), .ZN(W26647));
  NOR2X1 G10780 (.A1(W20303), .A2(W38694), .ZN(O16160));
  NOR2X1 G10781 (.A1(W19187), .A2(W13144), .ZN(W24110));
  NOR2X1 G10782 (.A1(I902), .A2(W20109), .ZN(O2973));
  NOR2X1 G10783 (.A1(W44296), .A2(W39880), .ZN(O16192));
  NOR2X1 G10784 (.A1(W18845), .A2(W21711), .ZN(O16194));
  NOR2X1 G10785 (.A1(W3754), .A2(W6040), .ZN(O16198));
  NOR2X1 G10786 (.A1(W31265), .A2(W42056), .ZN(O16199));
  NOR2X1 G10787 (.A1(W1669), .A2(I1585), .ZN(W3768));
  NOR2X1 G10788 (.A1(W5081), .A2(W5799), .ZN(W24108));
  NOR2X1 G10789 (.A1(W24920), .A2(W10391), .ZN(W26632));
  NOR2X1 G10790 (.A1(I1395), .A2(I930), .ZN(W3776));
  NOR2X1 G10791 (.A1(W31307), .A2(W7085), .ZN(O16204));
  NOR2X1 G10792 (.A1(W40111), .A2(W41432), .ZN(O16205));
  NOR2X1 G10793 (.A1(W24341), .A2(W35036), .ZN(O16206));
  NOR2X1 G10794 (.A1(W989), .A2(W28330), .ZN(O16208));
  NOR2X1 G10795 (.A1(I1065), .A2(W4149), .ZN(O16209));
  NOR2X1 G10796 (.A1(W1037), .A2(W917), .ZN(W3759));
  NOR2X1 G10797 (.A1(W1581), .A2(W2794), .ZN(O16210));
  NOR2X1 G10798 (.A1(W17696), .A2(W20409), .ZN(W26636));
  NOR2X1 G10799 (.A1(W2110), .A2(W3731), .ZN(W3792));
  NOR2X1 G10800 (.A1(W22206), .A2(W5669), .ZN(W24101));
  NOR2X1 G10801 (.A1(W40023), .A2(W12869), .ZN(O16180));
  NOR2X1 G10802 (.A1(I677), .A2(W2155), .ZN(W3789));
  NOR2X1 G10803 (.A1(W1466), .A2(W1018), .ZN(W3788));
  NOR2X1 G10804 (.A1(W1922), .A2(W18404), .ZN(W24102));
  NOR2X1 G10805 (.A1(W12066), .A2(I1382), .ZN(O16181));
  NOR2X1 G10806 (.A1(W2484), .A2(I1194), .ZN(W3785));
  NOR2X1 G10807 (.A1(W15056), .A2(W31978), .ZN(O16134));
  NOR2X1 G10808 (.A1(W2267), .A2(W2544), .ZN(W3783));
  NOR2X1 G10809 (.A1(W32249), .A2(W40257), .ZN(O16184));
  NOR2X1 G10810 (.A1(W25869), .A2(W42106), .ZN(W47185));
  NOR2X1 G10811 (.A1(W2380), .A2(W25343), .ZN(O16185));
  NOR2X1 G10812 (.A1(W18174), .A2(W21892), .ZN(W24104));
  NOR2X1 G10813 (.A1(W3650), .A2(I1388), .ZN(W3778));
  NOR2X1 G10814 (.A1(W2050), .A2(W3223), .ZN(W3777));
  NOR2X1 G10815 (.A1(W2042), .A2(W2991), .ZN(W3881));
  NOR2X1 G10816 (.A1(I1978), .A2(W2696), .ZN(W3889));
  NOR2X1 G10817 (.A1(W28360), .A2(W31914), .ZN(O16093));
  NOR2X1 G10818 (.A1(I1650), .A2(I1819), .ZN(W3887));
  NOR2X1 G10819 (.A1(W1731), .A2(W2937), .ZN(W3886));
  NOR2X1 G10820 (.A1(W3632), .A2(W2808), .ZN(W3885));
  NOR2X1 G10821 (.A1(W6592), .A2(W18612), .ZN(W24072));
  NOR2X1 G10822 (.A1(W18731), .A2(W6677), .ZN(O16095));
  NOR2X1 G10823 (.A1(W386), .A2(I614), .ZN(W3882));
  NOR2X1 G10824 (.A1(W1090), .A2(I840), .ZN(W3890));
  NOR2X1 G10825 (.A1(W24453), .A2(I575), .ZN(W26664));
  NOR2X1 G10826 (.A1(W1392), .A2(W3753), .ZN(W3878));
  NOR2X1 G10827 (.A1(W2662), .A2(I572), .ZN(W3877));
  NOR2X1 G10828 (.A1(W2075), .A2(W3191), .ZN(W3876));
  NOR2X1 G10829 (.A1(I764), .A2(W2364), .ZN(W3875));
  NOR2X1 G10830 (.A1(W19513), .A2(W8056), .ZN(W24075));
  NOR2X1 G10831 (.A1(W906), .A2(W3228), .ZN(W3873));
  NOR2X1 G10832 (.A1(W13900), .A2(W14223), .ZN(W26662));
  NOR2X1 G10833 (.A1(W34453), .A2(W41978), .ZN(O16080));
  NOR2X1 G10834 (.A1(W28397), .A2(W11106), .ZN(O16072));
  NOR2X1 G10835 (.A1(W2718), .A2(I597), .ZN(W3907));
  NOR2X1 G10836 (.A1(W13595), .A2(W17572), .ZN(W24067));
  NOR2X1 G10837 (.A1(W5913), .A2(W1155), .ZN(W26671));
  NOR2X1 G10838 (.A1(W44668), .A2(W40065), .ZN(O16077));
  NOR2X1 G10839 (.A1(W9870), .A2(W8011), .ZN(O3826));
  NOR2X1 G10840 (.A1(W3423), .A2(W17588), .ZN(W47066));
  NOR2X1 G10841 (.A1(W707), .A2(W24221), .ZN(W47067));
  NOR2X1 G10842 (.A1(W4835), .A2(W13381), .ZN(O3824));
  NOR2X1 G10843 (.A1(W23052), .A2(W25894), .ZN(O16081));
  NOR2X1 G10844 (.A1(W44645), .A2(W31816), .ZN(O16083));
  NOR2X1 G10845 (.A1(W5505), .A2(W4380), .ZN(O16084));
  NOR2X1 G10846 (.A1(I1400), .A2(W1836), .ZN(W3895));
  NOR2X1 G10847 (.A1(W32194), .A2(W39242), .ZN(W47074));
  NOR2X1 G10848 (.A1(I1167), .A2(W7926), .ZN(O16090));
  NOR2X1 G10849 (.A1(W22302), .A2(W23940), .ZN(O16091));
  NOR2X1 G10850 (.A1(W31585), .A2(W41532), .ZN(O16124));
  NOR2X1 G10851 (.A1(W2244), .A2(W3182), .ZN(W3852));
  NOR2X1 G10852 (.A1(W3351), .A2(W10366), .ZN(O3823));
  NOR2X1 G10853 (.A1(W1780), .A2(W3391), .ZN(W3850));
  NOR2X1 G10854 (.A1(W19199), .A2(W35570), .ZN(O16116));
  NOR2X1 G10855 (.A1(W10641), .A2(W11469), .ZN(O16117));
  NOR2X1 G10856 (.A1(I1812), .A2(W2749), .ZN(W24083));
  NOR2X1 G10857 (.A1(W10731), .A2(W25163), .ZN(O16122));
  NOR2X1 G10858 (.A1(W45121), .A2(W34317), .ZN(O16123));
  NOR2X1 G10859 (.A1(I686), .A2(W2112), .ZN(W3853));
  NOR2X1 G10860 (.A1(I1795), .A2(I1127), .ZN(W3843));
  NOR2X1 G10861 (.A1(W13541), .A2(W25409), .ZN(W26655));
  NOR2X1 G10862 (.A1(W20309), .A2(W36955), .ZN(W47126));
  NOR2X1 G10863 (.A1(W14199), .A2(W31725), .ZN(O16132));
  NOR2X1 G10864 (.A1(W1210), .A2(W1556), .ZN(W3838));
  NOR2X1 G10865 (.A1(W12333), .A2(W19536), .ZN(W24086));
  NOR2X1 G10866 (.A1(W2437), .A2(W420), .ZN(W3836));
  NOR2X1 G10867 (.A1(W1889), .A2(W3632), .ZN(W3861));
  NOR2X1 G10868 (.A1(W3724), .A2(I970), .ZN(W3870));
  NOR2X1 G10869 (.A1(W33365), .A2(W19258), .ZN(O16101));
  NOR2X1 G10870 (.A1(W12243), .A2(W8255), .ZN(W24078));
  NOR2X1 G10871 (.A1(W29326), .A2(W2391), .ZN(O16103));
  NOR2X1 G10872 (.A1(W2175), .A2(I1667), .ZN(W3866));
  NOR2X1 G10873 (.A1(W33586), .A2(W1191), .ZN(O16104));
  NOR2X1 G10874 (.A1(I1396), .A2(W1062), .ZN(W3864));
  NOR2X1 G10875 (.A1(W37637), .A2(W45837), .ZN(O16108));
  NOR2X1 G10876 (.A1(W26547), .A2(W4425), .ZN(O3847));
  NOR2X1 G10877 (.A1(W361), .A2(W35301), .ZN(O16109));
  NOR2X1 G10878 (.A1(W506), .A2(W1935), .ZN(W3859));
  NOR2X1 G10879 (.A1(W3764), .A2(W678), .ZN(W3858));
  NOR2X1 G10880 (.A1(W17940), .A2(W46459), .ZN(O16110));
  NOR2X1 G10881 (.A1(W1730), .A2(W3710), .ZN(W3856));
  NOR2X1 G10882 (.A1(W978), .A2(W22744), .ZN(W24080));
  NOR2X1 G10883 (.A1(W11552), .A2(W19173), .ZN(W26657));
  NOR2X1 G10884 (.A1(W14395), .A2(W8714), .ZN(W23936));
  NOR2X1 G10885 (.A1(W16102), .A2(W3446), .ZN(W23931));
  NOR2X1 G10886 (.A1(W4123), .A2(W2259), .ZN(W4275));
  NOR2X1 G10887 (.A1(W22546), .A2(W23903), .ZN(O15780));
  NOR2X1 G10888 (.A1(W17687), .A2(W15735), .ZN(W23932));
  NOR2X1 G10889 (.A1(W7933), .A2(I1594), .ZN(W26793));
  NOR2X1 G10890 (.A1(W25508), .A2(W15365), .ZN(W26792));
  NOR2X1 G10891 (.A1(W14064), .A2(W12262), .ZN(O3871));
  NOR2X1 G10892 (.A1(W17938), .A2(W705), .ZN(O15785));
  NOR2X1 G10893 (.A1(W45779), .A2(W46168), .ZN(O15777));
  NOR2X1 G10894 (.A1(W5337), .A2(W14045), .ZN(W23937));
  NOR2X1 G10895 (.A1(W20897), .A2(W8802), .ZN(O15788));
  NOR2X1 G10896 (.A1(W3672), .A2(W3526), .ZN(W4265));
  NOR2X1 G10897 (.A1(W14319), .A2(W5444), .ZN(W23938));
  NOR2X1 G10898 (.A1(W6748), .A2(W21179), .ZN(W23940));
  NOR2X1 G10899 (.A1(W12077), .A2(W13333), .ZN(W23941));
  NOR2X1 G10900 (.A1(W3801), .A2(W1296), .ZN(W4260));
  NOR2X1 G10901 (.A1(W428), .A2(W2095), .ZN(W4259));
  NOR2X1 G10902 (.A1(W18875), .A2(W1437), .ZN(O15773));
  NOR2X1 G10903 (.A1(W10376), .A2(W27052), .ZN(O15769));
  NOR2X1 G10904 (.A1(W3358), .A2(W3132), .ZN(W4294));
  NOR2X1 G10905 (.A1(W24620), .A2(W25115), .ZN(W26796));
  NOR2X1 G10906 (.A1(W4261), .A2(W1612), .ZN(W4292));
  NOR2X1 G10907 (.A1(W1613), .A2(I376), .ZN(W4290));
  NOR2X1 G10908 (.A1(W2008), .A2(W3738), .ZN(W4289));
  NOR2X1 G10909 (.A1(I1562), .A2(W2809), .ZN(W4288));
  NOR2X1 G10910 (.A1(W3152), .A2(W3355), .ZN(W4286));
  NOR2X1 G10911 (.A1(W16040), .A2(W20698), .ZN(W26784));
  NOR2X1 G10912 (.A1(I1858), .A2(W2541), .ZN(W4284));
  NOR2X1 G10913 (.A1(W15747), .A2(W34941), .ZN(O15774));
  NOR2X1 G10914 (.A1(W1004), .A2(I1195), .ZN(W4282));
  NOR2X1 G10915 (.A1(W37076), .A2(W11677), .ZN(O15775));
  NOR2X1 G10916 (.A1(W40813), .A2(W26644), .ZN(O15776));
  NOR2X1 G10917 (.A1(W18158), .A2(I362), .ZN(W23930));
  NOR2X1 G10918 (.A1(I937), .A2(W1185), .ZN(W4278));
  NOR2X1 G10919 (.A1(W3911), .A2(W3694), .ZN(O53));
  NOR2X1 G10920 (.A1(W3819), .A2(W347), .ZN(W4234));
  NOR2X1 G10921 (.A1(W2258), .A2(W4210), .ZN(W4233));
  NOR2X1 G10922 (.A1(W812), .A2(W4017), .ZN(W4232));
  NOR2X1 G10923 (.A1(W12850), .A2(W38152), .ZN(O15821));
  NOR2X1 G10924 (.A1(W3084), .A2(W711), .ZN(W4230));
  NOR2X1 G10925 (.A1(W26547), .A2(W1315), .ZN(O3865));
  NOR2X1 G10926 (.A1(I104), .A2(W1976), .ZN(W4228));
  NOR2X1 G10927 (.A1(W942), .A2(W4074), .ZN(W4227));
  NOR2X1 G10928 (.A1(W30850), .A2(W28239), .ZN(O15820));
  NOR2X1 G10929 (.A1(W107), .A2(W119), .ZN(W4225));
  NOR2X1 G10930 (.A1(W24101), .A2(W42967), .ZN(O15824));
  NOR2X1 G10931 (.A1(W3921), .A2(W3132), .ZN(W4222));
  NOR2X1 G10932 (.A1(W8659), .A2(I1003), .ZN(O3863));
  NOR2X1 G10933 (.A1(W20064), .A2(W17434), .ZN(W26770));
  NOR2X1 G10934 (.A1(W1682), .A2(I1325), .ZN(W4219));
  NOR2X1 G10935 (.A1(W9156), .A2(W23018), .ZN(O15827));
  NOR2X1 G10936 (.A1(W12610), .A2(W1179), .ZN(O15802));
  NOR2X1 G10937 (.A1(W21665), .A2(W22963), .ZN(W26783));
  NOR2X1 G10938 (.A1(W2772), .A2(W717), .ZN(W46733));
  NOR2X1 G10939 (.A1(W1053), .A2(W4108), .ZN(W4253));
  NOR2X1 G10940 (.A1(W26746), .A2(W12293), .ZN(W26780));
  NOR2X1 G10941 (.A1(W32064), .A2(W7041), .ZN(O15798));
  NOR2X1 G10942 (.A1(W19386), .A2(W19344), .ZN(W46739));
  NOR2X1 G10943 (.A1(I94), .A2(W6336), .ZN(W23948));
  NOR2X1 G10944 (.A1(W2094), .A2(W2213), .ZN(W4247));
  NOR2X1 G10945 (.A1(W2193), .A2(W23087), .ZN(O2924));
  NOR2X1 G10946 (.A1(W22918), .A2(W13001), .ZN(W26779));
  NOR2X1 G10947 (.A1(W9518), .A2(W9777), .ZN(O2929));
  NOR2X1 G10948 (.A1(W13214), .A2(W9013), .ZN(W26776));
  NOR2X1 G10949 (.A1(W16032), .A2(W16085), .ZN(W23954));
  NOR2X1 G10950 (.A1(W45525), .A2(I1430), .ZN(O15815));
  NOR2X1 G10951 (.A1(W14170), .A2(W6144), .ZN(O15818));
  NOR2X1 G10952 (.A1(W3813), .A2(W3323), .ZN(W4236));
  NOR2X1 G10953 (.A1(W13219), .A2(W10266), .ZN(W23914));
  NOR2X1 G10954 (.A1(W16964), .A2(W116), .ZN(W46648));
  NOR2X1 G10955 (.A1(W3528), .A2(W3064), .ZN(W4349));
  NOR2X1 G10956 (.A1(W3454), .A2(W2313), .ZN(W4348));
  NOR2X1 G10957 (.A1(W368), .A2(W3521), .ZN(W4347));
  NOR2X1 G10958 (.A1(W24256), .A2(W21473), .ZN(O3881));
  NOR2X1 G10959 (.A1(W5248), .A2(W18858), .ZN(W26808));
  NOR2X1 G10960 (.A1(W1330), .A2(W2813), .ZN(W4344));
  NOR2X1 G10961 (.A1(W3979), .A2(W3066), .ZN(W4343));
  NOR2X1 G10962 (.A1(W9275), .A2(W20738), .ZN(W23910));
  NOR2X1 G10963 (.A1(W3704), .A2(W192), .ZN(W4341));
  NOR2X1 G10964 (.A1(W24218), .A2(W37856), .ZN(O15730));
  NOR2X1 G10965 (.A1(I407), .A2(W87), .ZN(W4339));
  NOR2X1 G10966 (.A1(W18888), .A2(W19238), .ZN(O3880));
  NOR2X1 G10967 (.A1(W23783), .A2(W5837), .ZN(O15733));
  NOR2X1 G10968 (.A1(W39944), .A2(W12368), .ZN(W46661));
  NOR2X1 G10969 (.A1(W5616), .A2(W5037), .ZN(W26806));
  NOR2X1 G10970 (.A1(W777), .A2(W2849), .ZN(W4334));
  NOR2X1 G10971 (.A1(W178), .A2(I1803), .ZN(W4361));
  NOR2X1 G10972 (.A1(W45948), .A2(I486), .ZN(O15709));
  NOR2X1 G10973 (.A1(W1455), .A2(I1248), .ZN(W4371));
  NOR2X1 G10974 (.A1(W2948), .A2(W148), .ZN(W4370));
  NOR2X1 G10975 (.A1(I1994), .A2(I215), .ZN(W4369));
  NOR2X1 G10976 (.A1(W9502), .A2(W8887), .ZN(O15711));
  NOR2X1 G10977 (.A1(W39909), .A2(W35512), .ZN(O15713));
  NOR2X1 G10978 (.A1(W1148), .A2(W1780), .ZN(W4363));
  NOR2X1 G10979 (.A1(W5825), .A2(W12901), .ZN(W26813));
  NOR2X1 G10980 (.A1(W3483), .A2(W2388), .ZN(W4333));
  NOR2X1 G10981 (.A1(W15716), .A2(W15310), .ZN(O15715));
  NOR2X1 G10982 (.A1(W9682), .A2(W2693), .ZN(O3882));
  NOR2X1 G10983 (.A1(W13083), .A2(W14431), .ZN(W23909));
  NOR2X1 G10984 (.A1(I980), .A2(W3822), .ZN(W4356));
  NOR2X1 G10985 (.A1(W2005), .A2(W20788), .ZN(O15720));
  NOR2X1 G10986 (.A1(W43120), .A2(W5364), .ZN(O15721));
  NOR2X1 G10987 (.A1(W2767), .A2(W3640), .ZN(W4353));
  NOR2X1 G10988 (.A1(I875), .A2(W1062), .ZN(W4304));
  NOR2X1 G10989 (.A1(W166), .A2(W3507), .ZN(W4314));
  NOR2X1 G10990 (.A1(W9644), .A2(W7655), .ZN(O3876));
  NOR2X1 G10991 (.A1(W16827), .A2(W39074), .ZN(O15757));
  NOR2X1 G10992 (.A1(W4203), .A2(W3981), .ZN(W4309));
  NOR2X1 G10993 (.A1(W6486), .A2(I503), .ZN(W23924));
  NOR2X1 G10994 (.A1(W3451), .A2(I1055), .ZN(W4307));
  NOR2X1 G10995 (.A1(W6379), .A2(W37457), .ZN(O15760));
  NOR2X1 G10996 (.A1(I1245), .A2(W2424), .ZN(W4305));
  NOR2X1 G10997 (.A1(W2959), .A2(W2926), .ZN(O54));
  NOR2X1 G10998 (.A1(W3677), .A2(I371), .ZN(W4303));
  NOR2X1 G10999 (.A1(W181), .A2(W1362), .ZN(W4302));
  NOR2X1 G11000 (.A1(W2411), .A2(I294), .ZN(W4301));
  NOR2X1 G11001 (.A1(W12967), .A2(W3001), .ZN(O15763));
  NOR2X1 G11002 (.A1(W4268), .A2(W2442), .ZN(W4299));
  NOR2X1 G11003 (.A1(I1616), .A2(W613), .ZN(W4298));
  NOR2X1 G11004 (.A1(W7328), .A2(W6541), .ZN(W26797));
  NOR2X1 G11005 (.A1(W23210), .A2(W24109), .ZN(O15743));
  NOR2X1 G11006 (.A1(W701), .A2(W1849), .ZN(W4332));
  NOR2X1 G11007 (.A1(W3387), .A2(W3572), .ZN(W4331));
  NOR2X1 G11008 (.A1(W32366), .A2(W26538), .ZN(W46664));
  NOR2X1 G11009 (.A1(W4017), .A2(I1506), .ZN(W4329));
  NOR2X1 G11010 (.A1(W10245), .A2(W39575), .ZN(O15737));
  NOR2X1 G11011 (.A1(W58), .A2(I584), .ZN(W4327));
  NOR2X1 G11012 (.A1(W10179), .A2(W10605), .ZN(O2920));
  NOR2X1 G11013 (.A1(W44680), .A2(W29679), .ZN(O15742));
  NOR2X1 G11014 (.A1(W26), .A2(W716), .ZN(W4217));
  NOR2X1 G11015 (.A1(W30945), .A2(W21953), .ZN(O15744));
  NOR2X1 G11016 (.A1(W12509), .A2(W5983), .ZN(O3879));
  NOR2X1 G11017 (.A1(W30996), .A2(W34094), .ZN(O15746));
  NOR2X1 G11018 (.A1(W45245), .A2(W33494), .ZN(O15749));
  NOR2X1 G11019 (.A1(W45693), .A2(W1911), .ZN(O15750));
  NOR2X1 G11020 (.A1(I812), .A2(W1916), .ZN(W26803));
  NOR2X1 G11021 (.A1(W40276), .A2(W4480), .ZN(O15752));
  NOR2X1 G11022 (.A1(W21829), .A2(W20024), .ZN(O2942));
  NOR2X1 G11023 (.A1(W12682), .A2(W3805), .ZN(W23987));
  NOR2X1 G11024 (.A1(W1743), .A2(W3083), .ZN(W4124));
  NOR2X1 G11025 (.A1(W2293), .A2(W542), .ZN(W4123));
  NOR2X1 G11026 (.A1(I1075), .A2(W2181), .ZN(W4122));
  NOR2X1 G11027 (.A1(I114), .A2(W2967), .ZN(W4121));
  NOR2X1 G11028 (.A1(W11490), .A2(W11228), .ZN(W26742));
  NOR2X1 G11029 (.A1(W477), .A2(W16336), .ZN(O15894));
  NOR2X1 G11030 (.A1(W5234), .A2(W24039), .ZN(O15895));
  NOR2X1 G11031 (.A1(W24120), .A2(W2044), .ZN(W26745));
  NOR2X1 G11032 (.A1(W7132), .A2(W13428), .ZN(O3855));
  NOR2X1 G11033 (.A1(W11317), .A2(W4292), .ZN(W26740));
  NOR2X1 G11034 (.A1(W4974), .A2(W35084), .ZN(O15903));
  NOR2X1 G11035 (.A1(W3789), .A2(W1864), .ZN(W4113));
  NOR2X1 G11036 (.A1(W32262), .A2(W8924), .ZN(O15904));
  NOR2X1 G11037 (.A1(W4119), .A2(W15869), .ZN(O15905));
  NOR2X1 G11038 (.A1(W2745), .A2(W525), .ZN(W4110));
  NOR2X1 G11039 (.A1(W12573), .A2(W9058), .ZN(W23992));
  NOR2X1 G11040 (.A1(W2351), .A2(W16905), .ZN(W26749));
  NOR2X1 G11041 (.A1(W131), .A2(W438), .ZN(W4143));
  NOR2X1 G11042 (.A1(W7961), .A2(W27761), .ZN(W46833));
  NOR2X1 G11043 (.A1(W2626), .A2(W1215), .ZN(W4141));
  NOR2X1 G11044 (.A1(W16343), .A2(W34336), .ZN(W46834));
  NOR2X1 G11045 (.A1(W30330), .A2(W937), .ZN(O15880));
  NOR2X1 G11046 (.A1(W1743), .A2(W42453), .ZN(O15881));
  NOR2X1 G11047 (.A1(W812), .A2(W3455), .ZN(W4137));
  NOR2X1 G11048 (.A1(W3351), .A2(W1272), .ZN(W23980));
  NOR2X1 G11049 (.A1(W3724), .A2(W399), .ZN(W4108));
  NOR2X1 G11050 (.A1(W32643), .A2(W12723), .ZN(O15884));
  NOR2X1 G11051 (.A1(W14155), .A2(W4059), .ZN(W23982));
  NOR2X1 G11052 (.A1(W16343), .A2(W2358), .ZN(W26747));
  NOR2X1 G11053 (.A1(I1532), .A2(W570), .ZN(W4131));
  NOR2X1 G11054 (.A1(W24231), .A2(W20609), .ZN(W26746));
  NOR2X1 G11055 (.A1(W1065), .A2(W1942), .ZN(W4129));
  NOR2X1 G11056 (.A1(I1974), .A2(W4050), .ZN(W4128));
  NOR2X1 G11057 (.A1(W15779), .A2(W38504), .ZN(W46895));
  NOR2X1 G11058 (.A1(W3774), .A2(W2023), .ZN(W4089));
  NOR2X1 G11059 (.A1(W8856), .A2(W43835), .ZN(O15921));
  NOR2X1 G11060 (.A1(W14477), .A2(W1931), .ZN(W26733));
  NOR2X1 G11061 (.A1(I405), .A2(W4062), .ZN(W4085));
  NOR2X1 G11062 (.A1(W3315), .A2(W8495), .ZN(W23998));
  NOR2X1 G11063 (.A1(W9506), .A2(W13866), .ZN(W26731));
  NOR2X1 G11064 (.A1(W1132), .A2(W1197), .ZN(W4081));
  NOR2X1 G11065 (.A1(W17851), .A2(W35243), .ZN(W46894));
  NOR2X1 G11066 (.A1(W26626), .A2(W26588), .ZN(O15920));
  NOR2X1 G11067 (.A1(W33525), .A2(W5309), .ZN(O15930));
  NOR2X1 G11068 (.A1(W4172), .A2(W1910), .ZN(O2945));
  NOR2X1 G11069 (.A1(I267), .A2(W2356), .ZN(W4074));
  NOR2X1 G11070 (.A1(I941), .A2(W2189), .ZN(W4073));
  NOR2X1 G11071 (.A1(W45114), .A2(W15395), .ZN(O15935));
  NOR2X1 G11072 (.A1(W1262), .A2(W1142), .ZN(W4070));
  NOR2X1 G11073 (.A1(W2011), .A2(I1016), .ZN(W4068));
  NOR2X1 G11074 (.A1(W31634), .A2(W29808), .ZN(O15915));
  NOR2X1 G11075 (.A1(W2666), .A2(W2877), .ZN(W4107));
  NOR2X1 G11076 (.A1(W25598), .A2(W30886), .ZN(O15908));
  NOR2X1 G11077 (.A1(W11685), .A2(W23865), .ZN(O3852));
  NOR2X1 G11078 (.A1(I79), .A2(I204), .ZN(W4103));
  NOR2X1 G11079 (.A1(W33641), .A2(W32228), .ZN(O15912));
  NOR2X1 G11080 (.A1(W7562), .A2(W30121), .ZN(O15913));
  NOR2X1 G11081 (.A1(W37080), .A2(W36746), .ZN(O15914));
  NOR2X1 G11082 (.A1(W2636), .A2(I1681), .ZN(W4099));
  NOR2X1 G11083 (.A1(W26332), .A2(W23423), .ZN(W26751));
  NOR2X1 G11084 (.A1(W5252), .A2(W7878), .ZN(O2944));
  NOR2X1 G11085 (.A1(W7526), .A2(W15301), .ZN(O15917));
  NOR2X1 G11086 (.A1(I831), .A2(W44911), .ZN(W46881));
  NOR2X1 G11087 (.A1(W2673), .A2(W3181), .ZN(W4094));
  NOR2X1 G11088 (.A1(W1893), .A2(W647), .ZN(W4093));
  NOR2X1 G11089 (.A1(W24053), .A2(W39049), .ZN(O15919));
  NOR2X1 G11090 (.A1(W3599), .A2(I209), .ZN(W4091));
  NOR2X1 G11091 (.A1(W22964), .A2(W5310), .ZN(O2933));
  NOR2X1 G11092 (.A1(W28257), .A2(W22435), .ZN(O15847));
  NOR2X1 G11093 (.A1(W2417), .A2(W357), .ZN(W4197));
  NOR2X1 G11094 (.A1(I972), .A2(I1248), .ZN(W4196));
  NOR2X1 G11095 (.A1(W3473), .A2(W389), .ZN(W4195));
  NOR2X1 G11096 (.A1(W570), .A2(W3341), .ZN(W4194));
  NOR2X1 G11097 (.A1(W3540), .A2(W1700), .ZN(W4193));
  NOR2X1 G11098 (.A1(I681), .A2(W2432), .ZN(W4192));
  NOR2X1 G11099 (.A1(I66), .A2(W1519), .ZN(W4191));
  NOR2X1 G11100 (.A1(W18955), .A2(W13093), .ZN(W23965));
  NOR2X1 G11101 (.A1(W23349), .A2(W11381), .ZN(O15849));
  NOR2X1 G11102 (.A1(W3820), .A2(W1704), .ZN(W4188));
  NOR2X1 G11103 (.A1(W23526), .A2(W31186), .ZN(O15850));
  NOR2X1 G11104 (.A1(W14905), .A2(W10475), .ZN(O3861));
  NOR2X1 G11105 (.A1(W6365), .A2(W7304), .ZN(W26763));
  NOR2X1 G11106 (.A1(W18915), .A2(W6197), .ZN(O2935));
  NOR2X1 G11107 (.A1(W372), .A2(I603), .ZN(W4183));
  NOR2X1 G11108 (.A1(W35563), .A2(W1502), .ZN(O15855));
  NOR2X1 G11109 (.A1(W5451), .A2(W26957), .ZN(O15841));
  NOR2X1 G11110 (.A1(W21478), .A2(W10633), .ZN(W23960));
  NOR2X1 G11111 (.A1(W23), .A2(W372), .ZN(W4214));
  NOR2X1 G11112 (.A1(W26742), .A2(W23877), .ZN(O15830));
  NOR2X1 G11113 (.A1(W10825), .A2(W26687), .ZN(W26768));
  NOR2X1 G11114 (.A1(W25596), .A2(W21240), .ZN(O15832));
  NOR2X1 G11115 (.A1(W342), .A2(W14698), .ZN(W23963));
  NOR2X1 G11116 (.A1(W16604), .A2(W6767), .ZN(W26767));
  NOR2X1 G11117 (.A1(W3539), .A2(W41514), .ZN(W46786));
  NOR2X1 G11118 (.A1(W1925), .A2(I1952), .ZN(W4181));
  NOR2X1 G11119 (.A1(W942), .A2(I142), .ZN(W4206));
  NOR2X1 G11120 (.A1(W36063), .A2(W46560), .ZN(O15844));
  NOR2X1 G11121 (.A1(W21921), .A2(W25145), .ZN(O15846));
  NOR2X1 G11122 (.A1(W640), .A2(W3078), .ZN(W4203));
  NOR2X1 G11123 (.A1(W3560), .A2(W3603), .ZN(W4202));
  NOR2X1 G11124 (.A1(W1494), .A2(I947), .ZN(W4201));
  NOR2X1 G11125 (.A1(W144), .A2(W4197), .ZN(W4200));
  NOR2X1 G11126 (.A1(W1947), .A2(I1043), .ZN(W4153));
  NOR2X1 G11127 (.A1(I1604), .A2(W4000), .ZN(W4162));
  NOR2X1 G11128 (.A1(W13048), .A2(W4275), .ZN(O15868));
  NOR2X1 G11129 (.A1(W8026), .A2(W26821), .ZN(O15869));
  NOR2X1 G11130 (.A1(W612), .A2(I1970), .ZN(W4159));
  NOR2X1 G11131 (.A1(W11520), .A2(W4513), .ZN(O15871));
  NOR2X1 G11132 (.A1(W3385), .A2(W23322), .ZN(O15873));
  NOR2X1 G11133 (.A1(I659), .A2(W714), .ZN(W4155));
  NOR2X1 G11134 (.A1(W844), .A2(W82), .ZN(W26753));
  NOR2X1 G11135 (.A1(W39745), .A2(W1892), .ZN(W46817));
  NOR2X1 G11136 (.A1(I1343), .A2(W3677), .ZN(W4152));
  NOR2X1 G11137 (.A1(W2360), .A2(I730), .ZN(W4151));
  NOR2X1 G11138 (.A1(W35114), .A2(W35761), .ZN(O15874));
  NOR2X1 G11139 (.A1(W1913), .A2(W2230), .ZN(W4149));
  NOR2X1 G11140 (.A1(W7788), .A2(W16434), .ZN(O2937));
  NOR2X1 G11141 (.A1(W3200), .A2(I559), .ZN(W4146));
  NOR2X1 G11142 (.A1(W3537), .A2(W37572), .ZN(O15877));
  NOR2X1 G11143 (.A1(W13890), .A2(W21517), .ZN(W23971));
  NOR2X1 G11144 (.A1(W29715), .A2(W14485), .ZN(O15857));
  NOR2X1 G11145 (.A1(W16018), .A2(I1892), .ZN(W26761));
  NOR2X1 G11146 (.A1(W85), .A2(I948), .ZN(W4178));
  NOR2X1 G11147 (.A1(W4501), .A2(W4090), .ZN(O15860));
  NOR2X1 G11148 (.A1(W3251), .A2(I765), .ZN(W4176));
  NOR2X1 G11149 (.A1(W3764), .A2(W2791), .ZN(W4175));
  NOR2X1 G11150 (.A1(I950), .A2(W574), .ZN(W4174));
  NOR2X1 G11151 (.A1(W199), .A2(W2247), .ZN(W4173));
  NOR2X1 G11152 (.A1(W13359), .A2(W19300), .ZN(O17350));
  NOR2X1 G11153 (.A1(W5147), .A2(W71), .ZN(O15863));
  NOR2X1 G11154 (.A1(W14919), .A2(W9676), .ZN(O3859));
  NOR2X1 G11155 (.A1(W8447), .A2(W23871), .ZN(O2936));
  NOR2X1 G11156 (.A1(I943), .A2(I1105), .ZN(W4168));
  NOR2X1 G11157 (.A1(W29557), .A2(W45179), .ZN(W46815));
  NOR2X1 G11158 (.A1(W16194), .A2(W36926), .ZN(O15865));
  NOR2X1 G11159 (.A1(W376), .A2(W3965), .ZN(W4164));
  NOR2X1 G11160 (.A1(I1674), .A2(I1675), .ZN(W837));
  NOR2X1 G11161 (.A1(W7864), .A2(W13176), .ZN(O18923));
  NOR2X1 G11162 (.A1(W17413), .A2(W32826), .ZN(O18926));
  NOR2X1 G11163 (.A1(W4435), .A2(W19026), .ZN(O3281));
  NOR2X1 G11164 (.A1(I1686), .A2(I1687), .ZN(W843));
  NOR2X1 G11165 (.A1(W17499), .A2(W24622), .ZN(O3475));
  NOR2X1 G11166 (.A1(W7139), .A2(W34783), .ZN(O18931));
  NOR2X1 G11167 (.A1(W12349), .A2(I1638), .ZN(O3283));
  NOR2X1 G11168 (.A1(I1678), .A2(I1679), .ZN(W839));
  NOR2X1 G11169 (.A1(W18067), .A2(W3699), .ZN(W50148));
  NOR2X1 G11170 (.A1(W3973), .A2(W10795), .ZN(W25625));
  NOR2X1 G11171 (.A1(I1668), .A2(I1669), .ZN(W834));
  NOR2X1 G11172 (.A1(W11666), .A2(W10246), .ZN(O3473));
  NOR2X1 G11173 (.A1(W22404), .A2(W20088), .ZN(W25067));
  NOR2X1 G11174 (.A1(W25692), .A2(W1893), .ZN(O18943));
  NOR2X1 G11175 (.A1(I1658), .A2(I1659), .ZN(W829));
  NOR2X1 G11176 (.A1(I1656), .A2(I1657), .ZN(W828));
  NOR2X1 G11177 (.A1(W21255), .A2(W48788), .ZN(O18945));
  NOR2X1 G11178 (.A1(W12541), .A2(W22202), .ZN(W25051));
  NOR2X1 G11179 (.A1(I1738), .A2(I1739), .ZN(W869));
  NOR2X1 G11180 (.A1(W35033), .A2(W39099), .ZN(O18908));
  NOR2X1 G11181 (.A1(W10748), .A2(W19802), .ZN(O3478));
  NOR2X1 G11182 (.A1(I1732), .A2(I1733), .ZN(W866));
  NOR2X1 G11183 (.A1(I1730), .A2(I1731), .ZN(W865));
  NOR2X1 G11184 (.A1(I1728), .A2(I1729), .ZN(W864));
  NOR2X1 G11185 (.A1(I1724), .A2(I1725), .ZN(W862));
  NOR2X1 G11186 (.A1(W844), .A2(W43903), .ZN(O18912));
  NOR2X1 G11187 (.A1(I1650), .A2(I1651), .ZN(W825));
  NOR2X1 G11188 (.A1(W23375), .A2(W5587), .ZN(W25636));
  NOR2X1 G11189 (.A1(I1716), .A2(I1717), .ZN(W858));
  NOR2X1 G11190 (.A1(W43448), .A2(W16033), .ZN(O18915));
  NOR2X1 G11191 (.A1(I1710), .A2(I1711), .ZN(W855));
  NOR2X1 G11192 (.A1(W24800), .A2(W22329), .ZN(W25054));
  NOR2X1 G11193 (.A1(W17707), .A2(W48563), .ZN(O18921));
  NOR2X1 G11194 (.A1(I1702), .A2(I1703), .ZN(W851));
  NOR2X1 G11195 (.A1(W7029), .A2(I953), .ZN(O3466));
  NOR2X1 G11196 (.A1(W7595), .A2(W17060), .ZN(O3288));
  NOR2X1 G11197 (.A1(W16601), .A2(W9697), .ZN(O18963));
  NOR2X1 G11198 (.A1(W13928), .A2(W32395), .ZN(O18965));
  NOR2X1 G11199 (.A1(I1602), .A2(I1603), .ZN(W801));
  NOR2X1 G11200 (.A1(W8962), .A2(W14411), .ZN(W25080));
  NOR2X1 G11201 (.A1(I1598), .A2(I1599), .ZN(W799));
  NOR2X1 G11202 (.A1(I1596), .A2(I1597), .ZN(W798));
  NOR2X1 G11203 (.A1(I1592), .A2(I1593), .ZN(W796));
  NOR2X1 G11204 (.A1(W34097), .A2(W6526), .ZN(O18960));
  NOR2X1 G11205 (.A1(W604), .A2(W9835), .ZN(W25084));
  NOR2X1 G11206 (.A1(W45879), .A2(W45813), .ZN(O18975));
  NOR2X1 G11207 (.A1(W31257), .A2(W22705), .ZN(O18979));
  NOR2X1 G11208 (.A1(I1578), .A2(I1579), .ZN(W789));
  NOR2X1 G11209 (.A1(I1576), .A2(I1577), .ZN(W788));
  NOR2X1 G11210 (.A1(I1574), .A2(I1575), .ZN(W787));
  NOR2X1 G11211 (.A1(I1572), .A2(I1573), .ZN(O6));
  NOR2X1 G11212 (.A1(W48915), .A2(W9473), .ZN(O18980));
  NOR2X1 G11213 (.A1(I1632), .A2(I1633), .ZN(W816));
  NOR2X1 G11214 (.A1(W530), .A2(W9169), .ZN(W25069));
  NOR2X1 G11215 (.A1(I1646), .A2(I1647), .ZN(W823));
  NOR2X1 G11216 (.A1(I171), .A2(W14029), .ZN(W25619));
  NOR2X1 G11217 (.A1(I1201), .A2(W17090), .ZN(W25071));
  NOR2X1 G11218 (.A1(W1823), .A2(W16881), .ZN(W25616));
  NOR2X1 G11219 (.A1(I1638), .A2(I1639), .ZN(W819));
  NOR2X1 G11220 (.A1(I1636), .A2(I1637), .ZN(W818));
  NOR2X1 G11221 (.A1(W25099), .A2(W10534), .ZN(O3470));
  NOR2X1 G11222 (.A1(W37939), .A2(W29172), .ZN(O18905));
  NOR2X1 G11223 (.A1(W12248), .A2(W24629), .ZN(O18953));
  NOR2X1 G11224 (.A1(W15982), .A2(W21122), .ZN(W25613));
  NOR2X1 G11225 (.A1(W36091), .A2(W39925), .ZN(O18955));
  NOR2X1 G11226 (.A1(I482), .A2(W7235), .ZN(O18956));
  NOR2X1 G11227 (.A1(W14667), .A2(W23603), .ZN(O3287));
  NOR2X1 G11228 (.A1(W21771), .A2(W8222), .ZN(O18958));
  NOR2X1 G11229 (.A1(I1616), .A2(I1617), .ZN(W808));
  NOR2X1 G11230 (.A1(I1830), .A2(I1831), .ZN(W915));
  NOR2X1 G11231 (.A1(W45809), .A2(W19627), .ZN(O18851));
  NOR2X1 G11232 (.A1(I1846), .A2(I1847), .ZN(W923));
  NOR2X1 G11233 (.A1(W40800), .A2(I1233), .ZN(O18852));
  NOR2X1 G11234 (.A1(I1842), .A2(I1843), .ZN(W921));
  NOR2X1 G11235 (.A1(I1838), .A2(I1839), .ZN(W919));
  NOR2X1 G11236 (.A1(W23603), .A2(W25157), .ZN(O18854));
  NOR2X1 G11237 (.A1(I1834), .A2(I1835), .ZN(W917));
  NOR2X1 G11238 (.A1(W9912), .A2(W17345), .ZN(W25655));
  NOR2X1 G11239 (.A1(I1850), .A2(I1851), .ZN(W925));
  NOR2X1 G11240 (.A1(W15565), .A2(W3757), .ZN(W25036));
  NOR2X1 G11241 (.A1(W33137), .A2(W42453), .ZN(O18862));
  NOR2X1 G11242 (.A1(W10032), .A2(W48063), .ZN(O18863));
  NOR2X1 G11243 (.A1(W7888), .A2(W42177), .ZN(O18864));
  NOR2X1 G11244 (.A1(W22315), .A2(W4841), .ZN(O18865));
  NOR2X1 G11245 (.A1(W13509), .A2(W22797), .ZN(W25648));
  NOR2X1 G11246 (.A1(W4236), .A2(W26694), .ZN(O18869));
  NOR2X1 G11247 (.A1(W37945), .A2(W30316), .ZN(O18871));
  NOR2X1 G11248 (.A1(W15730), .A2(W12846), .ZN(O3272));
  NOR2X1 G11249 (.A1(I502), .A2(W16803), .ZN(O3489));
  NOR2X1 G11250 (.A1(I1886), .A2(I1887), .ZN(W943));
  NOR2X1 G11251 (.A1(W13334), .A2(W27551), .ZN(O18839));
  NOR2X1 G11252 (.A1(I1882), .A2(I1883), .ZN(W941));
  NOR2X1 G11253 (.A1(W22052), .A2(W1502), .ZN(O3487));
  NOR2X1 G11254 (.A1(W14590), .A2(W12054), .ZN(W25028));
  NOR2X1 G11255 (.A1(I1876), .A2(I1877), .ZN(W938));
  NOR2X1 G11256 (.A1(I1872), .A2(I1873), .ZN(W936));
  NOR2X1 G11257 (.A1(W8787), .A2(W17879), .ZN(O3482));
  NOR2X1 G11258 (.A1(W44337), .A2(W1949), .ZN(O18847));
  NOR2X1 G11259 (.A1(W20027), .A2(W19208), .ZN(W25031));
  NOR2X1 G11260 (.A1(I1864), .A2(I1865), .ZN(W932));
  NOR2X1 G11261 (.A1(W463), .A2(W3668), .ZN(O18849));
  NOR2X1 G11262 (.A1(I1860), .A2(I1861), .ZN(W930));
  NOR2X1 G11263 (.A1(I1858), .A2(I1859), .ZN(W929));
  NOR2X1 G11264 (.A1(I1852), .A2(I1853), .ZN(O7));
  NOR2X1 G11265 (.A1(W36076), .A2(W13131), .ZN(O18897));
  NOR2X1 G11266 (.A1(W17175), .A2(W558), .ZN(O18891));
  NOR2X1 G11267 (.A1(I1772), .A2(I1773), .ZN(W886));
  NOR2X1 G11268 (.A1(W9806), .A2(W12480), .ZN(W25047));
  NOR2X1 G11269 (.A1(W11373), .A2(W31299), .ZN(O18893));
  NOR2X1 G11270 (.A1(W42631), .A2(W24520), .ZN(O18894));
  NOR2X1 G11271 (.A1(W20600), .A2(W39661), .ZN(O18896));
  NOR2X1 G11272 (.A1(I1760), .A2(I1761), .ZN(W880));
  NOR2X1 G11273 (.A1(W23572), .A2(W19185), .ZN(W50121));
  NOR2X1 G11274 (.A1(W5319), .A2(W3888), .ZN(W25045));
  NOR2X1 G11275 (.A1(W48913), .A2(W25187), .ZN(W50123));
  NOR2X1 G11276 (.A1(I1752), .A2(I1753), .ZN(W876));
  NOR2X1 G11277 (.A1(W48235), .A2(W45367), .ZN(O18898));
  NOR2X1 G11278 (.A1(W24052), .A2(W7452), .ZN(O3278));
  NOR2X1 G11279 (.A1(I1746), .A2(I1747), .ZN(W873));
  NOR2X1 G11280 (.A1(W48274), .A2(W175), .ZN(O18902));
  NOR2X1 G11281 (.A1(W24044), .A2(W38579), .ZN(O18904));
  NOR2X1 G11282 (.A1(I1792), .A2(I1793), .ZN(W896));
  NOR2X1 G11283 (.A1(I1898), .A2(W15229), .ZN(W25645));
  NOR2X1 G11284 (.A1(W44821), .A2(W1694), .ZN(O18874));
  NOR2X1 G11285 (.A1(W39786), .A2(W38343), .ZN(O18876));
  NOR2X1 G11286 (.A1(W21492), .A2(W28763), .ZN(O18877));
  NOR2X1 G11287 (.A1(W1575), .A2(W10864), .ZN(O3480));
  NOR2X1 G11288 (.A1(I1798), .A2(I1799), .ZN(W899));
  NOR2X1 G11289 (.A1(W41648), .A2(W11933), .ZN(O18879));
  NOR2X1 G11290 (.A1(W42044), .A2(W20775), .ZN(O18880));
  NOR2X1 G11291 (.A1(I1568), .A2(I1569), .ZN(W784));
  NOR2X1 G11292 (.A1(W5176), .A2(W21904), .ZN(W25042));
  NOR2X1 G11293 (.A1(W44703), .A2(W35417), .ZN(O18882));
  NOR2X1 G11294 (.A1(W4899), .A2(W14501), .ZN(O3276));
  NOR2X1 G11295 (.A1(W2823), .A2(W26604), .ZN(O18886));
  NOR2X1 G11296 (.A1(W17951), .A2(W11098), .ZN(W25642));
  NOR2X1 G11297 (.A1(W12609), .A2(W10995), .ZN(O18888));
  NOR2X1 G11298 (.A1(W32328), .A2(W39052), .ZN(O18889));
  NOR2X1 G11299 (.A1(W14712), .A2(W24009), .ZN(O3308));
  NOR2X1 G11300 (.A1(I1372), .A2(I1373), .ZN(W686));
  NOR2X1 G11301 (.A1(W5299), .A2(W19675), .ZN(W25565));
  NOR2X1 G11302 (.A1(I1366), .A2(I1367), .ZN(W683));
  NOR2X1 G11303 (.A1(I1364), .A2(I1365), .ZN(W682));
  NOR2X1 G11304 (.A1(W23141), .A2(W45971), .ZN(O19098));
  NOR2X1 G11305 (.A1(I9), .A2(W6079), .ZN(O19099));
  NOR2X1 G11306 (.A1(W2090), .A2(W13641), .ZN(W25121));
  NOR2X1 G11307 (.A1(W9008), .A2(W19581), .ZN(W25122));
  NOR2X1 G11308 (.A1(W14465), .A2(I536), .ZN(O3459));
  NOR2X1 G11309 (.A1(I1352), .A2(I1353), .ZN(W676));
  NOR2X1 G11310 (.A1(W18614), .A2(W46833), .ZN(O19104));
  NOR2X1 G11311 (.A1(W32553), .A2(W17135), .ZN(O19105));
  NOR2X1 G11312 (.A1(I1346), .A2(I1347), .ZN(W673));
  NOR2X1 G11313 (.A1(W39408), .A2(W48706), .ZN(O19106));
  NOR2X1 G11314 (.A1(W5962), .A2(W13467), .ZN(O19108));
  NOR2X1 G11315 (.A1(W30819), .A2(W20456), .ZN(O19109));
  NOR2X1 G11316 (.A1(W14131), .A2(W21519), .ZN(O3309));
  NOR2X1 G11317 (.A1(I1392), .A2(I1393), .ZN(W696));
  NOR2X1 G11318 (.A1(W25054), .A2(W6829), .ZN(W25571));
  NOR2X1 G11319 (.A1(I1410), .A2(I1411), .ZN(W705));
  NOR2X1 G11320 (.A1(W38183), .A2(W23338), .ZN(O19070));
  NOR2X1 G11321 (.A1(I1402), .A2(I1403), .ZN(W701));
  NOR2X1 G11322 (.A1(I1400), .A2(I1401), .ZN(W700));
  NOR2X1 G11323 (.A1(I1398), .A2(I1399), .ZN(W699));
  NOR2X1 G11324 (.A1(W13491), .A2(W37987), .ZN(O19071));
  NOR2X1 G11325 (.A1(W23625), .A2(I1550), .ZN(W25114));
  NOR2X1 G11326 (.A1(W17368), .A2(W20633), .ZN(W25126));
  NOR2X1 G11327 (.A1(I1390), .A2(I1391), .ZN(W695));
  NOR2X1 G11328 (.A1(W8340), .A2(I1236), .ZN(O3460));
  NOR2X1 G11329 (.A1(W19363), .A2(W29213), .ZN(O19081));
  NOR2X1 G11330 (.A1(W47919), .A2(W35166), .ZN(O19085));
  NOR2X1 G11331 (.A1(I1380), .A2(I1381), .ZN(W690));
  NOR2X1 G11332 (.A1(W11763), .A2(W24664), .ZN(O19088));
  NOR2X1 G11333 (.A1(W20991), .A2(W12574), .ZN(O3306));
  NOR2X1 G11334 (.A1(W8888), .A2(W29029), .ZN(O19143));
  NOR2X1 G11335 (.A1(W38239), .A2(W9447), .ZN(O19132));
  NOR2X1 G11336 (.A1(W2010), .A2(W18508), .ZN(W25135));
  NOR2X1 G11337 (.A1(W19611), .A2(W21953), .ZN(O19136));
  NOR2X1 G11338 (.A1(I1288), .A2(I1289), .ZN(W644));
  NOR2X1 G11339 (.A1(W8945), .A2(W3979), .ZN(O19140));
  NOR2X1 G11340 (.A1(W33695), .A2(W45488), .ZN(O19141));
  NOR2X1 G11341 (.A1(I1282), .A2(I1283), .ZN(W641));
  NOR2X1 G11342 (.A1(I1280), .A2(I1281), .ZN(W640));
  NOR2X1 G11343 (.A1(W16019), .A2(W10415), .ZN(O3453));
  NOR2X1 G11344 (.A1(I1276), .A2(I1277), .ZN(W638));
  NOR2X1 G11345 (.A1(W1025), .A2(W23708), .ZN(O3452));
  NOR2X1 G11346 (.A1(I1272), .A2(I1273), .ZN(W636));
  NOR2X1 G11347 (.A1(I1599), .A2(I1226), .ZN(W25547));
  NOR2X1 G11348 (.A1(W8821), .A2(W23413), .ZN(W25140));
  NOR2X1 G11349 (.A1(W14103), .A2(W15580), .ZN(O3312));
  NOR2X1 G11350 (.A1(W36652), .A2(W33644), .ZN(O19150));
  NOR2X1 G11351 (.A1(I1316), .A2(I1317), .ZN(W658));
  NOR2X1 G11352 (.A1(I1332), .A2(I1333), .ZN(W666));
  NOR2X1 G11353 (.A1(W4142), .A2(W16486), .ZN(W25561));
  NOR2X1 G11354 (.A1(W43742), .A2(W5493), .ZN(O19114));
  NOR2X1 G11355 (.A1(W25538), .A2(W23971), .ZN(O19116));
  NOR2X1 G11356 (.A1(W22696), .A2(W18672), .ZN(W25128));
  NOR2X1 G11357 (.A1(W23662), .A2(W14914), .ZN(O3456));
  NOR2X1 G11358 (.A1(I1320), .A2(I1321), .ZN(W660));
  NOR2X1 G11359 (.A1(W1603), .A2(W23710), .ZN(O3455));
  NOR2X1 G11360 (.A1(I1414), .A2(I1415), .ZN(W707));
  NOR2X1 G11361 (.A1(W49353), .A2(W20054), .ZN(O19122));
  NOR2X1 G11362 (.A1(W49549), .A2(W13357), .ZN(O19123));
  NOR2X1 G11363 (.A1(W5620), .A2(W7464), .ZN(W25558));
  NOR2X1 G11364 (.A1(W503), .A2(W6488), .ZN(O19126));
  NOR2X1 G11365 (.A1(W34640), .A2(W19065), .ZN(O19128));
  NOR2X1 G11366 (.A1(W921), .A2(W5809), .ZN(W25133));
  NOR2X1 G11367 (.A1(I1300), .A2(I1301), .ZN(W650));
  NOR2X1 G11368 (.A1(W20665), .A2(W20065), .ZN(W25581));
  NOR2X1 G11369 (.A1(W14911), .A2(W18722), .ZN(O3463));
  NOR2X1 G11370 (.A1(W5619), .A2(W17434), .ZN(O19005));
  NOR2X1 G11371 (.A1(W22118), .A2(W34561), .ZN(O19006));
  NOR2X1 G11372 (.A1(W26301), .A2(W39572), .ZN(O19009));
  NOR2X1 G11373 (.A1(W44358), .A2(W46881), .ZN(O19012));
  NOR2X1 G11374 (.A1(W9454), .A2(W17702), .ZN(W25582));
  NOR2X1 G11375 (.A1(W17090), .A2(W48469), .ZN(O19014));
  NOR2X1 G11376 (.A1(I1508), .A2(I1509), .ZN(W754));
  NOR2X1 G11377 (.A1(W538), .A2(W15493), .ZN(O19000));
  NOR2X1 G11378 (.A1(W32373), .A2(W31672), .ZN(O19016));
  NOR2X1 G11379 (.A1(W30851), .A2(W6313), .ZN(O19018));
  NOR2X1 G11380 (.A1(W36017), .A2(W48541), .ZN(O19019));
  NOR2X1 G11381 (.A1(W43557), .A2(W2380), .ZN(W50250));
  NOR2X1 G11382 (.A1(W8038), .A2(W2737), .ZN(O19020));
  NOR2X1 G11383 (.A1(I1494), .A2(I1495), .ZN(W747));
  NOR2X1 G11384 (.A1(I1492), .A2(I1493), .ZN(W746));
  NOR2X1 G11385 (.A1(I1490), .A2(I1491), .ZN(W745));
  NOR2X1 G11386 (.A1(W43722), .A2(W45119), .ZN(O18992));
  NOR2X1 G11387 (.A1(I115), .A2(W8350), .ZN(W25601));
  NOR2X1 G11388 (.A1(W21505), .A2(W23269), .ZN(O18982));
  NOR2X1 G11389 (.A1(W171), .A2(W11321), .ZN(W25600));
  NOR2X1 G11390 (.A1(W39840), .A2(W21980), .ZN(O18984));
  NOR2X1 G11391 (.A1(I1556), .A2(I1557), .ZN(W778));
  NOR2X1 G11392 (.A1(I1033), .A2(W42773), .ZN(O18988));
  NOR2X1 G11393 (.A1(W18624), .A2(W854), .ZN(O3294));
  NOR2X1 G11394 (.A1(W10078), .A2(W15281), .ZN(W25597));
  NOR2X1 G11395 (.A1(I1626), .A2(W12684), .ZN(O3301));
  NOR2X1 G11396 (.A1(I1546), .A2(I1547), .ZN(W773));
  NOR2X1 G11397 (.A1(W18636), .A2(W14019), .ZN(W25594));
  NOR2X1 G11398 (.A1(I1540), .A2(I1541), .ZN(W770));
  NOR2X1 G11399 (.A1(I1822), .A2(W20233), .ZN(O3464));
  NOR2X1 G11400 (.A1(W18816), .A2(W25260), .ZN(W25591));
  NOR2X1 G11401 (.A1(W10015), .A2(W15315), .ZN(O3296));
  NOR2X1 G11402 (.A1(I1532), .A2(I1533), .ZN(W766));
  NOR2X1 G11403 (.A1(W48554), .A2(W18122), .ZN(O19051));
  NOR2X1 G11404 (.A1(W33757), .A2(W10191), .ZN(O19040));
  NOR2X1 G11405 (.A1(I1448), .A2(I1449), .ZN(W724));
  NOR2X1 G11406 (.A1(W20560), .A2(W30623), .ZN(O19045));
  NOR2X1 G11407 (.A1(I1444), .A2(I1445), .ZN(W722));
  NOR2X1 G11408 (.A1(W39352), .A2(W43224), .ZN(O19046));
  NOR2X1 G11409 (.A1(W24620), .A2(W1485), .ZN(O19048));
  NOR2X1 G11410 (.A1(I1438), .A2(I1439), .ZN(W719));
  NOR2X1 G11411 (.A1(W7710), .A2(W23692), .ZN(O3304));
  NOR2X1 G11412 (.A1(W6859), .A2(W25236), .ZN(O19039));
  NOR2X1 G11413 (.A1(I1430), .A2(I1431), .ZN(W715));
  NOR2X1 G11414 (.A1(I1428), .A2(I1429), .ZN(W714));
  NOR2X1 G11415 (.A1(I1426), .A2(I1427), .ZN(W713));
  NOR2X1 G11416 (.A1(I1424), .A2(I1425), .ZN(W712));
  NOR2X1 G11417 (.A1(W5211), .A2(W7712), .ZN(W25573));
  NOR2X1 G11418 (.A1(I1420), .A2(I1421), .ZN(W710));
  NOR2X1 G11419 (.A1(W9524), .A2(W5815), .ZN(O19057));
  NOR2X1 G11420 (.A1(W8939), .A2(W3218), .ZN(O19033));
  NOR2X1 G11421 (.A1(W3008), .A2(W45883), .ZN(O19022));
  NOR2X1 G11422 (.A1(W1722), .A2(W16506), .ZN(O19023));
  NOR2X1 G11423 (.A1(W48963), .A2(W29859), .ZN(O19024));
  NOR2X1 G11424 (.A1(W21401), .A2(W23890), .ZN(O19028));
  NOR2X1 G11425 (.A1(W27924), .A2(W29289), .ZN(O19029));
  NOR2X1 G11426 (.A1(W12269), .A2(W4065), .ZN(W25103));
  NOR2X1 G11427 (.A1(W25499), .A2(W13727), .ZN(O3462));
  NOR2X1 G11428 (.A1(I1472), .A2(I1473), .ZN(W736));
  NOR2X1 G11429 (.A1(I1892), .A2(I1893), .ZN(W946));
  NOR2X1 G11430 (.A1(W46948), .A2(W4224), .ZN(O19035));
  NOR2X1 G11431 (.A1(I1466), .A2(I1467), .ZN(W733));
  NOR2X1 G11432 (.A1(I1464), .A2(I1465), .ZN(W732));
  NOR2X1 G11433 (.A1(I1462), .A2(I1463), .ZN(W731));
  NOR2X1 G11434 (.A1(W24318), .A2(I1550), .ZN(W25578));
  NOR2X1 G11435 (.A1(I1458), .A2(I1459), .ZN(W729));
  NOR2X1 G11436 (.A1(W49495), .A2(W36687), .ZN(O19038));
  NOR2X1 G11437 (.A1(W30737), .A2(W6244), .ZN(O18651));
  NOR2X1 G11438 (.A1(W23000), .A2(I40), .ZN(O18643));
  NOR2X1 G11439 (.A1(W8039), .A2(W6682), .ZN(O3256));
  NOR2X1 G11440 (.A1(W10535), .A2(W46137), .ZN(O18645));
  NOR2X1 G11441 (.A1(W10880), .A2(W11793), .ZN(W24957));
  NOR2X1 G11442 (.A1(W12660), .A2(W31317), .ZN(O18648));
  NOR2X1 G11443 (.A1(W691), .A2(I568), .ZN(W1152));
  NOR2X1 G11444 (.A1(W177), .A2(I472), .ZN(W1150));
  NOR2X1 G11445 (.A1(W29668), .A2(W24529), .ZN(O18650));
  NOR2X1 G11446 (.A1(W14669), .A2(W8459), .ZN(O3513));
  NOR2X1 G11447 (.A1(W22204), .A2(W28974), .ZN(O18653));
  NOR2X1 G11448 (.A1(W31892), .A2(W16213), .ZN(O18654));
  NOR2X1 G11449 (.A1(W3724), .A2(W41035), .ZN(O18655));
  NOR2X1 G11450 (.A1(W33756), .A2(W5851), .ZN(O18656));
  NOR2X1 G11451 (.A1(I1602), .A2(W1119), .ZN(W1143));
  NOR2X1 G11452 (.A1(I920), .A2(W1042), .ZN(W1142));
  NOR2X1 G11453 (.A1(W837), .A2(W22374), .ZN(O18657));
  NOR2X1 G11454 (.A1(W8023), .A2(W15053), .ZN(O3511));
  NOR2X1 G11455 (.A1(W12587), .A2(W21041), .ZN(O3514));
  NOR2X1 G11456 (.A1(W1156), .A2(I248), .ZN(W1177));
  NOR2X1 G11457 (.A1(W5618), .A2(W5277), .ZN(O3251));
  NOR2X1 G11458 (.A1(I868), .A2(W234), .ZN(W1175));
  NOR2X1 G11459 (.A1(W27494), .A2(I882), .ZN(O18620));
  NOR2X1 G11460 (.A1(W28331), .A2(W23491), .ZN(O18623));
  NOR2X1 G11461 (.A1(W15052), .A2(W2058), .ZN(O18624));
  NOR2X1 G11462 (.A1(I280), .A2(I488), .ZN(W1171));
  NOR2X1 G11463 (.A1(I576), .A2(W11672), .ZN(W24949));
  NOR2X1 G11464 (.A1(W17198), .A2(W1933), .ZN(O18660));
  NOR2X1 G11465 (.A1(W4891), .A2(I1686), .ZN(W25746));
  NOR2X1 G11466 (.A1(W724), .A2(I1506), .ZN(O9));
  NOR2X1 G11467 (.A1(W30781), .A2(W23039), .ZN(O18631));
  NOR2X1 G11468 (.A1(W12533), .A2(W47287), .ZN(O18633));
  NOR2X1 G11469 (.A1(I365), .A2(I433), .ZN(W1163));
  NOR2X1 G11470 (.A1(I1628), .A2(I456), .ZN(W1161));
  NOR2X1 G11471 (.A1(W3350), .A2(W7229), .ZN(O3253));
  NOR2X1 G11472 (.A1(W22003), .A2(W4726), .ZN(O3507));
  NOR2X1 G11473 (.A1(I368), .A2(I1442), .ZN(W1116));
  NOR2X1 G11474 (.A1(W15196), .A2(W38220), .ZN(O18678));
  NOR2X1 G11475 (.A1(W8737), .A2(W48545), .ZN(O18679));
  NOR2X1 G11476 (.A1(I112), .A2(I1611), .ZN(W1113));
  NOR2X1 G11477 (.A1(W215), .A2(W1065), .ZN(W1112));
  NOR2X1 G11478 (.A1(W251), .A2(I366), .ZN(W1111));
  NOR2X1 G11479 (.A1(I446), .A2(I285), .ZN(W1110));
  NOR2X1 G11480 (.A1(I1442), .A2(I1612), .ZN(W1109));
  NOR2X1 G11481 (.A1(I1018), .A2(I1788), .ZN(W1117));
  NOR2X1 G11482 (.A1(W9000), .A2(W2885), .ZN(W24967));
  NOR2X1 G11483 (.A1(W27821), .A2(W4059), .ZN(O18685));
  NOR2X1 G11484 (.A1(I804), .A2(I435), .ZN(W1105));
  NOR2X1 G11485 (.A1(W5037), .A2(W18090), .ZN(O3260));
  NOR2X1 G11486 (.A1(I1921), .A2(I843), .ZN(W1103));
  NOR2X1 G11487 (.A1(W37161), .A2(W12454), .ZN(O18688));
  NOR2X1 G11488 (.A1(W620), .A2(I1862), .ZN(W1101));
  NOR2X1 G11489 (.A1(W38798), .A2(W11857), .ZN(O18671));
  NOR2X1 G11490 (.A1(I1255), .A2(I300), .ZN(W1138));
  NOR2X1 G11491 (.A1(W26977), .A2(W8176), .ZN(O18661));
  NOR2X1 G11492 (.A1(W14922), .A2(W18605), .ZN(O18662));
  NOR2X1 G11493 (.A1(W493), .A2(W539), .ZN(W1135));
  NOR2X1 G11494 (.A1(W7242), .A2(W16260), .ZN(O3509));
  NOR2X1 G11495 (.A1(W413), .A2(W890), .ZN(W1132));
  NOR2X1 G11496 (.A1(W28126), .A2(W19637), .ZN(O18667));
  NOR2X1 G11497 (.A1(W40679), .A2(W32992), .ZN(O18668));
  NOR2X1 G11498 (.A1(I1121), .A2(W667), .ZN(W1178));
  NOR2X1 G11499 (.A1(I590), .A2(I889), .ZN(W1127));
  NOR2X1 G11500 (.A1(W2774), .A2(W19175), .ZN(O18674));
  NOR2X1 G11501 (.A1(W905), .A2(I1608), .ZN(W1124));
  NOR2X1 G11502 (.A1(W950), .A2(I1801), .ZN(W1123));
  NOR2X1 G11503 (.A1(W9950), .A2(W18538), .ZN(O18675));
  NOR2X1 G11504 (.A1(W35388), .A2(W41582), .ZN(W49894));
  NOR2X1 G11505 (.A1(W99), .A2(I831), .ZN(W1118));
  NOR2X1 G11506 (.A1(W21668), .A2(W22559), .ZN(O3524));
  NOR2X1 G11507 (.A1(W34040), .A2(W28214), .ZN(O18551));
  NOR2X1 G11508 (.A1(W15373), .A2(W26648), .ZN(O18553));
  NOR2X1 G11509 (.A1(W46729), .A2(W16452), .ZN(O18555));
  NOR2X1 G11510 (.A1(W497), .A2(W1056), .ZN(O11));
  NOR2X1 G11511 (.A1(W20203), .A2(W49687), .ZN(O18557));
  NOR2X1 G11512 (.A1(W2440), .A2(W19221), .ZN(O18558));
  NOR2X1 G11513 (.A1(W540), .A2(W45718), .ZN(O18559));
  NOR2X1 G11514 (.A1(W494), .A2(W22909), .ZN(W49774));
  NOR2X1 G11515 (.A1(W796), .A2(I1841), .ZN(W1236));
  NOR2X1 G11516 (.A1(W3725), .A2(W32221), .ZN(O18564));
  NOR2X1 G11517 (.A1(W21076), .A2(W31445), .ZN(O18565));
  NOR2X1 G11518 (.A1(W92), .A2(I1717), .ZN(W1224));
  NOR2X1 G11519 (.A1(W865), .A2(W1181), .ZN(W1223));
  NOR2X1 G11520 (.A1(W477), .A2(I151), .ZN(W1222));
  NOR2X1 G11521 (.A1(W10286), .A2(W38529), .ZN(O18567));
  NOR2X1 G11522 (.A1(W5181), .A2(W5421), .ZN(W25769));
  NOR2X1 G11523 (.A1(W1139), .A2(I782), .ZN(W1219));
  NOR2X1 G11524 (.A1(W12234), .A2(W22195), .ZN(W25773));
  NOR2X1 G11525 (.A1(W953), .A2(W874), .ZN(W1255));
  NOR2X1 G11526 (.A1(W1163), .A2(W408), .ZN(W1253));
  NOR2X1 G11527 (.A1(W13017), .A2(W930), .ZN(O3243));
  NOR2X1 G11528 (.A1(W22922), .A2(W16199), .ZN(W25777));
  NOR2X1 G11529 (.A1(W2273), .A2(I541), .ZN(O18538));
  NOR2X1 G11530 (.A1(W6337), .A2(W39660), .ZN(O18542));
  NOR2X1 G11531 (.A1(I323), .A2(W298), .ZN(W1247));
  NOR2X1 G11532 (.A1(W27083), .A2(W15122), .ZN(O18543));
  NOR2X1 G11533 (.A1(W44560), .A2(W10092), .ZN(O18573));
  NOR2X1 G11534 (.A1(W667), .A2(I1506), .ZN(W1244));
  NOR2X1 G11535 (.A1(I889), .A2(W28051), .ZN(O18545));
  NOR2X1 G11536 (.A1(W11405), .A2(W43992), .ZN(W49756));
  NOR2X1 G11537 (.A1(W835), .A2(I1265), .ZN(W1241));
  NOR2X1 G11538 (.A1(I1620), .A2(W12591), .ZN(O18547));
  NOR2X1 G11539 (.A1(W6364), .A2(W7805), .ZN(W25771));
  NOR2X1 G11540 (.A1(W9082), .A2(W16060), .ZN(W24928));
  NOR2X1 G11541 (.A1(W23578), .A2(W21984), .ZN(W25755));
  NOR2X1 G11542 (.A1(W6259), .A2(W12857), .ZN(O18602));
  NOR2X1 G11543 (.A1(I1377), .A2(I1766), .ZN(W1194));
  NOR2X1 G11544 (.A1(W19789), .A2(W10581), .ZN(O3518));
  NOR2X1 G11545 (.A1(W33466), .A2(W35203), .ZN(O18603));
  NOR2X1 G11546 (.A1(W49660), .A2(W30105), .ZN(O18604));
  NOR2X1 G11547 (.A1(W467), .A2(I637), .ZN(W1190));
  NOR2X1 G11548 (.A1(W3912), .A2(W24191), .ZN(O18606));
  NOR2X1 G11549 (.A1(I862), .A2(W690), .ZN(W1188));
  NOR2X1 G11550 (.A1(W6197), .A2(W23639), .ZN(W25764));
  NOR2X1 G11551 (.A1(W5512), .A2(W21402), .ZN(W25753));
  NOR2X1 G11552 (.A1(I145), .A2(W16612), .ZN(W25752));
  NOR2X1 G11553 (.A1(W3628), .A2(W18689), .ZN(W24944));
  NOR2X1 G11554 (.A1(W14661), .A2(W47957), .ZN(O18615));
  NOR2X1 G11555 (.A1(I1450), .A2(I1003), .ZN(W1181));
  NOR2X1 G11556 (.A1(W767), .A2(W41735), .ZN(O18616));
  NOR2X1 G11557 (.A1(W1289), .A2(W18623), .ZN(W24946));
  NOR2X1 G11558 (.A1(I1040), .A2(I1544), .ZN(W1206));
  NOR2X1 G11559 (.A1(I1489), .A2(W152), .ZN(W1217));
  NOR2X1 G11560 (.A1(W563), .A2(W1594), .ZN(W24931));
  NOR2X1 G11561 (.A1(W3793), .A2(W20400), .ZN(O18577));
  NOR2X1 G11562 (.A1(W35875), .A2(W22066), .ZN(O18580));
  NOR2X1 G11563 (.A1(I1934), .A2(W16260), .ZN(O18581));
  NOR2X1 G11564 (.A1(W37456), .A2(W37942), .ZN(O18582));
  NOR2X1 G11565 (.A1(W4192), .A2(W21543), .ZN(W49796));
  NOR2X1 G11566 (.A1(W10265), .A2(W27523), .ZN(O18586));
  NOR2X1 G11567 (.A1(W37499), .A2(W46582), .ZN(O18689));
  NOR2X1 G11568 (.A1(W32635), .A2(W41056), .ZN(O18593));
  NOR2X1 G11569 (.A1(I1550), .A2(I718), .ZN(W1204));
  NOR2X1 G11570 (.A1(W8233), .A2(W22752), .ZN(O18594));
  NOR2X1 G11571 (.A1(W1011), .A2(W179), .ZN(W1202));
  NOR2X1 G11572 (.A1(W14699), .A2(W5936), .ZN(O3245));
  NOR2X1 G11573 (.A1(W7737), .A2(I1113), .ZN(W25765));
  NOR2X1 G11574 (.A1(I998), .A2(I1303), .ZN(W1199));
  NOR2X1 G11575 (.A1(I1990), .A2(I1991), .ZN(W995));
  NOR2X1 G11576 (.A1(I1284), .A2(I1611), .ZN(W1005));
  NOR2X1 G11577 (.A1(W49615), .A2(W47994), .ZN(O18787));
  NOR2X1 G11578 (.A1(W37198), .A2(W16614), .ZN(O18789));
  NOR2X1 G11579 (.A1(W10748), .A2(W30930), .ZN(O18791));
  NOR2X1 G11580 (.A1(W23881), .A2(W18564), .ZN(O18792));
  NOR2X1 G11581 (.A1(W36540), .A2(W33325), .ZN(O18793));
  NOR2X1 G11582 (.A1(I1996), .A2(I1997), .ZN(W998));
  NOR2X1 G11583 (.A1(W11623), .A2(W21668), .ZN(W25690));
  NOR2X1 G11584 (.A1(I204), .A2(I1672), .ZN(W1006));
  NOR2X1 G11585 (.A1(W2743), .A2(W23068), .ZN(W25009));
  NOR2X1 G11586 (.A1(I1984), .A2(I1985), .ZN(W992));
  NOR2X1 G11587 (.A1(I1982), .A2(I1983), .ZN(W991));
  NOR2X1 G11588 (.A1(I1980), .A2(I1981), .ZN(W990));
  NOR2X1 G11589 (.A1(I1978), .A2(I1979), .ZN(W989));
  NOR2X1 G11590 (.A1(I1976), .A2(I1977), .ZN(W988));
  NOR2X1 G11591 (.A1(I1259), .A2(W19951), .ZN(O18805));
  NOR2X1 G11592 (.A1(W15976), .A2(W10379), .ZN(O18806));
  NOR2X1 G11593 (.A1(W24071), .A2(W14610), .ZN(O3495));
  NOR2X1 G11594 (.A1(I1812), .A2(W952), .ZN(W1023));
  NOR2X1 G11595 (.A1(W9111), .A2(W16451), .ZN(W24999));
  NOR2X1 G11596 (.A1(I396), .A2(I765), .ZN(W1021));
  NOR2X1 G11597 (.A1(I926), .A2(I1105), .ZN(W1020));
  NOR2X1 G11598 (.A1(W3544), .A2(W14664), .ZN(O3496));
  NOR2X1 G11599 (.A1(W12961), .A2(W2569), .ZN(W25697));
  NOR2X1 G11600 (.A1(W10067), .A2(W15714), .ZN(W25002));
  NOR2X1 G11601 (.A1(I1377), .A2(I1831), .ZN(W1016));
  NOR2X1 G11602 (.A1(W1038), .A2(I1769), .ZN(W25683));
  NOR2X1 G11603 (.A1(W31595), .A2(W35333), .ZN(O18783));
  NOR2X1 G11604 (.A1(W406), .A2(I1233), .ZN(W1012));
  NOR2X1 G11605 (.A1(I1532), .A2(W312), .ZN(W1011));
  NOR2X1 G11606 (.A1(W36723), .A2(W39992), .ZN(O18784));
  NOR2X1 G11607 (.A1(I1681), .A2(I857), .ZN(W1009));
  NOR2X1 G11608 (.A1(W23031), .A2(W1738), .ZN(W25005));
  NOR2X1 G11609 (.A1(W540), .A2(I1828), .ZN(W1007));
  NOR2X1 G11610 (.A1(I1910), .A2(I1911), .ZN(W955));
  NOR2X1 G11611 (.A1(W6507), .A2(W1237), .ZN(W25022));
  NOR2X1 G11612 (.A1(W9513), .A2(W23463), .ZN(O3490));
  NOR2X1 G11613 (.A1(I1922), .A2(I1923), .ZN(W961));
  NOR2X1 G11614 (.A1(I1920), .A2(I1921), .ZN(W960));
  NOR2X1 G11615 (.A1(I1918), .A2(I1919), .ZN(W959));
  NOR2X1 G11616 (.A1(I1916), .A2(I1917), .ZN(W958));
  NOR2X1 G11617 (.A1(W37991), .A2(W30662), .ZN(O18834));
  NOR2X1 G11618 (.A1(I1912), .A2(I1913), .ZN(W956));
  NOR2X1 G11619 (.A1(I1930), .A2(I1931), .ZN(W965));
  NOR2X1 G11620 (.A1(I1908), .A2(I1909), .ZN(W954));
  NOR2X1 G11621 (.A1(I1906), .A2(I1907), .ZN(W953));
  NOR2X1 G11622 (.A1(W8192), .A2(W1385), .ZN(O18835));
  NOR2X1 G11623 (.A1(I1902), .A2(I1903), .ZN(W951));
  NOR2X1 G11624 (.A1(I1900), .A2(I1901), .ZN(W950));
  NOR2X1 G11625 (.A1(W44141), .A2(W24540), .ZN(O18837));
  NOR2X1 G11626 (.A1(I1894), .A2(I1895), .ZN(W947));
  NOR2X1 G11627 (.A1(W2901), .A2(W2800), .ZN(O18818));
  NOR2X1 G11628 (.A1(I1968), .A2(I1969), .ZN(W984));
  NOR2X1 G11629 (.A1(W4713), .A2(W8584), .ZN(W25012));
  NOR2X1 G11630 (.A1(W4898), .A2(W18300), .ZN(W25675));
  NOR2X1 G11631 (.A1(W10293), .A2(W12691), .ZN(W25015));
  NOR2X1 G11632 (.A1(W10097), .A2(W5408), .ZN(W25016));
  NOR2X1 G11633 (.A1(I1956), .A2(I1957), .ZN(W978));
  NOR2X1 G11634 (.A1(W24059), .A2(W49839), .ZN(O18816));
  NOR2X1 G11635 (.A1(W31477), .A2(W36505), .ZN(O18817));
  NOR2X1 G11636 (.A1(I324), .A2(I1187), .ZN(W1024));
  NOR2X1 G11637 (.A1(I521), .A2(W22430), .ZN(W25018));
  NOR2X1 G11638 (.A1(W3305), .A2(W19005), .ZN(W25671));
  NOR2X1 G11639 (.A1(I1942), .A2(I1943), .ZN(W971));
  NOR2X1 G11640 (.A1(I1940), .A2(I1941), .ZN(W970));
  NOR2X1 G11641 (.A1(W30084), .A2(W42900), .ZN(O18823));
  NOR2X1 G11642 (.A1(I1934), .A2(I1935), .ZN(W967));
  NOR2X1 G11643 (.A1(I1932), .A2(I1933), .ZN(W966));
  NOR2X1 G11644 (.A1(W3556), .A2(W8718), .ZN(O18719));
  NOR2X1 G11645 (.A1(I144), .A2(W384), .ZN(W1079));
  NOR2X1 G11646 (.A1(W42432), .A2(W16880), .ZN(O18711));
  NOR2X1 G11647 (.A1(W10207), .A2(I1331), .ZN(O18713));
  NOR2X1 G11648 (.A1(W527), .A2(W18183), .ZN(O3263));
  NOR2X1 G11649 (.A1(W6588), .A2(W47180), .ZN(O18716));
  NOR2X1 G11650 (.A1(I1333), .A2(W49), .ZN(W1074));
  NOR2X1 G11651 (.A1(I1934), .A2(I1030), .ZN(W1073));
  NOR2X1 G11652 (.A1(W985), .A2(W44), .ZN(O3264));
  NOR2X1 G11653 (.A1(W13264), .A2(W39424), .ZN(O18708));
  NOR2X1 G11654 (.A1(W418), .A2(I1395), .ZN(W1070));
  NOR2X1 G11655 (.A1(W12316), .A2(W23740), .ZN(O18721));
  NOR2X1 G11656 (.A1(W26011), .A2(W15197), .ZN(O18723));
  NOR2X1 G11657 (.A1(W13458), .A2(W25718), .ZN(O18724));
  NOR2X1 G11658 (.A1(W23791), .A2(W22926), .ZN(O18726));
  NOR2X1 G11659 (.A1(W43147), .A2(W33864), .ZN(O18727));
  NOR2X1 G11660 (.A1(W9006), .A2(W22481), .ZN(W24978));
  NOR2X1 G11661 (.A1(W36130), .A2(W36), .ZN(O18731));
  NOR2X1 G11662 (.A1(W608), .A2(I1769), .ZN(W1091));
  NOR2X1 G11663 (.A1(I581), .A2(W741), .ZN(W1099));
  NOR2X1 G11664 (.A1(I1283), .A2(I492), .ZN(W1098));
  NOR2X1 G11665 (.A1(W348), .A2(I1573), .ZN(W1097));
  NOR2X1 G11666 (.A1(W15117), .A2(W34311), .ZN(O18691));
  NOR2X1 G11667 (.A1(W10517), .A2(W13017), .ZN(W24969));
  NOR2X1 G11668 (.A1(W17905), .A2(W21518), .ZN(W24970));
  NOR2X1 G11669 (.A1(W11989), .A2(W46402), .ZN(O18694));
  NOR2X1 G11670 (.A1(W22898), .A2(W8299), .ZN(W24971));
  NOR2X1 G11671 (.A1(W996), .A2(W742), .ZN(W1061));
  NOR2X1 G11672 (.A1(I540), .A2(W320), .ZN(W1090));
  NOR2X1 G11673 (.A1(W10150), .A2(W35944), .ZN(O18700));
  NOR2X1 G11674 (.A1(W81), .A2(I598), .ZN(W1088));
  NOR2X1 G11675 (.A1(W33997), .A2(W38199), .ZN(O18702));
  NOR2X1 G11676 (.A1(W3700), .A2(W17655), .ZN(W25724));
  NOR2X1 G11677 (.A1(W837), .A2(W1001), .ZN(W1083));
  NOR2X1 G11678 (.A1(W23229), .A2(W44765), .ZN(O18706));
  NOR2X1 G11679 (.A1(W621), .A2(W672), .ZN(W1033));
  NOR2X1 G11680 (.A1(W20442), .A2(W11409), .ZN(W24987));
  NOR2X1 G11681 (.A1(W14589), .A2(W6757), .ZN(O3500));
  NOR2X1 G11682 (.A1(W453), .A2(I1416), .ZN(W1039));
  NOR2X1 G11683 (.A1(W46624), .A2(W40716), .ZN(O18759));
  NOR2X1 G11684 (.A1(W847), .A2(I404), .ZN(W1037));
  NOR2X1 G11685 (.A1(W3349), .A2(W23420), .ZN(W25706));
  NOR2X1 G11686 (.A1(I1196), .A2(W599), .ZN(W1035));
  NOR2X1 G11687 (.A1(W13677), .A2(W18794), .ZN(O18763));
  NOR2X1 G11688 (.A1(W33691), .A2(W13456), .ZN(O18754));
  NOR2X1 G11689 (.A1(W16377), .A2(W21061), .ZN(W24991));
  NOR2X1 G11690 (.A1(W3194), .A2(W6240), .ZN(W24993));
  NOR2X1 G11691 (.A1(W13441), .A2(W22515), .ZN(O3499));
  NOR2X1 G11692 (.A1(I1569), .A2(W10964), .ZN(W25700));
  NOR2X1 G11693 (.A1(W5636), .A2(W4764), .ZN(W25699));
  NOR2X1 G11694 (.A1(W1070), .A2(W19235), .ZN(W24997));
  NOR2X1 G11695 (.A1(W4532), .A2(W16027), .ZN(W24998));
  NOR2X1 G11696 (.A1(W974), .A2(I1106), .ZN(W1051));
  NOR2X1 G11697 (.A1(I1646), .A2(W463), .ZN(W1060));
  NOR2X1 G11698 (.A1(W21588), .A2(W37164), .ZN(O18735));
  NOR2X1 G11699 (.A1(W6117), .A2(W4308), .ZN(O18737));
  NOR2X1 G11700 (.A1(W10999), .A2(W9731), .ZN(W24980));
  NOR2X1 G11701 (.A1(W14397), .A2(W2171), .ZN(W25712));
  NOR2X1 G11702 (.A1(I1362), .A2(W663), .ZN(W1054));
  NOR2X1 G11703 (.A1(I511), .A2(I1893), .ZN(W1053));
  NOR2X1 G11704 (.A1(I29), .A2(W9125), .ZN(O18745));
  NOR2X1 G11705 (.A1(W20714), .A2(W21045), .ZN(W25546));
  NOR2X1 G11706 (.A1(I414), .A2(W48877), .ZN(O18746));
  NOR2X1 G11707 (.A1(W18440), .A2(W5163), .ZN(W24983));
  NOR2X1 G11708 (.A1(W15709), .A2(W3935), .ZN(W49966));
  NOR2X1 G11709 (.A1(W16164), .A2(W18353), .ZN(W24984));
  NOR2X1 G11710 (.A1(I506), .A2(W8543), .ZN(O3501));
  NOR2X1 G11711 (.A1(W232), .A2(W106), .ZN(W1045));
  NOR2X1 G11712 (.A1(W21556), .A2(W23652), .ZN(W24986));
  NOR2X1 G11713 (.A1(W1642), .A2(W783), .ZN(W25413));
  NOR2X1 G11714 (.A1(I442), .A2(I443), .ZN(W221));
  NOR2X1 G11715 (.A1(I440), .A2(I441), .ZN(W220));
  NOR2X1 G11716 (.A1(W4168), .A2(W11863), .ZN(W25419));
  NOR2X1 G11717 (.A1(I434), .A2(I435), .ZN(W217));
  NOR2X1 G11718 (.A1(W16677), .A2(W12812), .ZN(O19538));
  NOR2X1 G11719 (.A1(I430), .A2(I431), .ZN(W215));
  NOR2X1 G11720 (.A1(W10913), .A2(W47308), .ZN(O19540));
  NOR2X1 G11721 (.A1(W24928), .A2(W9342), .ZN(O3413));
  NOR2X1 G11722 (.A1(I444), .A2(I445), .ZN(W222));
  NOR2X1 G11723 (.A1(I420), .A2(I421), .ZN(W210));
  NOR2X1 G11724 (.A1(I416), .A2(I417), .ZN(W208));
  NOR2X1 G11725 (.A1(I414), .A2(I415), .ZN(W207));
  NOR2X1 G11726 (.A1(I412), .A2(I413), .ZN(W206));
  NOR2X1 G11727 (.A1(I406), .A2(I407), .ZN(W203));
  NOR2X1 G11728 (.A1(W36832), .A2(W43679), .ZN(O19550));
  NOR2X1 G11729 (.A1(W2759), .A2(W47886), .ZN(O19552));
  NOR2X1 G11730 (.A1(I400), .A2(I401), .ZN(W200));
  NOR2X1 G11731 (.A1(I462), .A2(I463), .ZN(W231));
  NOR2X1 G11732 (.A1(I480), .A2(I481), .ZN(W240));
  NOR2X1 G11733 (.A1(W42606), .A2(W29144), .ZN(O19512));
  NOR2X1 G11734 (.A1(W14932), .A2(W30268), .ZN(O19516));
  NOR2X1 G11735 (.A1(W23528), .A2(W15391), .ZN(O3347));
  NOR2X1 G11736 (.A1(W12023), .A2(W17217), .ZN(O19520));
  NOR2X1 G11737 (.A1(W21055), .A2(W13535), .ZN(O19521));
  NOR2X1 G11738 (.A1(I468), .A2(I469), .ZN(W234));
  NOR2X1 G11739 (.A1(I466), .A2(I467), .ZN(W233));
  NOR2X1 G11740 (.A1(W12459), .A2(W20902), .ZN(W25407));
  NOR2X1 G11741 (.A1(W24215), .A2(W24090), .ZN(W25422));
  NOR2X1 G11742 (.A1(I458), .A2(I459), .ZN(W229));
  NOR2X1 G11743 (.A1(W16702), .A2(W5158), .ZN(O19526));
  NOR2X1 G11744 (.A1(I454), .A2(I455), .ZN(W227));
  NOR2X1 G11745 (.A1(W47689), .A2(W14040), .ZN(O19529));
  NOR2X1 G11746 (.A1(W322), .A2(W36768), .ZN(O19533));
  NOR2X1 G11747 (.A1(I446), .A2(I447), .ZN(W223));
  NOR2X1 G11748 (.A1(I336), .A2(I337), .ZN(W168));
  NOR2X1 G11749 (.A1(I540), .A2(W21381), .ZN(W25280));
  NOR2X1 G11750 (.A1(W33470), .A2(W24687), .ZN(O19578));
  NOR2X1 G11751 (.A1(I1526), .A2(W10486), .ZN(W25401));
  NOR2X1 G11752 (.A1(W13464), .A2(W15664), .ZN(O3357));
  NOR2X1 G11753 (.A1(I346), .A2(I347), .ZN(W173));
  NOR2X1 G11754 (.A1(W12164), .A2(W20532), .ZN(W25285));
  NOR2X1 G11755 (.A1(W12794), .A2(W23621), .ZN(O3359));
  NOR2X1 G11756 (.A1(I338), .A2(I339), .ZN(W169));
  NOR2X1 G11757 (.A1(W27088), .A2(W1271), .ZN(O19576));
  NOR2X1 G11758 (.A1(I334), .A2(I335), .ZN(W167));
  NOR2X1 G11759 (.A1(I330), .A2(I331), .ZN(W165));
  NOR2X1 G11760 (.A1(W5927), .A2(W22854), .ZN(W25289));
  NOR2X1 G11761 (.A1(W8960), .A2(W14968), .ZN(O19592));
  NOR2X1 G11762 (.A1(W20182), .A2(W20409), .ZN(W25393));
  NOR2X1 G11763 (.A1(W38542), .A2(W11230), .ZN(O19594));
  NOR2X1 G11764 (.A1(W6218), .A2(W17721), .ZN(W25291));
  NOR2X1 G11765 (.A1(W19876), .A2(W23918), .ZN(W25392));
  NOR2X1 G11766 (.A1(W10904), .A2(W9985), .ZN(O3410));
  NOR2X1 G11767 (.A1(W36358), .A2(W3710), .ZN(O19554));
  NOR2X1 G11768 (.A1(W35845), .A2(W5519), .ZN(O19555));
  NOR2X1 G11769 (.A1(W15156), .A2(W23519), .ZN(W25406));
  NOR2X1 G11770 (.A1(W10341), .A2(W20039), .ZN(O19559));
  NOR2X1 G11771 (.A1(W39133), .A2(W1658), .ZN(O19560));
  NOR2X1 G11772 (.A1(W13837), .A2(W9802), .ZN(O3353));
  NOR2X1 G11773 (.A1(I384), .A2(I385), .ZN(W192));
  NOR2X1 G11774 (.A1(W11948), .A2(W16984), .ZN(O19562));
  NOR2X1 G11775 (.A1(W441), .A2(W8507), .ZN(O19511));
  NOR2X1 G11776 (.A1(W23998), .A2(W928), .ZN(W25276));
  NOR2X1 G11777 (.A1(I374), .A2(I375), .ZN(W187));
  NOR2X1 G11778 (.A1(W41194), .A2(W50148), .ZN(O19568));
  NOR2X1 G11779 (.A1(W12415), .A2(W11091), .ZN(W25278));
  NOR2X1 G11780 (.A1(W7495), .A2(W2650), .ZN(O3356));
  NOR2X1 G11781 (.A1(I364), .A2(I365), .ZN(W182));
  NOR2X1 G11782 (.A1(W48577), .A2(W7743), .ZN(O19575));
  NOR2X1 G11783 (.A1(I582), .A2(I583), .ZN(W291));
  NOR2X1 G11784 (.A1(W32169), .A2(W39644), .ZN(O19452));
  NOR2X1 G11785 (.A1(W9573), .A2(W45566), .ZN(O19456));
  NOR2X1 G11786 (.A1(W22867), .A2(W39600), .ZN(O19457));
  NOR2X1 G11787 (.A1(I812), .A2(W9265), .ZN(O19465));
  NOR2X1 G11788 (.A1(W2993), .A2(W42259), .ZN(O19468));
  NOR2X1 G11789 (.A1(W47260), .A2(W35409), .ZN(O19469));
  NOR2X1 G11790 (.A1(W14062), .A2(W868), .ZN(W25450));
  NOR2X1 G11791 (.A1(W12813), .A2(W16140), .ZN(O19471));
  NOR2X1 G11792 (.A1(W32879), .A2(W46213), .ZN(O19451));
  NOR2X1 G11793 (.A1(I578), .A2(I579), .ZN(W289));
  NOR2X1 G11794 (.A1(W6575), .A2(W18310), .ZN(W25445));
  NOR2X1 G11795 (.A1(W41290), .A2(W35564), .ZN(O19477));
  NOR2X1 G11796 (.A1(W19549), .A2(W12453), .ZN(W25444));
  NOR2X1 G11797 (.A1(W24040), .A2(W15), .ZN(O3425));
  NOR2X1 G11798 (.A1(W40805), .A2(I1025), .ZN(O19480));
  NOR2X1 G11799 (.A1(I566), .A2(I567), .ZN(W283));
  NOR2X1 G11800 (.A1(I562), .A2(I563), .ZN(W281));
  NOR2X1 G11801 (.A1(W4491), .A2(W20678), .ZN(W25236));
  NOR2X1 G11802 (.A1(I638), .A2(I639), .ZN(W319));
  NOR2X1 G11803 (.A1(I636), .A2(I637), .ZN(W318));
  NOR2X1 G11804 (.A1(I634), .A2(I635), .ZN(W317));
  NOR2X1 G11805 (.A1(I632), .A2(I633), .ZN(W316));
  NOR2X1 G11806 (.A1(I630), .A2(I631), .ZN(W315));
  NOR2X1 G11807 (.A1(I628), .A2(I629), .ZN(W314));
  NOR2X1 G11808 (.A1(W22238), .A2(W49262), .ZN(O19443));
  NOR2X1 G11809 (.A1(I624), .A2(I625), .ZN(W312));
  NOR2X1 G11810 (.A1(W21913), .A2(W489), .ZN(O19483));
  NOR2X1 G11811 (.A1(I620), .A2(I621), .ZN(W310));
  NOR2X1 G11812 (.A1(I618), .A2(I619), .ZN(W309));
  NOR2X1 G11813 (.A1(W49426), .A2(W43081), .ZN(O19446));
  NOR2X1 G11814 (.A1(I614), .A2(I615), .ZN(W307));
  NOR2X1 G11815 (.A1(I612), .A2(I613), .ZN(W306));
  NOR2X1 G11816 (.A1(W48183), .A2(W7170), .ZN(O19449));
  NOR2X1 G11817 (.A1(I606), .A2(I607), .ZN(W303));
  NOR2X1 G11818 (.A1(W10044), .A2(W14525), .ZN(O19500));
  NOR2X1 G11819 (.A1(I753), .A2(W17068), .ZN(O3422));
  NOR2X1 G11820 (.A1(I520), .A2(I521), .ZN(W260));
  NOR2X1 G11821 (.A1(I518), .A2(I519), .ZN(W259));
  NOR2X1 G11822 (.A1(I516), .A2(I517), .ZN(W258));
  NOR2X1 G11823 (.A1(W10765), .A2(W12902), .ZN(W25436));
  NOR2X1 G11824 (.A1(W4434), .A2(W19219), .ZN(O3420));
  NOR2X1 G11825 (.A1(I510), .A2(I511), .ZN(W255));
  NOR2X1 G11826 (.A1(W19629), .A2(W12692), .ZN(O19498));
  NOR2X1 G11827 (.A1(I524), .A2(I525), .ZN(W262));
  NOR2X1 G11828 (.A1(W8963), .A2(W2999), .ZN(O3345));
  NOR2X1 G11829 (.A1(W23126), .A2(W5906), .ZN(W25254));
  NOR2X1 G11830 (.A1(W16655), .A2(W20431), .ZN(O19505));
  NOR2X1 G11831 (.A1(I494), .A2(I495), .ZN(W247));
  NOR2X1 G11832 (.A1(I492), .A2(I493), .ZN(W246));
  NOR2X1 G11833 (.A1(W586), .A2(W19439), .ZN(W25257));
  NOR2X1 G11834 (.A1(I484), .A2(I485), .ZN(W242));
  NOR2X1 G11835 (.A1(I540), .A2(I541), .ZN(W270));
  NOR2X1 G11836 (.A1(I558), .A2(I559), .ZN(W279));
  NOR2X1 G11837 (.A1(I556), .A2(I557), .ZN(W278));
  NOR2X1 G11838 (.A1(I554), .A2(I555), .ZN(W277));
  NOR2X1 G11839 (.A1(W49942), .A2(W5099), .ZN(O19484));
  NOR2X1 G11840 (.A1(I550), .A2(I551), .ZN(W275));
  NOR2X1 G11841 (.A1(I548), .A2(I549), .ZN(W274));
  NOR2X1 G11842 (.A1(I546), .A2(I547), .ZN(W273));
  NOR2X1 G11843 (.A1(W6578), .A2(W26593), .ZN(O19485));
  NOR2X1 G11844 (.A1(I316), .A2(I317), .ZN(W158));
  NOR2X1 G11845 (.A1(I538), .A2(I539), .ZN(W269));
  NOR2X1 G11846 (.A1(W23696), .A2(W3303), .ZN(W25440));
  NOR2X1 G11847 (.A1(W5227), .A2(W47518), .ZN(O19488));
  NOR2X1 G11848 (.A1(W19157), .A2(I893), .ZN(W25248));
  NOR2X1 G11849 (.A1(I530), .A2(I531), .ZN(W265));
  NOR2X1 G11850 (.A1(W11113), .A2(W2666), .ZN(O19490));
  NOR2X1 G11851 (.A1(I526), .A2(I527), .ZN(W263));
  NOR2X1 G11852 (.A1(W9204), .A2(W33446), .ZN(O19705));
  NOR2X1 G11853 (.A1(I120), .A2(I121), .ZN(W60));
  NOR2X1 G11854 (.A1(W13563), .A2(W9143), .ZN(W25324));
  NOR2X1 G11855 (.A1(I114), .A2(I115), .ZN(W57));
  NOR2X1 G11856 (.A1(I112), .A2(I113), .ZN(W56));
  NOR2X1 G11857 (.A1(I110), .A2(I111), .ZN(W55));
  NOR2X1 G11858 (.A1(W22489), .A2(W16582), .ZN(W25325));
  NOR2X1 G11859 (.A1(W17376), .A2(W615), .ZN(O19703));
  NOR2X1 G11860 (.A1(W43645), .A2(W24544), .ZN(O19704));
  NOR2X1 G11861 (.A1(I122), .A2(I123), .ZN(W61));
  NOR2X1 G11862 (.A1(W25262), .A2(W20777), .ZN(O3392));
  NOR2X1 G11863 (.A1(W1223), .A2(W38454), .ZN(O19710));
  NOR2X1 G11864 (.A1(W3539), .A2(W23264), .ZN(O3391));
  NOR2X1 G11865 (.A1(W36648), .A2(W892), .ZN(O19712));
  NOR2X1 G11866 (.A1(W31566), .A2(W26004), .ZN(O19713));
  NOR2X1 G11867 (.A1(I90), .A2(I91), .ZN(W45));
  NOR2X1 G11868 (.A1(W19353), .A2(W20710), .ZN(O19714));
  NOR2X1 G11869 (.A1(W12589), .A2(W32866), .ZN(O19716));
  NOR2X1 G11870 (.A1(W22635), .A2(W1024), .ZN(W25370));
  NOR2X1 G11871 (.A1(W6575), .A2(W22631), .ZN(W25316));
  NOR2X1 G11872 (.A1(W19720), .A2(W42320), .ZN(O19670));
  NOR2X1 G11873 (.A1(I152), .A2(I153), .ZN(W76));
  NOR2X1 G11874 (.A1(I150), .A2(I151), .ZN(W75));
  NOR2X1 G11875 (.A1(W26038), .A2(W25731), .ZN(O19673));
  NOR2X1 G11876 (.A1(I146), .A2(I147), .ZN(W73));
  NOR2X1 G11877 (.A1(W8775), .A2(W23978), .ZN(O19674));
  NOR2X1 G11878 (.A1(W18443), .A2(W10932), .ZN(O19675));
  NOR2X1 G11879 (.A1(W8562), .A2(W22407), .ZN(O19719));
  NOR2X1 G11880 (.A1(W17603), .A2(W30560), .ZN(O19681));
  NOR2X1 G11881 (.A1(W14817), .A2(W37755), .ZN(O19682));
  NOR2X1 G11882 (.A1(W7894), .A2(W33325), .ZN(O19683));
  NOR2X1 G11883 (.A1(W9857), .A2(W24483), .ZN(W25368));
  NOR2X1 G11884 (.A1(W11580), .A2(W14288), .ZN(W25321));
  NOR2X1 G11885 (.A1(I1783), .A2(W16514), .ZN(O19688));
  NOR2X1 G11886 (.A1(W592), .A2(I1202), .ZN(O3374));
  NOR2X1 G11887 (.A1(I20), .A2(I21), .ZN(W10));
  NOR2X1 G11888 (.A1(I42), .A2(I43), .ZN(W21));
  NOR2X1 G11889 (.A1(W20799), .A2(W24542), .ZN(W25350));
  NOR2X1 G11890 (.A1(W18928), .A2(W18230), .ZN(O3384));
  NOR2X1 G11891 (.A1(I30), .A2(I31), .ZN(W15));
  NOR2X1 G11892 (.A1(W32064), .A2(I721), .ZN(O19748));
  NOR2X1 G11893 (.A1(I26), .A2(I27), .ZN(W13));
  NOR2X1 G11894 (.A1(W16977), .A2(W22642), .ZN(O3382));
  NOR2X1 G11895 (.A1(W17265), .A2(W47027), .ZN(O19752));
  NOR2X1 G11896 (.A1(W21608), .A2(I376), .ZN(O3386));
  NOR2X1 G11897 (.A1(W31414), .A2(W29558), .ZN(O19753));
  NOR2X1 G11898 (.A1(W21328), .A2(W46985), .ZN(O19754));
  NOR2X1 G11899 (.A1(I10), .A2(I11), .ZN(W5));
  NOR2X1 G11900 (.A1(I8), .A2(I9), .ZN(W4));
  NOR2X1 G11901 (.A1(I6), .A2(I7), .ZN(W3));
  NOR2X1 G11902 (.A1(W20140), .A2(W9887), .ZN(O19759));
  NOR2X1 G11903 (.A1(W11680), .A2(I615), .ZN(W25343));
  NOR2X1 G11904 (.A1(I64), .A2(I65), .ZN(W32));
  NOR2X1 G11905 (.A1(I80), .A2(I81), .ZN(W40));
  NOR2X1 G11906 (.A1(I78), .A2(I79), .ZN(W39));
  NOR2X1 G11907 (.A1(W8617), .A2(W24908), .ZN(O19721));
  NOR2X1 G11908 (.A1(I74), .A2(I75), .ZN(W37));
  NOR2X1 G11909 (.A1(W10305), .A2(W43681), .ZN(O19722));
  NOR2X1 G11910 (.A1(I70), .A2(I71), .ZN(W35));
  NOR2X1 G11911 (.A1(W32089), .A2(W5269), .ZN(O19724));
  NOR2X1 G11912 (.A1(W9815), .A2(W49007), .ZN(O19726));
  NOR2X1 G11913 (.A1(I160), .A2(I161), .ZN(W80));
  NOR2X1 G11914 (.A1(W5528), .A2(W17202), .ZN(O3388));
  NOR2X1 G11915 (.A1(W1643), .A2(W11990), .ZN(W25330));
  NOR2X1 G11916 (.A1(W5654), .A2(W39785), .ZN(O19731));
  NOR2X1 G11917 (.A1(I56), .A2(I57), .ZN(W28));
  NOR2X1 G11918 (.A1(I50), .A2(I51), .ZN(W25));
  NOR2X1 G11919 (.A1(I48), .A2(I49), .ZN(W24));
  NOR2X1 G11920 (.A1(W49234), .A2(W32042), .ZN(O19737));
  NOR2X1 G11921 (.A1(W6423), .A2(W728), .ZN(W25305));
  NOR2X1 G11922 (.A1(I270), .A2(I271), .ZN(W135));
  NOR2X1 G11923 (.A1(I266), .A2(I267), .ZN(W133));
  NOR2X1 G11924 (.A1(I262), .A2(I263), .ZN(W131));
  NOR2X1 G11925 (.A1(I260), .A2(I261), .ZN(W130));
  NOR2X1 G11926 (.A1(W42854), .A2(W33609), .ZN(O19631));
  NOR2X1 G11927 (.A1(I256), .A2(I257), .ZN(W128));
  NOR2X1 G11928 (.A1(W49538), .A2(W26129), .ZN(O19632));
  NOR2X1 G11929 (.A1(I252), .A2(I253), .ZN(W126));
  NOR2X1 G11930 (.A1(W3266), .A2(W23361), .ZN(O3366));
  NOR2X1 G11931 (.A1(I248), .A2(I249), .ZN(W124));
  NOR2X1 G11932 (.A1(I246), .A2(I247), .ZN(W123));
  NOR2X1 G11933 (.A1(I244), .A2(I245), .ZN(W122));
  NOR2X1 G11934 (.A1(W2868), .A2(W4844), .ZN(W25306));
  NOR2X1 G11935 (.A1(I240), .A2(I241), .ZN(W120));
  NOR2X1 G11936 (.A1(W4105), .A2(W20465), .ZN(O3368));
  NOR2X1 G11937 (.A1(W12254), .A2(W10521), .ZN(O19637));
  NOR2X1 G11938 (.A1(I234), .A2(I235), .ZN(W117));
  NOR2X1 G11939 (.A1(W2012), .A2(W17063), .ZN(O19609));
  NOR2X1 G11940 (.A1(W3463), .A2(W20296), .ZN(O3403));
  NOR2X1 G11941 (.A1(W29188), .A2(W45751), .ZN(O19600));
  NOR2X1 G11942 (.A1(W34237), .A2(W48569), .ZN(O19601));
  NOR2X1 G11943 (.A1(W3286), .A2(W7782), .ZN(O3402));
  NOR2X1 G11944 (.A1(W18243), .A2(W5904), .ZN(O3362));
  NOR2X1 G11945 (.A1(W27444), .A2(W8971), .ZN(O19605));
  NOR2X1 G11946 (.A1(W8153), .A2(W48106), .ZN(O19607));
  NOR2X1 G11947 (.A1(W6567), .A2(W1883), .ZN(O19608));
  NOR2X1 G11948 (.A1(W11633), .A2(W18300), .ZN(O3395));
  NOR2X1 G11949 (.A1(W9321), .A2(W14437), .ZN(O19611));
  NOR2X1 G11950 (.A1(W6646), .A2(W33645), .ZN(O19613));
  NOR2X1 G11951 (.A1(W2023), .A2(W15944), .ZN(O19614));
  NOR2X1 G11952 (.A1(W8839), .A2(W9994), .ZN(W25298));
  NOR2X1 G11953 (.A1(I282), .A2(I283), .ZN(W141));
  NOR2X1 G11954 (.A1(W6373), .A2(W49966), .ZN(O19618));
  NOR2X1 G11955 (.A1(W39432), .A2(W16974), .ZN(O19621));
  NOR2X1 G11956 (.A1(I178), .A2(I179), .ZN(W89));
  NOR2X1 G11957 (.A1(W18288), .A2(W23007), .ZN(O19654));
  NOR2X1 G11958 (.A1(W23164), .A2(I657), .ZN(W25312));
  NOR2X1 G11959 (.A1(I192), .A2(I193), .ZN(W96));
  NOR2X1 G11960 (.A1(I190), .A2(I191), .ZN(W95));
  NOR2X1 G11961 (.A1(W14493), .A2(W49068), .ZN(O19657));
  NOR2X1 G11962 (.A1(I184), .A2(I185), .ZN(W92));
  NOR2X1 G11963 (.A1(I1141), .A2(W14678), .ZN(O19659));
  NOR2X1 G11964 (.A1(I180), .A2(I181), .ZN(W90));
  NOR2X1 G11965 (.A1(W14223), .A2(W8578), .ZN(W25376));
  NOR2X1 G11966 (.A1(W45437), .A2(W44154), .ZN(O19661));
  NOR2X1 G11967 (.A1(I174), .A2(I175), .ZN(W87));
  NOR2X1 G11968 (.A1(I170), .A2(I171), .ZN(W85));
  NOR2X1 G11969 (.A1(I168), .A2(I169), .ZN(W84));
  NOR2X1 G11970 (.A1(W44949), .A2(W28817), .ZN(O19666));
  NOR2X1 G11971 (.A1(W2553), .A2(W13214), .ZN(W25372));
  NOR2X1 G11972 (.A1(I162), .A2(I163), .ZN(W81));
  NOR2X1 G11973 (.A1(W4663), .A2(W18948), .ZN(W25309));
  NOR2X1 G11974 (.A1(I230), .A2(I231), .ZN(W115));
  NOR2X1 G11975 (.A1(W24748), .A2(W12809), .ZN(O19640));
  NOR2X1 G11976 (.A1(W24907), .A2(W41305), .ZN(O19641));
  NOR2X1 G11977 (.A1(I224), .A2(I225), .ZN(W112));
  NOR2X1 G11978 (.A1(W36396), .A2(W7984), .ZN(O19642));
  NOR2X1 G11979 (.A1(W41699), .A2(W26415), .ZN(O19643));
  NOR2X1 G11980 (.A1(I218), .A2(I219), .ZN(W109));
  NOR2X1 G11981 (.A1(I216), .A2(I217), .ZN(W108));
  NOR2X1 G11982 (.A1(I640), .A2(I641), .ZN(W320));
  NOR2X1 G11983 (.A1(W15865), .A2(W26164), .ZN(O19646));
  NOR2X1 G11984 (.A1(W12614), .A2(W5442), .ZN(W25310));
  NOR2X1 G11985 (.A1(W2209), .A2(W35335), .ZN(O19648));
  NOR2X1 G11986 (.A1(W8031), .A2(W48663), .ZN(O19649));
  NOR2X1 G11987 (.A1(I1646), .A2(W22381), .ZN(O19650));
  NOR2X1 G11988 (.A1(W50627), .A2(W39695), .ZN(O19651));
  NOR2X1 G11989 (.A1(W44501), .A2(W29406), .ZN(O19652));
  NOR2X1 G11990 (.A1(I1048), .A2(I1049), .ZN(W524));
  NOR2X1 G11991 (.A1(W23682), .A2(W19008), .ZN(O19238));
  NOR2X1 G11992 (.A1(I1066), .A2(I1067), .ZN(W533));
  NOR2X1 G11993 (.A1(I1064), .A2(I1065), .ZN(W532));
  NOR2X1 G11994 (.A1(W20289), .A2(W9593), .ZN(O3320));
  NOR2X1 G11995 (.A1(W11653), .A2(W25437), .ZN(O3444));
  NOR2X1 G11996 (.A1(W3044), .A2(W34088), .ZN(O19246));
  NOR2X1 G11997 (.A1(W44307), .A2(W13279), .ZN(O19247));
  NOR2X1 G11998 (.A1(I619), .A2(W16866), .ZN(O19248));
  NOR2X1 G11999 (.A1(W11597), .A2(W132), .ZN(O3319));
  NOR2X1 G12000 (.A1(W2392), .A2(W22217), .ZN(O19252));
  NOR2X1 G12001 (.A1(W23163), .A2(W28270), .ZN(O19255));
  NOR2X1 G12002 (.A1(W46834), .A2(W14556), .ZN(O19260));
  NOR2X1 G12003 (.A1(W23569), .A2(W44594), .ZN(O19262));
  NOR2X1 G12004 (.A1(I1032), .A2(I1033), .ZN(W516));
  NOR2X1 G12005 (.A1(I1030), .A2(I1031), .ZN(W515));
  NOR2X1 G12006 (.A1(I1028), .A2(I1029), .ZN(W514));
  NOR2X1 G12007 (.A1(W32859), .A2(W34373), .ZN(O19263));
  NOR2X1 G12008 (.A1(W1494), .A2(W9676), .ZN(W25167));
  NOR2X1 G12009 (.A1(I1104), .A2(I1105), .ZN(W552));
  NOR2X1 G12010 (.A1(W32015), .A2(W27063), .ZN(O19222));
  NOR2X1 G12011 (.A1(W22081), .A2(W4855), .ZN(W25527));
  NOR2X1 G12012 (.A1(W5141), .A2(W37889), .ZN(O19225));
  NOR2X1 G12013 (.A1(W33061), .A2(I1694), .ZN(O19226));
  NOR2X1 G12014 (.A1(I1094), .A2(I1095), .ZN(W547));
  NOR2X1 G12015 (.A1(W39039), .A2(W16147), .ZN(O19227));
  NOR2X1 G12016 (.A1(I1090), .A2(I1091), .ZN(W545));
  NOR2X1 G12017 (.A1(I1024), .A2(I1025), .ZN(W512));
  NOR2X1 G12018 (.A1(W18730), .A2(W254), .ZN(W25526));
  NOR2X1 G12019 (.A1(W28909), .A2(W12726), .ZN(O19232));
  NOR2X1 G12020 (.A1(W29833), .A2(W1692), .ZN(O19233));
  NOR2X1 G12021 (.A1(W35954), .A2(W10429), .ZN(O19234));
  NOR2X1 G12022 (.A1(I1078), .A2(I1079), .ZN(W539));
  NOR2X1 G12023 (.A1(W16481), .A2(W7350), .ZN(W25169));
  NOR2X1 G12024 (.A1(I1072), .A2(I1073), .ZN(W536));
  NOR2X1 G12025 (.A1(I968), .A2(I969), .ZN(W484));
  NOR2X1 G12026 (.A1(W17677), .A2(W4414), .ZN(W25183));
  NOR2X1 G12027 (.A1(I982), .A2(I983), .ZN(W491));
  NOR2X1 G12028 (.A1(W33531), .A2(W28673), .ZN(O19281));
  NOR2X1 G12029 (.A1(W37923), .A2(W25388), .ZN(O19282));
  NOR2X1 G12030 (.A1(W3032), .A2(W4423), .ZN(O19283));
  NOR2X1 G12031 (.A1(I974), .A2(I975), .ZN(W487));
  NOR2X1 G12032 (.A1(W11228), .A2(W33912), .ZN(O19285));
  NOR2X1 G12033 (.A1(W19937), .A2(W16332), .ZN(W25184));
  NOR2X1 G12034 (.A1(W17496), .A2(W24460), .ZN(O19279));
  NOR2X1 G12035 (.A1(W9379), .A2(I736), .ZN(W25506));
  NOR2X1 G12036 (.A1(W21688), .A2(W1729), .ZN(O19293));
  NOR2X1 G12037 (.A1(W27596), .A2(W1316), .ZN(O19297));
  NOR2X1 G12038 (.A1(I956), .A2(I957), .ZN(W478));
  NOR2X1 G12039 (.A1(W42599), .A2(W12630), .ZN(O19298));
  NOR2X1 G12040 (.A1(W7907), .A2(W24892), .ZN(W25504));
  NOR2X1 G12041 (.A1(W18729), .A2(W19498), .ZN(W25503));
  NOR2X1 G12042 (.A1(W11460), .A2(W12710), .ZN(W25180));
  NOR2X1 G12043 (.A1(W30965), .A2(W3487), .ZN(O19265));
  NOR2X1 G12044 (.A1(I1020), .A2(I1021), .ZN(W510));
  NOR2X1 G12045 (.A1(W26675), .A2(W22906), .ZN(O19266));
  NOR2X1 G12046 (.A1(W31724), .A2(W44995), .ZN(O19267));
  NOR2X1 G12047 (.A1(I1014), .A2(I1015), .ZN(W507));
  NOR2X1 G12048 (.A1(I1010), .A2(I1011), .ZN(W505));
  NOR2X1 G12049 (.A1(W32266), .A2(W2855), .ZN(O19269));
  NOR2X1 G12050 (.A1(W39587), .A2(W39790), .ZN(O19270));
  NOR2X1 G12051 (.A1(I1106), .A2(I1107), .ZN(W553));
  NOR2X1 G12052 (.A1(W20059), .A2(W15803), .ZN(O19274));
  NOR2X1 G12053 (.A1(I1000), .A2(I1001), .ZN(W500));
  NOR2X1 G12054 (.A1(I998), .A2(I999), .ZN(W499));
  NOR2X1 G12055 (.A1(W11722), .A2(W22083), .ZN(W25508));
  NOR2X1 G12056 (.A1(W49341), .A2(W41926), .ZN(O19278));
  NOR2X1 G12057 (.A1(I990), .A2(I991), .ZN(W495));
  NOR2X1 G12058 (.A1(I988), .A2(I989), .ZN(W494));
  NOR2X1 G12059 (.A1(W5695), .A2(W23215), .ZN(W25538));
  NOR2X1 G12060 (.A1(I1220), .A2(I1221), .ZN(W610));
  NOR2X1 G12061 (.A1(W35207), .A2(W26559), .ZN(O19167));
  NOR2X1 G12062 (.A1(W38828), .A2(W11646), .ZN(O19169));
  NOR2X1 G12063 (.A1(W15851), .A2(W28182), .ZN(O19170));
  NOR2X1 G12064 (.A1(I1212), .A2(I1213), .ZN(W606));
  NOR2X1 G12065 (.A1(I1210), .A2(I1211), .ZN(W605));
  NOR2X1 G12066 (.A1(W7986), .A2(W23076), .ZN(W25540));
  NOR2X1 G12067 (.A1(W7846), .A2(W23435), .ZN(W25148));
  NOR2X1 G12068 (.A1(I1224), .A2(I1225), .ZN(W612));
  NOR2X1 G12069 (.A1(W9352), .A2(W20328), .ZN(W25152));
  NOR2X1 G12070 (.A1(W22041), .A2(W11140), .ZN(O19179));
  NOR2X1 G12071 (.A1(I1194), .A2(I1195), .ZN(W597));
  NOR2X1 G12072 (.A1(W6939), .A2(W10244), .ZN(W25153));
  NOR2X1 G12073 (.A1(W27010), .A2(W39215), .ZN(O19181));
  NOR2X1 G12074 (.A1(W7679), .A2(W2354), .ZN(O19183));
  NOR2X1 G12075 (.A1(W3122), .A2(W39906), .ZN(O19189));
  NOR2X1 G12076 (.A1(W18360), .A2(W2840), .ZN(O19194));
  NOR2X1 G12077 (.A1(W29900), .A2(W10913), .ZN(O19162));
  NOR2X1 G12078 (.A1(W39235), .A2(W13639), .ZN(O19158));
  NOR2X1 G12079 (.A1(W22057), .A2(W9371), .ZN(W25143));
  NOR2X1 G12080 (.A1(I1254), .A2(I1255), .ZN(W627));
  NOR2X1 G12081 (.A1(I1252), .A2(I1253), .ZN(W626));
  NOR2X1 G12082 (.A1(W49437), .A2(W32434), .ZN(O19161));
  NOR2X1 G12083 (.A1(I1246), .A2(I1247), .ZN(W623));
  NOR2X1 G12084 (.A1(I1244), .A2(I1245), .ZN(W622));
  NOR2X1 G12085 (.A1(I1242), .A2(I1243), .ZN(W621));
  NOR2X1 G12086 (.A1(W39394), .A2(W5748), .ZN(O19196));
  NOR2X1 G12087 (.A1(I1238), .A2(I1239), .ZN(W619));
  NOR2X1 G12088 (.A1(W23737), .A2(W12724), .ZN(O3451));
  NOR2X1 G12089 (.A1(I1234), .A2(I1235), .ZN(W617));
  NOR2X1 G12090 (.A1(I1232), .A2(I1233), .ZN(W616));
  NOR2X1 G12091 (.A1(I1230), .A2(I1231), .ZN(W615));
  NOR2X1 G12092 (.A1(I1228), .A2(I1229), .ZN(W614));
  NOR2X1 G12093 (.A1(W18088), .A2(W39987), .ZN(O19164));
  NOR2X1 G12094 (.A1(I1122), .A2(I1123), .ZN(W561));
  NOR2X1 G12095 (.A1(I1138), .A2(I1139), .ZN(W569));
  NOR2X1 G12096 (.A1(W3859), .A2(W1227), .ZN(W25162));
  NOR2X1 G12097 (.A1(W23237), .A2(W49816), .ZN(W50445));
  NOR2X1 G12098 (.A1(W6756), .A2(W31570), .ZN(O19212));
  NOR2X1 G12099 (.A1(W21884), .A2(W18321), .ZN(W25529));
  NOR2X1 G12100 (.A1(W37611), .A2(W35022), .ZN(O19214));
  NOR2X1 G12101 (.A1(I1126), .A2(I1127), .ZN(W563));
  NOR2X1 G12102 (.A1(W38143), .A2(W25967), .ZN(O19215));
  NOR2X1 G12103 (.A1(W13225), .A2(W22386), .ZN(O19208));
  NOR2X1 G12104 (.A1(I1120), .A2(I1121), .ZN(W560));
  NOR2X1 G12105 (.A1(I1118), .A2(I1119), .ZN(W559));
  NOR2X1 G12106 (.A1(W25746), .A2(W42499), .ZN(O19217));
  NOR2X1 G12107 (.A1(W2146), .A2(W15561), .ZN(W25528));
  NOR2X1 G12108 (.A1(W21023), .A2(W6011), .ZN(W25165));
  NOR2X1 G12109 (.A1(I1110), .A2(I1111), .ZN(W555));
  NOR2X1 G12110 (.A1(W49774), .A2(W36317), .ZN(O19221));
  NOR2X1 G12111 (.A1(I1160), .A2(I1161), .ZN(W580));
  NOR2X1 G12112 (.A1(W40335), .A2(W13919), .ZN(O19197));
  NOR2X1 G12113 (.A1(W14628), .A2(W15001), .ZN(W25156));
  NOR2X1 G12114 (.A1(I1172), .A2(I1173), .ZN(W586));
  NOR2X1 G12115 (.A1(I1170), .A2(I1171), .ZN(W585));
  NOR2X1 G12116 (.A1(I1806), .A2(W13805), .ZN(O3448));
  NOR2X1 G12117 (.A1(I1166), .A2(I1167), .ZN(W583));
  NOR2X1 G12118 (.A1(I1164), .A2(I1165), .ZN(W582));
  NOR2X1 G12119 (.A1(I1162), .A2(I1163), .ZN(W581));
  NOR2X1 G12120 (.A1(W11466), .A2(W4300), .ZN(O3325));
  NOR2X1 G12121 (.A1(W35874), .A2(W41300), .ZN(O19201));
  NOR2X1 G12122 (.A1(W8540), .A2(W18675), .ZN(W25159));
  NOR2X1 G12123 (.A1(W10757), .A2(W14140), .ZN(W50437));
  NOR2X1 G12124 (.A1(I1150), .A2(I1151), .ZN(W575));
  NOR2X1 G12125 (.A1(I1148), .A2(I1149), .ZN(W574));
  NOR2X1 G12126 (.A1(I1144), .A2(I1145), .ZN(W572));
  NOR2X1 G12127 (.A1(W23083), .A2(W19413), .ZN(O3317));
  NOR2X1 G12128 (.A1(I736), .A2(I737), .ZN(W368));
  NOR2X1 G12129 (.A1(W20760), .A2(W22725), .ZN(W25218));
  NOR2X1 G12130 (.A1(W47309), .A2(W4878), .ZN(O19389));
  NOR2X1 G12131 (.A1(I752), .A2(I753), .ZN(W376));
  NOR2X1 G12132 (.A1(W42299), .A2(W20582), .ZN(O19390));
  NOR2X1 G12133 (.A1(I744), .A2(I745), .ZN(W372));
  NOR2X1 G12134 (.A1(W42317), .A2(W41587), .ZN(O19399));
  NOR2X1 G12135 (.A1(W2749), .A2(W15649), .ZN(O3333));
  NOR2X1 G12136 (.A1(W31384), .A2(I96), .ZN(O19402));
  NOR2X1 G12137 (.A1(W22129), .A2(W17809), .ZN(W25217));
  NOR2X1 G12138 (.A1(W49237), .A2(W40905), .ZN(O19403));
  NOR2X1 G12139 (.A1(W7370), .A2(W16123), .ZN(W25222));
  NOR2X1 G12140 (.A1(I730), .A2(I731), .ZN(W365));
  NOR2X1 G12141 (.A1(I728), .A2(I729), .ZN(W364));
  NOR2X1 G12142 (.A1(I726), .A2(I727), .ZN(W363));
  NOR2X1 G12143 (.A1(I724), .A2(I725), .ZN(W362));
  NOR2X1 G12144 (.A1(I722), .A2(I723), .ZN(W361));
  NOR2X1 G12145 (.A1(W31753), .A2(W17173), .ZN(O19405));
  NOR2X1 G12146 (.A1(W48478), .A2(W47372), .ZN(O19377));
  NOR2X1 G12147 (.A1(I792), .A2(I793), .ZN(W396));
  NOR2X1 G12148 (.A1(I790), .A2(I791), .ZN(W395));
  NOR2X1 G12149 (.A1(I786), .A2(I787), .ZN(W393));
  NOR2X1 G12150 (.A1(I784), .A2(I785), .ZN(W392));
  NOR2X1 G12151 (.A1(W3686), .A2(W23422), .ZN(W25474));
  NOR2X1 G12152 (.A1(I780), .A2(I781), .ZN(W390));
  NOR2X1 G12153 (.A1(I778), .A2(I779), .ZN(W389));
  NOR2X1 G12154 (.A1(I776), .A2(I777), .ZN(W388));
  NOR2X1 G12155 (.A1(W1619), .A2(W13661), .ZN(W25223));
  NOR2X1 G12156 (.A1(W6063), .A2(W10548), .ZN(O3331));
  NOR2X1 G12157 (.A1(W40303), .A2(W36988), .ZN(O19379));
  NOR2X1 G12158 (.A1(W45558), .A2(I1446), .ZN(O19380));
  NOR2X1 G12159 (.A1(I766), .A2(I767), .ZN(W383));
  NOR2X1 G12160 (.A1(I764), .A2(I765), .ZN(W382));
  NOR2X1 G12161 (.A1(I842), .A2(W11883), .ZN(W25216));
  NOR2X1 G12162 (.A1(W11218), .A2(W37351), .ZN(O19383));
  NOR2X1 G12163 (.A1(W20753), .A2(W6753), .ZN(W25233));
  NOR2X1 G12164 (.A1(I678), .A2(I679), .ZN(W339));
  NOR2X1 G12165 (.A1(I676), .A2(I677), .ZN(W338));
  NOR2X1 G12166 (.A1(I674), .A2(I675), .ZN(W337));
  NOR2X1 G12167 (.A1(I672), .A2(I673), .ZN(O4));
  NOR2X1 G12168 (.A1(I670), .A2(I671), .ZN(W335));
  NOR2X1 G12169 (.A1(I668), .A2(I669), .ZN(W334));
  NOR2X1 G12170 (.A1(W40813), .A2(W14779), .ZN(O19428));
  NOR2X1 G12171 (.A1(W37448), .A2(W46372), .ZN(O19429));
  NOR2X1 G12172 (.A1(I680), .A2(I681), .ZN(W340));
  NOR2X1 G12173 (.A1(I658), .A2(I659), .ZN(W329));
  NOR2X1 G12174 (.A1(W44587), .A2(W29258), .ZN(O19433));
  NOR2X1 G12175 (.A1(W21727), .A2(W4434), .ZN(O19434));
  NOR2X1 G12176 (.A1(W16376), .A2(W16843), .ZN(O19435));
  NOR2X1 G12177 (.A1(I648), .A2(I649), .ZN(W324));
  NOR2X1 G12178 (.A1(I646), .A2(I647), .ZN(W323));
  NOR2X1 G12179 (.A1(W27638), .A2(W14302), .ZN(O19438));
  NOR2X1 G12180 (.A1(I700), .A2(I701), .ZN(W350));
  NOR2X1 G12181 (.A1(W40215), .A2(W172), .ZN(O19408));
  NOR2X1 G12182 (.A1(W13622), .A2(W13517), .ZN(W25470));
  NOR2X1 G12183 (.A1(I712), .A2(I713), .ZN(W356));
  NOR2X1 G12184 (.A1(I710), .A2(I711), .ZN(W355));
  NOR2X1 G12185 (.A1(W5855), .A2(W6398), .ZN(W25469));
  NOR2X1 G12186 (.A1(I706), .A2(I707), .ZN(W353));
  NOR2X1 G12187 (.A1(W23153), .A2(W25177), .ZN(O3335));
  NOR2X1 G12188 (.A1(W19598), .A2(I49), .ZN(O3336));
  NOR2X1 G12189 (.A1(W65), .A2(W16041), .ZN(O19371));
  NOR2X1 G12190 (.A1(W14076), .A2(W38656), .ZN(O19418));
  NOR2X1 G12191 (.A1(I694), .A2(I695), .ZN(W347));
  NOR2X1 G12192 (.A1(W23484), .A2(W25673), .ZN(O19419));
  NOR2X1 G12193 (.A1(W23677), .A2(I1746), .ZN(W25465));
  NOR2X1 G12194 (.A1(W12300), .A2(W7085), .ZN(W25464));
  NOR2X1 G12195 (.A1(W17489), .A2(W46518), .ZN(O19424));
  NOR2X1 G12196 (.A1(I682), .A2(I683), .ZN(W341));
  NOR2X1 G12197 (.A1(I894), .A2(I895), .ZN(W447));
  NOR2X1 G12198 (.A1(I910), .A2(I911), .ZN(W455));
  NOR2X1 G12199 (.A1(I908), .A2(I909), .ZN(W454));
  NOR2X1 G12200 (.A1(W838), .A2(W764), .ZN(W25194));
  NOR2X1 G12201 (.A1(W47239), .A2(W45920), .ZN(O19317));
  NOR2X1 G12202 (.A1(I514), .A2(W13833), .ZN(W25195));
  NOR2X1 G12203 (.A1(W37950), .A2(W8589), .ZN(O19319));
  NOR2X1 G12204 (.A1(W18900), .A2(W12539), .ZN(O19320));
  NOR2X1 G12205 (.A1(W29883), .A2(W13904), .ZN(O19321));
  NOR2X1 G12206 (.A1(I912), .A2(I913), .ZN(W456));
  NOR2X1 G12207 (.A1(W17720), .A2(W2381), .ZN(O3327));
  NOR2X1 G12208 (.A1(I888), .A2(I889), .ZN(W444));
  NOR2X1 G12209 (.A1(I884), .A2(I885), .ZN(W442));
  NOR2X1 G12210 (.A1(W13020), .A2(W16004), .ZN(O19325));
  NOR2X1 G12211 (.A1(I880), .A2(I881), .ZN(W440));
  NOR2X1 G12212 (.A1(W28964), .A2(W15557), .ZN(O19327));
  NOR2X1 G12213 (.A1(W2455), .A2(W6570), .ZN(W25495));
  NOR2X1 G12214 (.A1(I874), .A2(I875), .ZN(W437));
  NOR2X1 G12215 (.A1(I928), .A2(I929), .ZN(W464));
  NOR2X1 G12216 (.A1(W3741), .A2(W27311), .ZN(O19303));
  NOR2X1 G12217 (.A1(I942), .A2(I943), .ZN(W471));
  NOR2X1 G12218 (.A1(W24876), .A2(W19756), .ZN(O3437));
  NOR2X1 G12219 (.A1(W45855), .A2(W4551), .ZN(O19305));
  NOR2X1 G12220 (.A1(I936), .A2(I937), .ZN(W468));
  NOR2X1 G12221 (.A1(W28579), .A2(W26999), .ZN(O19306));
  NOR2X1 G12222 (.A1(W19812), .A2(W9764), .ZN(O19307));
  NOR2X1 G12223 (.A1(W29483), .A2(W18561), .ZN(O19311));
  NOR2X1 G12224 (.A1(W7611), .A2(W14401), .ZN(O19331));
  NOR2X1 G12225 (.A1(W21040), .A2(W9915), .ZN(W25499));
  NOR2X1 G12226 (.A1(I924), .A2(I925), .ZN(W462));
  NOR2X1 G12227 (.A1(I922), .A2(I923), .ZN(W461));
  NOR2X1 G12228 (.A1(W48022), .A2(W48705), .ZN(O19313));
  NOR2X1 G12229 (.A1(W14342), .A2(W50242), .ZN(O19314));
  NOR2X1 G12230 (.A1(I916), .A2(I917), .ZN(W458));
  NOR2X1 G12231 (.A1(I914), .A2(I915), .ZN(W457));
  NOR2X1 G12232 (.A1(I816), .A2(I817), .ZN(W408));
  NOR2X1 G12233 (.A1(W6100), .A2(W9061), .ZN(W25203));
  NOR2X1 G12234 (.A1(I832), .A2(I833), .ZN(W416));
  NOR2X1 G12235 (.A1(I830), .A2(I831), .ZN(W415));
  NOR2X1 G12236 (.A1(W6681), .A2(W1824), .ZN(W25204));
  NOR2X1 G12237 (.A1(I614), .A2(W24075), .ZN(W25488));
  NOR2X1 G12238 (.A1(I824), .A2(I825), .ZN(W412));
  NOR2X1 G12239 (.A1(W9764), .A2(W31850), .ZN(O19353));
  NOR2X1 G12240 (.A1(I818), .A2(I819), .ZN(W409));
  NOR2X1 G12241 (.A1(W684), .A2(W19536), .ZN(W25490));
  NOR2X1 G12242 (.A1(I814), .A2(I815), .ZN(W407));
  NOR2X1 G12243 (.A1(W14267), .A2(W28793), .ZN(O19356));
  NOR2X1 G12244 (.A1(W19457), .A2(W1273), .ZN(W25485));
  NOR2X1 G12245 (.A1(I808), .A2(I809), .ZN(W404));
  NOR2X1 G12246 (.A1(W21422), .A2(W6921), .ZN(O3433));
  NOR2X1 G12247 (.A1(W22195), .A2(W18097), .ZN(W25479));
  NOR2X1 G12248 (.A1(I1466), .A2(W7199), .ZN(O19368));
  NOR2X1 G12249 (.A1(W15186), .A2(W50539), .ZN(O19338));
  NOR2X1 G12250 (.A1(I870), .A2(I871), .ZN(W435));
  NOR2X1 G12251 (.A1(W48469), .A2(W48553), .ZN(O19333));
  NOR2X1 G12252 (.A1(W21171), .A2(W4140), .ZN(O19335));
  NOR2X1 G12253 (.A1(W9904), .A2(W27569), .ZN(O19337));
  NOR2X1 G12254 (.A1(I862), .A2(I863), .ZN(W431));
  NOR2X1 G12255 (.A1(I860), .A2(I861), .ZN(W430));
  NOR2X1 G12256 (.A1(I858), .A2(I859), .ZN(W429));
  NOR2X1 G12257 (.A1(I856), .A2(I857), .ZN(W428));
  NOR2X1 G12258 (.A1(I646), .A2(I983), .ZN(W1257));
  NOR2X1 G12259 (.A1(I852), .A2(I853), .ZN(W426));
  NOR2X1 G12260 (.A1(W49528), .A2(W20832), .ZN(O19339));
  NOR2X1 G12261 (.A1(W8825), .A2(W15472), .ZN(W25493));
  NOR2X1 G12262 (.A1(W1239), .A2(W31367), .ZN(O19342));
  NOR2X1 G12263 (.A1(W30312), .A2(W33840), .ZN(O19343));
  NOR2X1 G12264 (.A1(W50123), .A2(W48234), .ZN(O19346));
  NOR2X1 G12265 (.A1(I838), .A2(I839), .ZN(W419));
  NOR2X1 G12266 (.A1(I1470), .A2(W1335), .ZN(W2093));
  NOR2X1 G12267 (.A1(W24438), .A2(W6454), .ZN(W26101));
  NOR2X1 G12268 (.A1(I1462), .A2(W1974), .ZN(W2100));
  NOR2X1 G12269 (.A1(W22165), .A2(W38151), .ZN(O17737));
  NOR2X1 G12270 (.A1(I115), .A2(I527), .ZN(W2098));
  NOR2X1 G12271 (.A1(W45984), .A2(W7582), .ZN(O17738));
  NOR2X1 G12272 (.A1(I109), .A2(W131), .ZN(W2096));
  NOR2X1 G12273 (.A1(W1298), .A2(W587), .ZN(W2095));
  NOR2X1 G12274 (.A1(W35862), .A2(W10855), .ZN(O17740));
  NOR2X1 G12275 (.A1(W1450), .A2(I407), .ZN(W2102));
  NOR2X1 G12276 (.A1(W1633), .A2(W1759), .ZN(W2092));
  NOR2X1 G12277 (.A1(W14512), .A2(W20186), .ZN(O17742));
  NOR2X1 G12278 (.A1(W23790), .A2(W35373), .ZN(O17743));
  NOR2X1 G12279 (.A1(W7136), .A2(W8937), .ZN(W26092));
  NOR2X1 G12280 (.A1(W15753), .A2(W8555), .ZN(W26091));
  NOR2X1 G12281 (.A1(W28172), .A2(W4939), .ZN(O17748));
  NOR2X1 G12282 (.A1(W21411), .A2(W37771), .ZN(O17750));
  NOR2X1 G12283 (.A1(W24456), .A2(I409), .ZN(O17751));
  NOR2X1 G12284 (.A1(W1066), .A2(I1310), .ZN(W2110));
  NOR2X1 G12285 (.A1(W44864), .A2(W18601), .ZN(O17726));
  NOR2X1 G12286 (.A1(I1115), .A2(W1661), .ZN(W2117));
  NOR2X1 G12287 (.A1(W10183), .A2(W14380), .ZN(W26103));
  NOR2X1 G12288 (.A1(W842), .A2(I549), .ZN(W2115));
  NOR2X1 G12289 (.A1(W575), .A2(I6), .ZN(W2114));
  NOR2X1 G12290 (.A1(I744), .A2(W861), .ZN(W2113));
  NOR2X1 G12291 (.A1(W43755), .A2(W42893), .ZN(O17728));
  NOR2X1 G12292 (.A1(I229), .A2(I420), .ZN(O17));
  NOR2X1 G12293 (.A1(I1983), .A2(W904), .ZN(W2082));
  NOR2X1 G12294 (.A1(W5082), .A2(W22790), .ZN(O3632));
  NOR2X1 G12295 (.A1(W33929), .A2(W22597), .ZN(O17731));
  NOR2X1 G12296 (.A1(W25764), .A2(W14752), .ZN(O17733));
  NOR2X1 G12297 (.A1(I1454), .A2(W14), .ZN(W2106));
  NOR2X1 G12298 (.A1(W788), .A2(I804), .ZN(W2105));
  NOR2X1 G12299 (.A1(I24), .A2(I438), .ZN(W2104));
  NOR2X1 G12300 (.A1(W40647), .A2(W26913), .ZN(O17735));
  NOR2X1 G12301 (.A1(W48567), .A2(W26094), .ZN(O17782));
  NOR2X1 G12302 (.A1(W14802), .A2(I817), .ZN(W26083));
  NOR2X1 G12303 (.A1(W37255), .A2(W43431), .ZN(O17771));
  NOR2X1 G12304 (.A1(W45529), .A2(W45761), .ZN(O17775));
  NOR2X1 G12305 (.A1(W592), .A2(W8060), .ZN(O17776));
  NOR2X1 G12306 (.A1(I353), .A2(W1372), .ZN(W2056));
  NOR2X1 G12307 (.A1(W5283), .A2(W17058), .ZN(W24651));
  NOR2X1 G12308 (.A1(W14621), .A2(W18849), .ZN(W24652));
  NOR2X1 G12309 (.A1(W398), .A2(W1884), .ZN(W2051));
  NOR2X1 G12310 (.A1(W7239), .A2(W10150), .ZN(O17768));
  NOR2X1 G12311 (.A1(I952), .A2(I7), .ZN(W2049));
  NOR2X1 G12312 (.A1(W12054), .A2(W2050), .ZN(O17783));
  NOR2X1 G12313 (.A1(W38488), .A2(W27865), .ZN(O17784));
  NOR2X1 G12314 (.A1(W16671), .A2(W40169), .ZN(O17785));
  NOR2X1 G12315 (.A1(W35152), .A2(W6891), .ZN(O17786));
  NOR2X1 G12316 (.A1(W3181), .A2(W47775), .ZN(O17787));
  NOR2X1 G12317 (.A1(I1427), .A2(W286), .ZN(W2043));
  NOR2X1 G12318 (.A1(W2732), .A2(W19346), .ZN(W26080));
  NOR2X1 G12319 (.A1(I222), .A2(I479), .ZN(W2073));
  NOR2X1 G12320 (.A1(I254), .A2(I1570), .ZN(W2081));
  NOR2X1 G12321 (.A1(I162), .A2(W3045), .ZN(O3150));
  NOR2X1 G12322 (.A1(W1373), .A2(W190), .ZN(W2079));
  NOR2X1 G12323 (.A1(W497), .A2(W253), .ZN(W2078));
  NOR2X1 G12324 (.A1(W957), .A2(W15576), .ZN(W24638));
  NOR2X1 G12325 (.A1(I814), .A2(I1952), .ZN(W2076));
  NOR2X1 G12326 (.A1(W11200), .A2(W8201), .ZN(O3627));
  NOR2X1 G12327 (.A1(W10898), .A2(W24333), .ZN(W24640));
  NOR2X1 G12328 (.A1(W5150), .A2(W48396), .ZN(O17724));
  NOR2X1 G12329 (.A1(W43523), .A2(W34766), .ZN(W48913));
  NOR2X1 G12330 (.A1(I1697), .A2(I1590), .ZN(W2067));
  NOR2X1 G12331 (.A1(W1843), .A2(W18379), .ZN(O17762));
  NOR2X1 G12332 (.A1(W9611), .A2(W9775), .ZN(O3624));
  NOR2X1 G12333 (.A1(W34441), .A2(W32734), .ZN(O17764));
  NOR2X1 G12334 (.A1(W20499), .A2(W22349), .ZN(O3153));
  NOR2X1 G12335 (.A1(W23356), .A2(W5832), .ZN(O3154));
  NOR2X1 G12336 (.A1(W372), .A2(W1975), .ZN(W2164));
  NOR2X1 G12337 (.A1(W5215), .A2(W38337), .ZN(O17677));
  NOR2X1 G12338 (.A1(W10875), .A2(W9549), .ZN(O3143));
  NOR2X1 G12339 (.A1(W12096), .A2(W1444), .ZN(O17682));
  NOR2X1 G12340 (.A1(W918), .A2(W1582), .ZN(W2169));
  NOR2X1 G12341 (.A1(I1410), .A2(I137), .ZN(W2168));
  NOR2X1 G12342 (.A1(W7733), .A2(W15310), .ZN(W26111));
  NOR2X1 G12343 (.A1(W11409), .A2(W5259), .ZN(O3635));
  NOR2X1 G12344 (.A1(W48073), .A2(W14688), .ZN(O17686));
  NOR2X1 G12345 (.A1(I1688), .A2(W11180), .ZN(O17675));
  NOR2X1 G12346 (.A1(W13642), .A2(W25708), .ZN(W26109));
  NOR2X1 G12347 (.A1(I533), .A2(W701), .ZN(W2161));
  NOR2X1 G12348 (.A1(W543), .A2(W34549), .ZN(O17693));
  NOR2X1 G12349 (.A1(I164), .A2(W1604), .ZN(W2159));
  NOR2X1 G12350 (.A1(W24088), .A2(W11181), .ZN(O17695));
  NOR2X1 G12351 (.A1(W22866), .A2(W9822), .ZN(O3145));
  NOR2X1 G12352 (.A1(W21021), .A2(W20015), .ZN(O3146));
  NOR2X1 G12353 (.A1(I909), .A2(W718), .ZN(W2155));
  NOR2X1 G12354 (.A1(W40323), .A2(W22396), .ZN(O17664));
  NOR2X1 G12355 (.A1(W1132), .A2(W799), .ZN(W2191));
  NOR2X1 G12356 (.A1(W9597), .A2(W7992), .ZN(W26115));
  NOR2X1 G12357 (.A1(I1509), .A2(I1375), .ZN(W2189));
  NOR2X1 G12358 (.A1(W34018), .A2(W16008), .ZN(O17658));
  NOR2X1 G12359 (.A1(W21420), .A2(W22044), .ZN(O3140));
  NOR2X1 G12360 (.A1(W30012), .A2(W11077), .ZN(O17663));
  NOR2X1 G12361 (.A1(I1679), .A2(I1586), .ZN(W2185));
  NOR2X1 G12362 (.A1(W1009), .A2(I909), .ZN(W2184));
  NOR2X1 G12363 (.A1(I871), .A2(I874), .ZN(W2154));
  NOR2X1 G12364 (.A1(W27841), .A2(W30633), .ZN(O17668));
  NOR2X1 G12365 (.A1(W17718), .A2(W12308), .ZN(W24615));
  NOR2X1 G12366 (.A1(W532), .A2(W1412), .ZN(W2179));
  NOR2X1 G12367 (.A1(W306), .A2(I1695), .ZN(W2177));
  NOR2X1 G12368 (.A1(W2683), .A2(W1542), .ZN(O3142));
  NOR2X1 G12369 (.A1(W32479), .A2(W38272), .ZN(O17674));
  NOR2X1 G12370 (.A1(W812), .A2(I903), .ZN(W2174));
  NOR2X1 G12371 (.A1(W82), .A2(W24363), .ZN(O17720));
  NOR2X1 G12372 (.A1(I986), .A2(W2098), .ZN(O17711));
  NOR2X1 G12373 (.A1(W36149), .A2(W28641), .ZN(O17712));
  NOR2X1 G12374 (.A1(W23389), .A2(W12142), .ZN(O17713));
  NOR2X1 G12375 (.A1(W23127), .A2(W6593), .ZN(W24627));
  NOR2X1 G12376 (.A1(I1570), .A2(W216), .ZN(W2132));
  NOR2X1 G12377 (.A1(W31361), .A2(W36532), .ZN(O17716));
  NOR2X1 G12378 (.A1(W32510), .A2(W16862), .ZN(O17718));
  NOR2X1 G12379 (.A1(W3956), .A2(W17500), .ZN(W26106));
  NOR2X1 G12380 (.A1(W21373), .A2(W23450), .ZN(O17710));
  NOR2X1 G12381 (.A1(I1395), .A2(I1533), .ZN(W2127));
  NOR2X1 G12382 (.A1(W2062), .A2(I1565), .ZN(W2126));
  NOR2X1 G12383 (.A1(W21554), .A2(W40516), .ZN(W48877));
  NOR2X1 G12384 (.A1(W11558), .A2(W5154), .ZN(O17723));
  NOR2X1 G12385 (.A1(W1332), .A2(W924), .ZN(W2123));
  NOR2X1 G12386 (.A1(W1608), .A2(W206), .ZN(W2122));
  NOR2X1 G12387 (.A1(W1599), .A2(I1720), .ZN(W2121));
  NOR2X1 G12388 (.A1(I412), .A2(W1285), .ZN(W2145));
  NOR2X1 G12389 (.A1(W15406), .A2(W2065), .ZN(W24625));
  NOR2X1 G12390 (.A1(W20235), .A2(W43200), .ZN(O17699));
  NOR2X1 G12391 (.A1(I336), .A2(W1247), .ZN(W2151));
  NOR2X1 G12392 (.A1(W4695), .A2(W23012), .ZN(O17700));
  NOR2X1 G12393 (.A1(W30), .A2(W1837), .ZN(W2149));
  NOR2X1 G12394 (.A1(W13443), .A2(W21171), .ZN(O17701));
  NOR2X1 G12395 (.A1(W48848), .A2(W24566), .ZN(O17703));
  NOR2X1 G12396 (.A1(W11556), .A2(W33215), .ZN(O17704));
  NOR2X1 G12397 (.A1(W1174), .A2(W486), .ZN(W2041));
  NOR2X1 G12398 (.A1(W695), .A2(I1245), .ZN(W2144));
  NOR2X1 G12399 (.A1(W42797), .A2(W7996), .ZN(O17705));
  NOR2X1 G12400 (.A1(W17513), .A2(W18518), .ZN(O3634));
  NOR2X1 G12401 (.A1(W1852), .A2(W1285), .ZN(W2141));
  NOR2X1 G12402 (.A1(W10577), .A2(W14781), .ZN(O17709));
  NOR2X1 G12403 (.A1(I385), .A2(I1591), .ZN(W2139));
  NOR2X1 G12404 (.A1(W1640), .A2(W1182), .ZN(W2138));
  NOR2X1 G12405 (.A1(I1800), .A2(W1506), .ZN(W1932));
  NOR2X1 G12406 (.A1(I1378), .A2(I632), .ZN(W1943));
  NOR2X1 G12407 (.A1(W31842), .A2(W28542), .ZN(W49055));
  NOR2X1 G12408 (.A1(W17776), .A2(W9772), .ZN(W26042));
  NOR2X1 G12409 (.A1(I1306), .A2(W4762), .ZN(O3607));
  NOR2X1 G12410 (.A1(W16866), .A2(W36758), .ZN(O17890));
  NOR2X1 G12411 (.A1(I1646), .A2(W35732), .ZN(O17891));
  NOR2X1 G12412 (.A1(W14085), .A2(W11138), .ZN(O17893));
  NOR2X1 G12413 (.A1(W7687), .A2(W36509), .ZN(O17894));
  NOR2X1 G12414 (.A1(W637), .A2(W474), .ZN(W1944));
  NOR2X1 G12415 (.A1(W40999), .A2(W18887), .ZN(O17895));
  NOR2X1 G12416 (.A1(W1541), .A2(W255), .ZN(W1930));
  NOR2X1 G12417 (.A1(W10509), .A2(W31764), .ZN(O17897));
  NOR2X1 G12418 (.A1(W17520), .A2(W12388), .ZN(W24690));
  NOR2X1 G12419 (.A1(W8955), .A2(I55), .ZN(W24692));
  NOR2X1 G12420 (.A1(I1976), .A2(W1866), .ZN(W1924));
  NOR2X1 G12421 (.A1(I1211), .A2(W1866), .ZN(W1923));
  NOR2X1 G12422 (.A1(W45209), .A2(W5934), .ZN(O17903));
  NOR2X1 G12423 (.A1(W15251), .A2(W3680), .ZN(O17873));
  NOR2X1 G12424 (.A1(W6339), .A2(W38818), .ZN(O17863));
  NOR2X1 G12425 (.A1(I720), .A2(W25423), .ZN(W26055));
  NOR2X1 G12426 (.A1(I283), .A2(I904), .ZN(W1961));
  NOR2X1 G12427 (.A1(I925), .A2(W545), .ZN(W1960));
  NOR2X1 G12428 (.A1(W29308), .A2(W27168), .ZN(O17868));
  NOR2X1 G12429 (.A1(I412), .A2(W1630), .ZN(W1958));
  NOR2X1 G12430 (.A1(I364), .A2(W232), .ZN(W1957));
  NOR2X1 G12431 (.A1(W983), .A2(W22300), .ZN(O17872));
  NOR2X1 G12432 (.A1(W37890), .A2(W44497), .ZN(O17904));
  NOR2X1 G12433 (.A1(I1029), .A2(I1572), .ZN(W1953));
  NOR2X1 G12434 (.A1(W1721), .A2(W891), .ZN(W1951));
  NOR2X1 G12435 (.A1(I26), .A2(W16652), .ZN(W24681));
  NOR2X1 G12436 (.A1(W47547), .A2(W5884), .ZN(O17877));
  NOR2X1 G12437 (.A1(W14063), .A2(W21149), .ZN(W26044));
  NOR2X1 G12438 (.A1(W11947), .A2(W29011), .ZN(O17884));
  NOR2X1 G12439 (.A1(W208), .A2(I491), .ZN(W1945));
  NOR2X1 G12440 (.A1(W1287), .A2(W1168), .ZN(W1889));
  NOR2X1 G12441 (.A1(W24778), .A2(W29543), .ZN(O17921));
  NOR2X1 G12442 (.A1(W1519), .A2(W1258), .ZN(W1897));
  NOR2X1 G12443 (.A1(W10091), .A2(W4208), .ZN(W26020));
  NOR2X1 G12444 (.A1(I1263), .A2(W359), .ZN(W1895));
  NOR2X1 G12445 (.A1(W45720), .A2(W36216), .ZN(O17923));
  NOR2X1 G12446 (.A1(W39013), .A2(W40537), .ZN(O17925));
  NOR2X1 G12447 (.A1(W33127), .A2(W36663), .ZN(O17927));
  NOR2X1 G12448 (.A1(W10624), .A2(W22355), .ZN(W24707));
  NOR2X1 G12449 (.A1(W375), .A2(I1935), .ZN(W1899));
  NOR2X1 G12450 (.A1(I339), .A2(I1441), .ZN(W1888));
  NOR2X1 G12451 (.A1(W11205), .A2(W37990), .ZN(O17930));
  NOR2X1 G12452 (.A1(I1110), .A2(W20663), .ZN(W24709));
  NOR2X1 G12453 (.A1(W32830), .A2(W43635), .ZN(O17934));
  NOR2X1 G12454 (.A1(W21114), .A2(W25764), .ZN(W26014));
  NOR2X1 G12455 (.A1(W10412), .A2(W38992), .ZN(O17938));
  NOR2X1 G12456 (.A1(W1122), .A2(I1392), .ZN(W1880));
  NOR2X1 G12457 (.A1(W20905), .A2(W10695), .ZN(W26027));
  NOR2X1 G12458 (.A1(W13587), .A2(W21666), .ZN(W24693));
  NOR2X1 G12459 (.A1(W1049), .A2(I916), .ZN(W1919));
  NOR2X1 G12460 (.A1(W1431), .A2(W1340), .ZN(W1918));
  NOR2X1 G12461 (.A1(I79), .A2(W520), .ZN(W1916));
  NOR2X1 G12462 (.A1(W639), .A2(W760), .ZN(W1914));
  NOR2X1 G12463 (.A1(W827), .A2(W1793), .ZN(W1913));
  NOR2X1 G12464 (.A1(I1193), .A2(W17580), .ZN(O3605));
  NOR2X1 G12465 (.A1(W23394), .A2(W21207), .ZN(W24697));
  NOR2X1 G12466 (.A1(W11573), .A2(W28354), .ZN(W49029));
  NOR2X1 G12467 (.A1(W12381), .A2(W17966), .ZN(O3168));
  NOR2X1 G12468 (.A1(W5070), .A2(W13953), .ZN(W24701));
  NOR2X1 G12469 (.A1(W167), .A2(W1727), .ZN(W1906));
  NOR2X1 G12470 (.A1(W21796), .A2(W12216), .ZN(O17915));
  NOR2X1 G12471 (.A1(W1003), .A2(I271), .ZN(W1903));
  NOR2X1 G12472 (.A1(W3845), .A2(W6473), .ZN(W26023));
  NOR2X1 G12473 (.A1(W205), .A2(I574), .ZN(W1900));
  NOR2X1 G12474 (.A1(W30089), .A2(W8423), .ZN(O17814));
  NOR2X1 G12475 (.A1(W47381), .A2(W24532), .ZN(O17805));
  NOR2X1 G12476 (.A1(W19819), .A2(W8129), .ZN(O3157));
  NOR2X1 G12477 (.A1(W48557), .A2(W30465), .ZN(W48969));
  NOR2X1 G12478 (.A1(W19030), .A2(W44088), .ZN(O17807));
  NOR2X1 G12479 (.A1(W1465), .A2(I1578), .ZN(W2016));
  NOR2X1 G12480 (.A1(W38094), .A2(W28832), .ZN(O17811));
  NOR2X1 G12481 (.A1(W41981), .A2(W9714), .ZN(W48976));
  NOR2X1 G12482 (.A1(W1466), .A2(I444), .ZN(W2011));
  NOR2X1 G12483 (.A1(W22147), .A2(W2033), .ZN(O3619));
  NOR2X1 G12484 (.A1(W1963), .A2(I1928), .ZN(W2008));
  NOR2X1 G12485 (.A1(W937), .A2(W17088), .ZN(W24665));
  NOR2X1 G12486 (.A1(W674), .A2(W763), .ZN(W2006));
  NOR2X1 G12487 (.A1(W21070), .A2(W346), .ZN(W24666));
  NOR2X1 G12488 (.A1(W22190), .A2(W25776), .ZN(W26069));
  NOR2X1 G12489 (.A1(W742), .A2(I1552), .ZN(W2003));
  NOR2X1 G12490 (.A1(W492), .A2(W75), .ZN(W2002));
  NOR2X1 G12491 (.A1(W1526), .A2(W1063), .ZN(W2001));
  NOR2X1 G12492 (.A1(W1163), .A2(W401), .ZN(W2031));
  NOR2X1 G12493 (.A1(W672), .A2(I1303), .ZN(W2040));
  NOR2X1 G12494 (.A1(W38738), .A2(W35421), .ZN(O17790));
  NOR2X1 G12495 (.A1(W1651), .A2(W2002), .ZN(W2037));
  NOR2X1 G12496 (.A1(I140), .A2(I1358), .ZN(W2036));
  NOR2X1 G12497 (.A1(W176), .A2(I71), .ZN(W2035));
  NOR2X1 G12498 (.A1(W42104), .A2(W7382), .ZN(O17792));
  NOR2X1 G12499 (.A1(W4282), .A2(W22087), .ZN(O17793));
  NOR2X1 G12500 (.A1(W37752), .A2(W31067), .ZN(O17794));
  NOR2X1 G12501 (.A1(I1068), .A2(W1522), .ZN(W2000));
  NOR2X1 G12502 (.A1(W3395), .A2(W43726), .ZN(O17795));
  NOR2X1 G12503 (.A1(W19885), .A2(W2169), .ZN(O17799));
  NOR2X1 G12504 (.A1(I1561), .A2(I1490), .ZN(W2026));
  NOR2X1 G12505 (.A1(W420), .A2(W1790), .ZN(W2025));
  NOR2X1 G12506 (.A1(W21499), .A2(W21647), .ZN(O3621));
  NOR2X1 G12507 (.A1(W23087), .A2(W13154), .ZN(O3155));
  NOR2X1 G12508 (.A1(W17085), .A2(W20322), .ZN(O3156));
  NOR2X1 G12509 (.A1(I1321), .A2(I1148), .ZN(W1973));
  NOR2X1 G12510 (.A1(I1247), .A2(W1590), .ZN(W1982));
  NOR2X1 G12511 (.A1(I1345), .A2(I86), .ZN(W1981));
  NOR2X1 G12512 (.A1(W44075), .A2(W44153), .ZN(O17850));
  NOR2X1 G12513 (.A1(W17), .A2(I1542), .ZN(W1979));
  NOR2X1 G12514 (.A1(W14832), .A2(W9849), .ZN(W26063));
  NOR2X1 G12515 (.A1(I1220), .A2(W1281), .ZN(W1976));
  NOR2X1 G12516 (.A1(W42065), .A2(W6224), .ZN(O17855));
  NOR2X1 G12517 (.A1(I1493), .A2(W1170), .ZN(W1974));
  NOR2X1 G12518 (.A1(W12865), .A2(W200), .ZN(W26064));
  NOR2X1 G12519 (.A1(I163), .A2(I358), .ZN(W1972));
  NOR2X1 G12520 (.A1(W161), .A2(I1975), .ZN(W1971));
  NOR2X1 G12521 (.A1(W12011), .A2(W9354), .ZN(O3160));
  NOR2X1 G12522 (.A1(W1680), .A2(W36931), .ZN(O17859));
  NOR2X1 G12523 (.A1(I1552), .A2(W42585), .ZN(O17860));
  NOR2X1 G12524 (.A1(W1062), .A2(W799), .ZN(W1967));
  NOR2X1 G12525 (.A1(W634), .A2(W2980), .ZN(W26060));
  NOR2X1 G12526 (.A1(W5760), .A2(I330), .ZN(O17837));
  NOR2X1 G12527 (.A1(I31), .A2(W46025), .ZN(O17822));
  NOR2X1 G12528 (.A1(W2576), .A2(W44699), .ZN(O17823));
  NOR2X1 G12529 (.A1(W42274), .A2(W47162), .ZN(O17825));
  NOR2X1 G12530 (.A1(W40025), .A2(W17365), .ZN(O17826));
  NOR2X1 G12531 (.A1(W14388), .A2(W6590), .ZN(W26068));
  NOR2X1 G12532 (.A1(W9882), .A2(W25403), .ZN(O17832));
  NOR2X1 G12533 (.A1(W11455), .A2(W24587), .ZN(O17834));
  NOR2X1 G12534 (.A1(W12702), .A2(W12454), .ZN(W24669));
  NOR2X1 G12535 (.A1(W12738), .A2(I1513), .ZN(W24611));
  NOR2X1 G12536 (.A1(W16436), .A2(W18980), .ZN(W26067));
  NOR2X1 G12537 (.A1(I1195), .A2(W4114), .ZN(O17840));
  NOR2X1 G12538 (.A1(W586), .A2(I36), .ZN(W1988));
  NOR2X1 G12539 (.A1(W29751), .A2(W13290), .ZN(O17841));
  NOR2X1 G12540 (.A1(W1239), .A2(W262), .ZN(W1986));
  NOR2X1 G12541 (.A1(W7536), .A2(W22320), .ZN(W26065));
  NOR2X1 G12542 (.A1(W30691), .A2(W46615), .ZN(W49007));
  NOR2X1 G12543 (.A1(W17733), .A2(W46475), .ZN(O17450));
  NOR2X1 G12544 (.A1(I305), .A2(W698), .ZN(W2408));
  NOR2X1 G12545 (.A1(W38751), .A2(W16668), .ZN(O17441));
  NOR2X1 G12546 (.A1(I831), .A2(W1865), .ZN(W2406));
  NOR2X1 G12547 (.A1(W17973), .A2(W16749), .ZN(O17442));
  NOR2X1 G12548 (.A1(W1800), .A2(W714), .ZN(W2404));
  NOR2X1 G12549 (.A1(W37000), .A2(W43618), .ZN(O17443));
  NOR2X1 G12550 (.A1(W8216), .A2(W20060), .ZN(O17445));
  NOR2X1 G12551 (.A1(I1040), .A2(W1454), .ZN(O3110));
  NOR2X1 G12552 (.A1(W22743), .A2(W26616), .ZN(W48567));
  NOR2X1 G12553 (.A1(I1803), .A2(W24104), .ZN(O3111));
  NOR2X1 G12554 (.A1(I74), .A2(W1465), .ZN(W2397));
  NOR2X1 G12555 (.A1(W39877), .A2(W43587), .ZN(O17452));
  NOR2X1 G12556 (.A1(W1677), .A2(W1208), .ZN(W2395));
  NOR2X1 G12557 (.A1(W2041), .A2(I1571), .ZN(W2394));
  NOR2X1 G12558 (.A1(W4000), .A2(W28825), .ZN(O17456));
  NOR2X1 G12559 (.A1(W36222), .A2(W33578), .ZN(O17459));
  NOR2X1 G12560 (.A1(W266), .A2(I1944), .ZN(W2390));
  NOR2X1 G12561 (.A1(I868), .A2(W26), .ZN(W2417));
  NOR2X1 G12562 (.A1(W185), .A2(W1590), .ZN(W2426));
  NOR2X1 G12563 (.A1(W888), .A2(W1815), .ZN(W2425));
  NOR2X1 G12564 (.A1(W23307), .A2(I622), .ZN(W48553));
  NOR2X1 G12565 (.A1(W832), .A2(W1768), .ZN(W2423));
  NOR2X1 G12566 (.A1(W47815), .A2(W46895), .ZN(O17433));
  NOR2X1 G12567 (.A1(I622), .A2(W29220), .ZN(W48557));
  NOR2X1 G12568 (.A1(I1523), .A2(W18963), .ZN(W24538));
  NOR2X1 G12569 (.A1(I1298), .A2(W5309), .ZN(W24539));
  NOR2X1 G12570 (.A1(W22279), .A2(W12708), .ZN(O17464));
  NOR2X1 G12571 (.A1(I714), .A2(W958), .ZN(W2416));
  NOR2X1 G12572 (.A1(W74), .A2(W1778), .ZN(W2415));
  NOR2X1 G12573 (.A1(W13987), .A2(W32370), .ZN(W48563));
  NOR2X1 G12574 (.A1(W2296), .A2(W2219), .ZN(W2413));
  NOR2X1 G12575 (.A1(I1252), .A2(W14116), .ZN(O3670));
  NOR2X1 G12576 (.A1(W24071), .A2(W29023), .ZN(O17440));
  NOR2X1 G12577 (.A1(W1400), .A2(W6), .ZN(W2410));
  NOR2X1 G12578 (.A1(W24731), .A2(W24036), .ZN(O3663));
  NOR2X1 G12579 (.A1(W20301), .A2(W44682), .ZN(O17484));
  NOR2X1 G12580 (.A1(W42187), .A2(W9092), .ZN(O17485));
  NOR2X1 G12581 (.A1(W9200), .A2(W29161), .ZN(O17487));
  NOR2X1 G12582 (.A1(W33425), .A2(W17077), .ZN(O17488));
  NOR2X1 G12583 (.A1(W9112), .A2(W13798), .ZN(W26173));
  NOR2X1 G12584 (.A1(W3319), .A2(W14039), .ZN(O17493));
  NOR2X1 G12585 (.A1(W13485), .A2(W13527), .ZN(O17494));
  NOR2X1 G12586 (.A1(W23312), .A2(W2168), .ZN(O17495));
  NOR2X1 G12587 (.A1(W122), .A2(W729), .ZN(W2370));
  NOR2X1 G12588 (.A1(W1523), .A2(I916), .ZN(W2359));
  NOR2X1 G12589 (.A1(W19456), .A2(W21951), .ZN(W24555));
  NOR2X1 G12590 (.A1(W134), .A2(W1474), .ZN(W2357));
  NOR2X1 G12591 (.A1(W11312), .A2(W18385), .ZN(O3115));
  NOR2X1 G12592 (.A1(I324), .A2(W9495), .ZN(W24557));
  NOR2X1 G12593 (.A1(W29855), .A2(W28611), .ZN(O17504));
  NOR2X1 G12594 (.A1(W1), .A2(W9768), .ZN(O3662));
  NOR2X1 G12595 (.A1(W107), .A2(W2220), .ZN(W2379));
  NOR2X1 G12596 (.A1(W2348), .A2(W291), .ZN(W2388));
  NOR2X1 G12597 (.A1(W5844), .A2(W7421), .ZN(O3112));
  NOR2X1 G12598 (.A1(W13333), .A2(W4028), .ZN(O17467));
  NOR2X1 G12599 (.A1(W14596), .A2(W10022), .ZN(O3666));
  NOR2X1 G12600 (.A1(W22706), .A2(W45918), .ZN(W48602));
  NOR2X1 G12601 (.A1(W43798), .A2(W36956), .ZN(O17474));
  NOR2X1 G12602 (.A1(W16923), .A2(W19255), .ZN(O3114));
  NOR2X1 G12603 (.A1(W17037), .A2(W19873), .ZN(W26177));
  NOR2X1 G12604 (.A1(W44762), .A2(W40238), .ZN(O17430));
  NOR2X1 G12605 (.A1(I1332), .A2(W2327), .ZN(W2377));
  NOR2X1 G12606 (.A1(W21631), .A2(W23407), .ZN(W24551));
  NOR2X1 G12607 (.A1(W24077), .A2(W21022), .ZN(W48614));
  NOR2X1 G12608 (.A1(W11070), .A2(W20521), .ZN(O17483));
  NOR2X1 G12609 (.A1(W1455), .A2(W2036), .ZN(W2373));
  NOR2X1 G12610 (.A1(I1332), .A2(I994), .ZN(W2372));
  NOR2X1 G12611 (.A1(I827), .A2(W26), .ZN(W2371));
  NOR2X1 G12612 (.A1(W8063), .A2(W23479), .ZN(W24516));
  NOR2X1 G12613 (.A1(W27435), .A2(W25599), .ZN(O17370));
  NOR2X1 G12614 (.A1(W16341), .A2(W30277), .ZN(O17372));
  NOR2X1 G12615 (.A1(W1189), .A2(I794), .ZN(W2489));
  NOR2X1 G12616 (.A1(I1254), .A2(W1493), .ZN(W2488));
  NOR2X1 G12617 (.A1(I1144), .A2(I390), .ZN(W2487));
  NOR2X1 G12618 (.A1(I527), .A2(I23), .ZN(W2486));
  NOR2X1 G12619 (.A1(W4861), .A2(W22637), .ZN(O17373));
  NOR2X1 G12620 (.A1(W769), .A2(I1802), .ZN(O3680));
  NOR2X1 G12621 (.A1(W13124), .A2(W2029), .ZN(O17368));
  NOR2X1 G12622 (.A1(W18820), .A2(W20825), .ZN(W26213));
  NOR2X1 G12623 (.A1(W1656), .A2(W18737), .ZN(O17378));
  NOR2X1 G12624 (.A1(W22400), .A2(W19064), .ZN(W24518));
  NOR2X1 G12625 (.A1(W423), .A2(W10308), .ZN(W24519));
  NOR2X1 G12626 (.A1(I1188), .A2(I1501), .ZN(W2478));
  NOR2X1 G12627 (.A1(W20186), .A2(W5745), .ZN(W24520));
  NOR2X1 G12628 (.A1(W1523), .A2(W1443), .ZN(W2475));
  NOR2X1 G12629 (.A1(W295), .A2(W193), .ZN(O3676));
  NOR2X1 G12630 (.A1(W510), .A2(W844), .ZN(W2503));
  NOR2X1 G12631 (.A1(W2384), .A2(W2239), .ZN(W2514));
  NOR2X1 G12632 (.A1(W30195), .A2(W47007), .ZN(O17351));
  NOR2X1 G12633 (.A1(W45543), .A2(W3460), .ZN(O17353));
  NOR2X1 G12634 (.A1(W28015), .A2(W34018), .ZN(O17355));
  NOR2X1 G12635 (.A1(W44326), .A2(W46219), .ZN(W48469));
  NOR2X1 G12636 (.A1(W1146), .A2(W489), .ZN(W2506));
  NOR2X1 G12637 (.A1(W26401), .A2(W39887), .ZN(O17357));
  NOR2X1 G12638 (.A1(W17360), .A2(W17056), .ZN(O3684));
  NOR2X1 G12639 (.A1(W1037), .A2(I518), .ZN(W2471));
  NOR2X1 G12640 (.A1(W48136), .A2(W35300), .ZN(O17361));
  NOR2X1 G12641 (.A1(W27631), .A2(W41778), .ZN(O17362));
  NOR2X1 G12642 (.A1(W25571), .A2(W21339), .ZN(O17365));
  NOR2X1 G12643 (.A1(W37773), .A2(W18487), .ZN(O17366));
  NOR2X1 G12644 (.A1(I840), .A2(I1714), .ZN(W2497));
  NOR2X1 G12645 (.A1(W38599), .A2(W17595), .ZN(O17367));
  NOR2X1 G12646 (.A1(I1330), .A2(W295), .ZN(W2495));
  NOR2X1 G12647 (.A1(I1982), .A2(I1390), .ZN(W2436));
  NOR2X1 G12648 (.A1(I1266), .A2(I724), .ZN(W2445));
  NOR2X1 G12649 (.A1(W13046), .A2(W15514), .ZN(O17420));
  NOR2X1 G12650 (.A1(W2168), .A2(W1767), .ZN(W2443));
  NOR2X1 G12651 (.A1(I418), .A2(W1258), .ZN(W2442));
  NOR2X1 G12652 (.A1(W2585), .A2(W5737), .ZN(O17421));
  NOR2X1 G12653 (.A1(W1981), .A2(W737), .ZN(W2439));
  NOR2X1 G12654 (.A1(W19130), .A2(W21751), .ZN(O17422));
  NOR2X1 G12655 (.A1(W664), .A2(I1026), .ZN(W2437));
  NOR2X1 G12656 (.A1(W20845), .A2(W25153), .ZN(O17415));
  NOR2X1 G12657 (.A1(W2153), .A2(W1468), .ZN(W2435));
  NOR2X1 G12658 (.A1(W651), .A2(I1245), .ZN(W2434));
  NOR2X1 G12659 (.A1(I1339), .A2(W5609), .ZN(W26193));
  NOR2X1 G12660 (.A1(W29500), .A2(W37006), .ZN(O17423));
  NOR2X1 G12661 (.A1(W4842), .A2(W7940), .ZN(W26192));
  NOR2X1 G12662 (.A1(I1119), .A2(W36804), .ZN(O17425));
  NOR2X1 G12663 (.A1(W21020), .A2(W38722), .ZN(O17428));
  NOR2X1 G12664 (.A1(W165), .A2(W119), .ZN(W2459));
  NOR2X1 G12665 (.A1(W2332), .A2(W1310), .ZN(W2470));
  NOR2X1 G12666 (.A1(W17230), .A2(W3572), .ZN(O17389));
  NOR2X1 G12667 (.A1(I544), .A2(W107), .ZN(O17390));
  NOR2X1 G12668 (.A1(W34466), .A2(W48325), .ZN(O17392));
  NOR2X1 G12669 (.A1(W44415), .A2(W22984), .ZN(O17393));
  NOR2X1 G12670 (.A1(W15918), .A2(W31710), .ZN(O17394));
  NOR2X1 G12671 (.A1(W36071), .A2(W34905), .ZN(O17398));
  NOR2X1 G12672 (.A1(I695), .A2(I1692), .ZN(W2461));
  NOR2X1 G12673 (.A1(W574), .A2(W1428), .ZN(W2352));
  NOR2X1 G12674 (.A1(W40771), .A2(W37425), .ZN(O17400));
  NOR2X1 G12675 (.A1(W1151), .A2(I56), .ZN(W2457));
  NOR2X1 G12676 (.A1(W3377), .A2(I908), .ZN(O17401));
  NOR2X1 G12677 (.A1(W4033), .A2(W35011), .ZN(O17402));
  NOR2X1 G12678 (.A1(W27256), .A2(W10732), .ZN(O17409));
  NOR2X1 G12679 (.A1(W45449), .A2(W35714), .ZN(O17413));
  NOR2X1 G12680 (.A1(W375), .A2(W519), .ZN(W2448));
  NOR2X1 G12681 (.A1(W21445), .A2(W9409), .ZN(W24599));
  NOR2X1 G12682 (.A1(I811), .A2(I1381), .ZN(W2248));
  NOR2X1 G12683 (.A1(W3865), .A2(W23493), .ZN(O17606));
  NOR2X1 G12684 (.A1(I13), .A2(W1275), .ZN(W2246));
  NOR2X1 G12685 (.A1(W16064), .A2(W3980), .ZN(W24597));
  NOR2X1 G12686 (.A1(W25801), .A2(W13544), .ZN(O3644));
  NOR2X1 G12687 (.A1(I4), .A2(I500), .ZN(W2242));
  NOR2X1 G12688 (.A1(W10700), .A2(W35844), .ZN(O17611));
  NOR2X1 G12689 (.A1(I797), .A2(W1391), .ZN(W2240));
  NOR2X1 G12690 (.A1(I636), .A2(I560), .ZN(W2249));
  NOR2X1 G12691 (.A1(W4880), .A2(W17727), .ZN(O17614));
  NOR2X1 G12692 (.A1(W17850), .A2(W17014), .ZN(O3133));
  NOR2X1 G12693 (.A1(I1042), .A2(W548), .ZN(W2236));
  NOR2X1 G12694 (.A1(W1895), .A2(W1534), .ZN(W2235));
  NOR2X1 G12695 (.A1(W2134), .A2(W2219), .ZN(W2234));
  NOR2X1 G12696 (.A1(W29549), .A2(W26397), .ZN(O17616));
  NOR2X1 G12697 (.A1(I1928), .A2(I1959), .ZN(W2232));
  NOR2X1 G12698 (.A1(W707), .A2(W673), .ZN(W2231));
  NOR2X1 G12699 (.A1(W9030), .A2(W41485), .ZN(O17596));
  NOR2X1 G12700 (.A1(I246), .A2(W2125), .ZN(W2269));
  NOR2X1 G12701 (.A1(W6169), .A2(W39038), .ZN(O17585));
  NOR2X1 G12702 (.A1(W11783), .A2(I1834), .ZN(O17589));
  NOR2X1 G12703 (.A1(W352), .A2(W4573), .ZN(W24592));
  NOR2X1 G12704 (.A1(W6478), .A2(I526), .ZN(O17593));
  NOR2X1 G12705 (.A1(W14501), .A2(W45141), .ZN(O17595));
  NOR2X1 G12706 (.A1(I928), .A2(I1149), .ZN(W2261));
  NOR2X1 G12707 (.A1(W13962), .A2(W6490), .ZN(W26135));
  NOR2X1 G12708 (.A1(W12013), .A2(W35255), .ZN(O17617));
  NOR2X1 G12709 (.A1(W35236), .A2(W15576), .ZN(O17598));
  NOR2X1 G12710 (.A1(W2043), .A2(I1440), .ZN(W2257));
  NOR2X1 G12711 (.A1(W47853), .A2(W44163), .ZN(O17600));
  NOR2X1 G12712 (.A1(W31564), .A2(W42369), .ZN(O17602));
  NOR2X1 G12713 (.A1(W29580), .A2(W44588), .ZN(O17604));
  NOR2X1 G12714 (.A1(I451), .A2(W820), .ZN(O18));
  NOR2X1 G12715 (.A1(W951), .A2(W1999), .ZN(W2250));
  NOR2X1 G12716 (.A1(W23796), .A2(W13556), .ZN(O17643));
  NOR2X1 G12717 (.A1(W24671), .A2(W27819), .ZN(O17632));
  NOR2X1 G12718 (.A1(W29129), .A2(W3456), .ZN(O17633));
  NOR2X1 G12719 (.A1(W13630), .A2(W14663), .ZN(O3137));
  NOR2X1 G12720 (.A1(W11892), .A2(W43186), .ZN(O17637));
  NOR2X1 G12721 (.A1(W44029), .A2(W38024), .ZN(O17639));
  NOR2X1 G12722 (.A1(W1339), .A2(W30), .ZN(W2204));
  NOR2X1 G12723 (.A1(W14522), .A2(W31764), .ZN(O17640));
  NOR2X1 G12724 (.A1(W14760), .A2(W42573), .ZN(W48788));
  NOR2X1 G12725 (.A1(W645), .A2(W1130), .ZN(W2213));
  NOR2X1 G12726 (.A1(W44824), .A2(W32667), .ZN(O17645));
  NOR2X1 G12727 (.A1(W29396), .A2(W45470), .ZN(O17648));
  NOR2X1 G12728 (.A1(W25490), .A2(W47008), .ZN(O17649));
  NOR2X1 G12729 (.A1(W1432), .A2(W24888), .ZN(O17650));
  NOR2X1 G12730 (.A1(W20801), .A2(W17314), .ZN(W24610));
  NOR2X1 G12731 (.A1(W32658), .A2(W43094), .ZN(O17653));
  NOR2X1 G12732 (.A1(W30860), .A2(W39323), .ZN(O17654));
  NOR2X1 G12733 (.A1(W1161), .A2(I1548), .ZN(W2221));
  NOR2X1 G12734 (.A1(W8460), .A2(W1415), .ZN(O3643));
  NOR2X1 G12735 (.A1(W21991), .A2(W48322), .ZN(O17623));
  NOR2X1 G12736 (.A1(W3190), .A2(W11905), .ZN(O3642));
  NOR2X1 G12737 (.A1(I1795), .A2(I1317), .ZN(W2226));
  NOR2X1 G12738 (.A1(W1059), .A2(I1079), .ZN(W2225));
  NOR2X1 G12739 (.A1(W2356), .A2(W34367), .ZN(O17627));
  NOR2X1 G12740 (.A1(W178), .A2(W1975), .ZN(W2223));
  NOR2X1 G12741 (.A1(I1931), .A2(W1341), .ZN(W2222));
  NOR2X1 G12742 (.A1(W1546), .A2(W5613), .ZN(O3130));
  NOR2X1 G12743 (.A1(W33488), .A2(W17906), .ZN(O17629));
  NOR2X1 G12744 (.A1(W19387), .A2(W24216), .ZN(W24603));
  NOR2X1 G12745 (.A1(W5563), .A2(I227), .ZN(W48775));
  NOR2X1 G12746 (.A1(W41142), .A2(W42385), .ZN(O17631));
  NOR2X1 G12747 (.A1(W8983), .A2(W20730), .ZN(W26124));
  NOR2X1 G12748 (.A1(W754), .A2(W1905), .ZN(W2215));
  NOR2X1 G12749 (.A1(W120), .A2(W800), .ZN(W2214));
  NOR2X1 G12750 (.A1(W33702), .A2(W42385), .ZN(O17540));
  NOR2X1 G12751 (.A1(W23620), .A2(W30339), .ZN(O17530));
  NOR2X1 G12752 (.A1(W36736), .A2(W45171), .ZN(O17533));
  NOR2X1 G12753 (.A1(W7250), .A2(W19036), .ZN(W26160));
  NOR2X1 G12754 (.A1(W33728), .A2(W12629), .ZN(W48670));
  NOR2X1 G12755 (.A1(I1760), .A2(W316), .ZN(W2325));
  NOR2X1 G12756 (.A1(W24862), .A2(W2354), .ZN(W26158));
  NOR2X1 G12757 (.A1(I534), .A2(W16235), .ZN(O3656));
  NOR2X1 G12758 (.A1(W30672), .A2(W46489), .ZN(O17538));
  NOR2X1 G12759 (.A1(W35939), .A2(W1044), .ZN(O17529));
  NOR2X1 G12760 (.A1(W14212), .A2(W14482), .ZN(O3655));
  NOR2X1 G12761 (.A1(W7339), .A2(W7280), .ZN(W26152));
  NOR2X1 G12762 (.A1(W2202), .A2(W379), .ZN(W2316));
  NOR2X1 G12763 (.A1(I755), .A2(I968), .ZN(W2315));
  NOR2X1 G12764 (.A1(W26610), .A2(W25139), .ZN(O17547));
  NOR2X1 G12765 (.A1(W6203), .A2(I1777), .ZN(O3654));
  NOR2X1 G12766 (.A1(W1023), .A2(W1958), .ZN(W2312));
  NOR2X1 G12767 (.A1(W8351), .A2(W15903), .ZN(W24574));
  NOR2X1 G12768 (.A1(W1084), .A2(W1862), .ZN(W2342));
  NOR2X1 G12769 (.A1(W43818), .A2(W38681), .ZN(O17506));
  NOR2X1 G12770 (.A1(W1548), .A2(W11071), .ZN(O17507));
  NOR2X1 G12771 (.A1(W31537), .A2(W6280), .ZN(O17508));
  NOR2X1 G12772 (.A1(W28000), .A2(W20890), .ZN(O17509));
  NOR2X1 G12773 (.A1(W8718), .A2(W37341), .ZN(O17510));
  NOR2X1 G12774 (.A1(W32989), .A2(W40655), .ZN(W48645));
  NOR2X1 G12775 (.A1(W859), .A2(I1027), .ZN(W2344));
  NOR2X1 G12776 (.A1(W8645), .A2(W46664), .ZN(O17518));
  NOR2X1 G12777 (.A1(W17542), .A2(W17395), .ZN(O17550));
  NOR2X1 G12778 (.A1(W9372), .A2(W27295), .ZN(O17520));
  NOR2X1 G12779 (.A1(W1198), .A2(W5911), .ZN(O17521));
  NOR2X1 G12780 (.A1(I1600), .A2(W259), .ZN(W2338));
  NOR2X1 G12781 (.A1(W21211), .A2(W22762), .ZN(W26167));
  NOR2X1 G12782 (.A1(W36125), .A2(W25195), .ZN(O17525));
  NOR2X1 G12783 (.A1(W15444), .A2(W11511), .ZN(W24564));
  NOR2X1 G12784 (.A1(I876), .A2(W572), .ZN(W2332));
  NOR2X1 G12785 (.A1(W1357), .A2(I812), .ZN(W2278));
  NOR2X1 G12786 (.A1(W1474), .A2(W73), .ZN(W2290));
  NOR2X1 G12787 (.A1(W21404), .A2(W20741), .ZN(O17570));
  NOR2X1 G12788 (.A1(W1041), .A2(W435), .ZN(W2288));
  NOR2X1 G12789 (.A1(W2070), .A2(I1399), .ZN(W2287));
  NOR2X1 G12790 (.A1(W38177), .A2(W22419), .ZN(O17572));
  NOR2X1 G12791 (.A1(I426), .A2(W450), .ZN(W2284));
  NOR2X1 G12792 (.A1(W21140), .A2(W12543), .ZN(W26143));
  NOR2X1 G12793 (.A1(I1165), .A2(W1578), .ZN(W2280));
  NOR2X1 G12794 (.A1(W25076), .A2(W34362), .ZN(O17568));
  NOR2X1 G12795 (.A1(W37595), .A2(W32617), .ZN(O17579));
  NOR2X1 G12796 (.A1(I1964), .A2(W747), .ZN(W2276));
  NOR2X1 G12797 (.A1(W46546), .A2(W15757), .ZN(O17580));
  NOR2X1 G12798 (.A1(W6304), .A2(W8736), .ZN(W24587));
  NOR2X1 G12799 (.A1(W1359), .A2(W903), .ZN(W2273));
  NOR2X1 G12800 (.A1(W14868), .A2(W3605), .ZN(W24588));
  NOR2X1 G12801 (.A1(W32915), .A2(W37698), .ZN(O17583));
  NOR2X1 G12802 (.A1(W16194), .A2(I112), .ZN(O3125));
  NOR2X1 G12803 (.A1(W9509), .A2(W24260), .ZN(O3124));
  NOR2X1 G12804 (.A1(I0), .A2(I640), .ZN(W2308));
  NOR2X1 G12805 (.A1(W1781), .A2(I1182), .ZN(W2307));
  NOR2X1 G12806 (.A1(W491), .A2(I735), .ZN(W2306));
  NOR2X1 G12807 (.A1(I494), .A2(W1799), .ZN(W24577));
  NOR2X1 G12808 (.A1(W39314), .A2(W38592), .ZN(O17555));
  NOR2X1 G12809 (.A1(W778), .A2(W1579), .ZN(W24578));
  NOR2X1 G12810 (.A1(W1034), .A2(W47892), .ZN(O17557));
  NOR2X1 G12811 (.A1(W1659), .A2(I1075), .ZN(W1879));
  NOR2X1 G12812 (.A1(W37538), .A2(W28006), .ZN(O17558));
  NOR2X1 G12813 (.A1(W24527), .A2(W21728), .ZN(W26147));
  NOR2X1 G12814 (.A1(W33049), .A2(W45606), .ZN(O17564));
  NOR2X1 G12815 (.A1(I1996), .A2(W1829), .ZN(W2295));
  NOR2X1 G12816 (.A1(W35769), .A2(W3858), .ZN(O17567));
  NOR2X1 G12817 (.A1(I1903), .A2(I1118), .ZN(W2293));
  NOR2X1 G12818 (.A1(W43135), .A2(W27750), .ZN(W48708));
  NOR2X1 G12819 (.A1(W5795), .A2(W16209), .ZN(O3549));
  NOR2X1 G12820 (.A1(W1056), .A2(W423), .ZN(W1465));
  NOR2X1 G12821 (.A1(W46100), .A2(I217), .ZN(O18341));
  NOR2X1 G12822 (.A1(W8830), .A2(W4444), .ZN(O3550));
  NOR2X1 G12823 (.A1(W47624), .A2(W41278), .ZN(O18348));
  NOR2X1 G12824 (.A1(W23903), .A2(W10142), .ZN(W24851));
  NOR2X1 G12825 (.A1(I456), .A2(W900), .ZN(W1460));
  NOR2X1 G12826 (.A1(W40643), .A2(W19880), .ZN(O18352));
  NOR2X1 G12827 (.A1(I124), .A2(W161), .ZN(W1457));
  NOR2X1 G12828 (.A1(W30825), .A2(W39799), .ZN(O18339));
  NOR2X1 G12829 (.A1(I1408), .A2(I1154), .ZN(W1455));
  NOR2X1 G12830 (.A1(W10850), .A2(W15111), .ZN(W24854));
  NOR2X1 G12831 (.A1(W696), .A2(W150), .ZN(W1453));
  NOR2X1 G12832 (.A1(W521), .A2(I1626), .ZN(W1452));
  NOR2X1 G12833 (.A1(W13695), .A2(W2672), .ZN(W24855));
  NOR2X1 G12834 (.A1(W11107), .A2(W52), .ZN(O3218));
  NOR2X1 G12835 (.A1(I137), .A2(I750), .ZN(W1449));
  NOR2X1 G12836 (.A1(W23775), .A2(W9012), .ZN(O18360));
  NOR2X1 G12837 (.A1(W12794), .A2(W21850), .ZN(W25861));
  NOR2X1 G12838 (.A1(I1065), .A2(W30760), .ZN(O18324));
  NOR2X1 G12839 (.A1(W1088), .A2(I1132), .ZN(W1484));
  NOR2X1 G12840 (.A1(W841), .A2(I370), .ZN(W1483));
  NOR2X1 G12841 (.A1(W17731), .A2(W4728), .ZN(O18325));
  NOR2X1 G12842 (.A1(W14622), .A2(W7383), .ZN(O18326));
  NOR2X1 G12843 (.A1(W8474), .A2(W14200), .ZN(O3212));
  NOR2X1 G12844 (.A1(W730), .A2(I1072), .ZN(W1478));
  NOR2X1 G12845 (.A1(W16424), .A2(W12354), .ZN(W24844));
  NOR2X1 G12846 (.A1(I791), .A2(I1162), .ZN(W1446));
  NOR2X1 G12847 (.A1(I519), .A2(I1700), .ZN(W1474));
  NOR2X1 G12848 (.A1(W18959), .A2(W9598), .ZN(O3554));
  NOR2X1 G12849 (.A1(I342), .A2(I246), .ZN(W1472));
  NOR2X1 G12850 (.A1(W14736), .A2(W43511), .ZN(O18336));
  NOR2X1 G12851 (.A1(W22711), .A2(W6298), .ZN(W25853));
  NOR2X1 G12852 (.A1(I632), .A2(W480), .ZN(W1469));
  NOR2X1 G12853 (.A1(W38415), .A2(W30058), .ZN(W49538));
  NOR2X1 G12854 (.A1(W572), .A2(W1259), .ZN(W1418));
  NOR2X1 G12855 (.A1(W830), .A2(I1911), .ZN(W1427));
  NOR2X1 G12856 (.A1(W3592), .A2(W18602), .ZN(W25839));
  NOR2X1 G12857 (.A1(I1958), .A2(W464), .ZN(W1425));
  NOR2X1 G12858 (.A1(W14394), .A2(W34890), .ZN(O18381));
  NOR2X1 G12859 (.A1(W38294), .A2(W48958), .ZN(O18385));
  NOR2X1 G12860 (.A1(W17208), .A2(W19618), .ZN(O3546));
  NOR2X1 G12861 (.A1(W15237), .A2(W13688), .ZN(W24866));
  NOR2X1 G12862 (.A1(W13420), .A2(W17534), .ZN(O3545));
  NOR2X1 G12863 (.A1(W44545), .A2(W7928), .ZN(O18379));
  NOR2X1 G12864 (.A1(W212), .A2(I1181), .ZN(W1417));
  NOR2X1 G12865 (.A1(I270), .A2(W470), .ZN(W1416));
  NOR2X1 G12866 (.A1(W1302), .A2(I1431), .ZN(W1415));
  NOR2X1 G12867 (.A1(W35728), .A2(W24502), .ZN(O18391));
  NOR2X1 G12868 (.A1(W44852), .A2(W25217), .ZN(O18392));
  NOR2X1 G12869 (.A1(W27078), .A2(W18810), .ZN(O18394));
  NOR2X1 G12870 (.A1(W44255), .A2(W12072), .ZN(O18398));
  NOR2X1 G12871 (.A1(W17838), .A2(W35453), .ZN(O18399));
  NOR2X1 G12872 (.A1(I1337), .A2(W453), .ZN(W1437));
  NOR2X1 G12873 (.A1(W48645), .A2(W42423), .ZN(O18362));
  NOR2X1 G12874 (.A1(W11116), .A2(W16977), .ZN(W24858));
  NOR2X1 G12875 (.A1(W23882), .A2(W16069), .ZN(O3548));
  NOR2X1 G12876 (.A1(W39541), .A2(W26748), .ZN(O18367));
  NOR2X1 G12877 (.A1(W17408), .A2(W6033), .ZN(O3219));
  NOR2X1 G12878 (.A1(W2296), .A2(W45232), .ZN(O18369));
  NOR2X1 G12879 (.A1(I398), .A2(I21), .ZN(W1439));
  NOR2X1 G12880 (.A1(W45861), .A2(W49116), .ZN(O18371));
  NOR2X1 G12881 (.A1(W18023), .A2(W15516), .ZN(W25864));
  NOR2X1 G12882 (.A1(W483), .A2(W47584), .ZN(O18373));
  NOR2X1 G12883 (.A1(W1330), .A2(I1282), .ZN(W1435));
  NOR2X1 G12884 (.A1(W8237), .A2(W16497), .ZN(O3547));
  NOR2X1 G12885 (.A1(W35729), .A2(W47626), .ZN(O18377));
  NOR2X1 G12886 (.A1(W7312), .A2(W14136), .ZN(O18378));
  NOR2X1 G12887 (.A1(W274), .A2(W58), .ZN(W1430));
  NOR2X1 G12888 (.A1(I755), .A2(I839), .ZN(W1429));
  NOR2X1 G12889 (.A1(I1835), .A2(W264), .ZN(W1535));
  NOR2X1 G12890 (.A1(W36047), .A2(W13388), .ZN(O18257));
  NOR2X1 G12891 (.A1(W8836), .A2(I11), .ZN(O18258));
  NOR2X1 G12892 (.A1(I793), .A2(W49174), .ZN(O18260));
  NOR2X1 G12893 (.A1(W33205), .A2(W34458), .ZN(O18262));
  NOR2X1 G12894 (.A1(I911), .A2(W899), .ZN(W1540));
  NOR2X1 G12895 (.A1(W12560), .A2(W12720), .ZN(W25879));
  NOR2X1 G12896 (.A1(W798), .A2(I1145), .ZN(W1537));
  NOR2X1 G12897 (.A1(I793), .A2(W288), .ZN(W1536));
  NOR2X1 G12898 (.A1(W32837), .A2(W902), .ZN(O18255));
  NOR2X1 G12899 (.A1(W47285), .A2(W30925), .ZN(O18268));
  NOR2X1 G12900 (.A1(W46121), .A2(W2136), .ZN(O18269));
  NOR2X1 G12901 (.A1(W19135), .A2(I1599), .ZN(W24824));
  NOR2X1 G12902 (.A1(W28647), .A2(W14322), .ZN(O18271));
  NOR2X1 G12903 (.A1(W45286), .A2(W34596), .ZN(O18272));
  NOR2X1 G12904 (.A1(I625), .A2(W401), .ZN(W1529));
  NOR2X1 G12905 (.A1(W22719), .A2(W12909), .ZN(O3204));
  NOR2X1 G12906 (.A1(W322), .A2(I575), .ZN(W1527));
  NOR2X1 G12907 (.A1(I938), .A2(I840), .ZN(W1555));
  NOR2X1 G12908 (.A1(W18038), .A2(W22099), .ZN(W25890));
  NOR2X1 G12909 (.A1(W9339), .A2(W42575), .ZN(O18240));
  NOR2X1 G12910 (.A1(W17777), .A2(W18169), .ZN(W24817));
  NOR2X1 G12911 (.A1(W743), .A2(I1949), .ZN(W1560));
  NOR2X1 G12912 (.A1(W913), .A2(W1465), .ZN(W1559));
  NOR2X1 G12913 (.A1(W12379), .A2(W6809), .ZN(W25889));
  NOR2X1 G12914 (.A1(W13604), .A2(W15139), .ZN(O18244));
  NOR2X1 G12915 (.A1(W46282), .A2(W11972), .ZN(O18245));
  NOR2X1 G12916 (.A1(W21696), .A2(W23461), .ZN(O18275));
  NOR2X1 G12917 (.A1(W1481), .A2(W1167), .ZN(W1553));
  NOR2X1 G12918 (.A1(W3334), .A2(W16696), .ZN(O18248));
  NOR2X1 G12919 (.A1(W37435), .A2(W35655), .ZN(O18250));
  NOR2X1 G12920 (.A1(I1931), .A2(W22144), .ZN(W49448));
  NOR2X1 G12921 (.A1(W796), .A2(W79), .ZN(W1548));
  NOR2X1 G12922 (.A1(I288), .A2(I1774), .ZN(W1547));
  NOR2X1 G12923 (.A1(W944), .A2(W2171), .ZN(W25881));
  NOR2X1 G12924 (.A1(W113), .A2(W31123), .ZN(O18312));
  NOR2X1 G12925 (.A1(W13052), .A2(W9027), .ZN(O18305));
  NOR2X1 G12926 (.A1(I707), .A2(I1414), .ZN(W1502));
  NOR2X1 G12927 (.A1(W23890), .A2(W7519), .ZN(O3210));
  NOR2X1 G12928 (.A1(W180), .A2(I1841), .ZN(W1500));
  NOR2X1 G12929 (.A1(I1739), .A2(W251), .ZN(W1499));
  NOR2X1 G12930 (.A1(W451), .A2(W1036), .ZN(W1498));
  NOR2X1 G12931 (.A1(I1264), .A2(I1423), .ZN(W1496));
  NOR2X1 G12932 (.A1(W9322), .A2(W22554), .ZN(O18310));
  NOR2X1 G12933 (.A1(W6690), .A2(I1457), .ZN(O3209));
  NOR2X1 G12934 (.A1(W13059), .A2(W24156), .ZN(O18313));
  NOR2X1 G12935 (.A1(I572), .A2(I1463), .ZN(W1492));
  NOR2X1 G12936 (.A1(W44820), .A2(W996), .ZN(O18314));
  NOR2X1 G12937 (.A1(W9613), .A2(W3206), .ZN(W24840));
  NOR2X1 G12938 (.A1(W12773), .A2(W7119), .ZN(O18320));
  NOR2X1 G12939 (.A1(W42629), .A2(W496), .ZN(O18321));
  NOR2X1 G12940 (.A1(W1163), .A2(W505), .ZN(W1487));
  NOR2X1 G12941 (.A1(W29503), .A2(W16090), .ZN(O18287));
  NOR2X1 G12942 (.A1(W22529), .A2(W21639), .ZN(O18276));
  NOR2X1 G12943 (.A1(W21437), .A2(W45413), .ZN(O18278));
  NOR2X1 G12944 (.A1(W1060), .A2(W937), .ZN(W1523));
  NOR2X1 G12945 (.A1(W16270), .A2(W21293), .ZN(W25878));
  NOR2X1 G12946 (.A1(W9811), .A2(W15501), .ZN(W24828));
  NOR2X1 G12947 (.A1(W5736), .A2(W7461), .ZN(O18283));
  NOR2X1 G12948 (.A1(W19609), .A2(W30773), .ZN(O18284));
  NOR2X1 G12949 (.A1(W16892), .A2(W20636), .ZN(O3206));
  NOR2X1 G12950 (.A1(I28), .A2(I1980), .ZN(W1409));
  NOR2X1 G12951 (.A1(W20256), .A2(W7360), .ZN(W24831));
  NOR2X1 G12952 (.A1(W20965), .A2(W4307), .ZN(O3207));
  NOR2X1 G12953 (.A1(W22537), .A2(W18125), .ZN(O3561));
  NOR2X1 G12954 (.A1(W12390), .A2(W45841), .ZN(O18295));
  NOR2X1 G12955 (.A1(W47854), .A2(W5673), .ZN(W49495));
  NOR2X1 G12956 (.A1(W39304), .A2(W37551), .ZN(O18299));
  NOR2X1 G12957 (.A1(W7249), .A2(W43012), .ZN(O18301));
  NOR2X1 G12958 (.A1(W8142), .A2(W26604), .ZN(O18485));
  NOR2X1 G12959 (.A1(W23700), .A2(W22217), .ZN(O18479));
  NOR2X1 G12960 (.A1(W42534), .A2(W20920), .ZN(O18480));
  NOR2X1 G12961 (.A1(W1251), .A2(W1130), .ZN(W1311));
  NOR2X1 G12962 (.A1(I930), .A2(I1646), .ZN(W1310));
  NOR2X1 G12963 (.A1(W21089), .A2(W16482), .ZN(O18481));
  NOR2X1 G12964 (.A1(W38576), .A2(W34275), .ZN(O18484));
  NOR2X1 G12965 (.A1(I1161), .A2(W1243), .ZN(W1307));
  NOR2X1 G12966 (.A1(I995), .A2(I861), .ZN(W1306));
  NOR2X1 G12967 (.A1(W14751), .A2(W7017), .ZN(O3234));
  NOR2X1 G12968 (.A1(W464), .A2(I1535), .ZN(W1304));
  NOR2X1 G12969 (.A1(W5551), .A2(W24123), .ZN(O18487));
  NOR2X1 G12970 (.A1(W42254), .A2(W28289), .ZN(O18491));
  NOR2X1 G12971 (.A1(I11), .A2(I39), .ZN(W1301));
  NOR2X1 G12972 (.A1(W48695), .A2(W2397), .ZN(O18493));
  NOR2X1 G12973 (.A1(W49029), .A2(W4437), .ZN(O18496));
  NOR2X1 G12974 (.A1(W3131), .A2(W11877), .ZN(O3236));
  NOR2X1 G12975 (.A1(W22435), .A2(W10140), .ZN(W25790));
  NOR2X1 G12976 (.A1(W147), .A2(I1697), .ZN(W1322));
  NOR2X1 G12977 (.A1(I676), .A2(I348), .ZN(W1330));
  NOR2X1 G12978 (.A1(W1064), .A2(I462), .ZN(W1329));
  NOR2X1 G12979 (.A1(W42773), .A2(W39667), .ZN(O18470));
  NOR2X1 G12980 (.A1(I1570), .A2(I1988), .ZN(W1327));
  NOR2X1 G12981 (.A1(W3861), .A2(W893), .ZN(W49678));
  NOR2X1 G12982 (.A1(I1895), .A2(W438), .ZN(W1325));
  NOR2X1 G12983 (.A1(W23247), .A2(W14273), .ZN(W24897));
  NOR2X1 G12984 (.A1(W404), .A2(I0), .ZN(W1323));
  NOR2X1 G12985 (.A1(W26017), .A2(W30514), .ZN(O18499));
  NOR2X1 G12986 (.A1(W42276), .A2(W4044), .ZN(O18473));
  NOR2X1 G12987 (.A1(W18716), .A2(W40923), .ZN(O18474));
  NOR2X1 G12988 (.A1(W19290), .A2(W20540), .ZN(W24898));
  NOR2X1 G12989 (.A1(I1067), .A2(I609), .ZN(W1318));
  NOR2X1 G12990 (.A1(W5659), .A2(W12405), .ZN(W25801));
  NOR2X1 G12991 (.A1(W190), .A2(I1928), .ZN(W1316));
  NOR2X1 G12992 (.A1(W6771), .A2(W33), .ZN(W25798));
  NOR2X1 G12993 (.A1(W1194), .A2(W728), .ZN(W1266));
  NOR2X1 G12994 (.A1(W23074), .A2(W17901), .ZN(W24913));
  NOR2X1 G12995 (.A1(W11018), .A2(W2039), .ZN(W24914));
  NOR2X1 G12996 (.A1(W10090), .A2(W11775), .ZN(O18523));
  NOR2X1 G12997 (.A1(I759), .A2(I799), .ZN(W1272));
  NOR2X1 G12998 (.A1(I918), .A2(I1738), .ZN(W1271));
  NOR2X1 G12999 (.A1(W70), .A2(I1557), .ZN(W1269));
  NOR2X1 G13000 (.A1(W10565), .A2(W6308), .ZN(O3529));
  NOR2X1 G13001 (.A1(I169), .A2(I1866), .ZN(W1267));
  NOR2X1 G13002 (.A1(W24555), .A2(W4672), .ZN(W25787));
  NOR2X1 G13003 (.A1(W22352), .A2(W12891), .ZN(O18527));
  NOR2X1 G13004 (.A1(I1620), .A2(I613), .ZN(W1264));
  NOR2X1 G13005 (.A1(W44907), .A2(W10059), .ZN(O18528));
  NOR2X1 G13006 (.A1(W13289), .A2(W17415), .ZN(W25783));
  NOR2X1 G13007 (.A1(W8961), .A2(W3071), .ZN(O3242));
  NOR2X1 G13008 (.A1(W385), .A2(I541), .ZN(W1260));
  NOR2X1 G13009 (.A1(I1171), .A2(W628), .ZN(W1259));
  NOR2X1 G13010 (.A1(W28374), .A2(W11699), .ZN(O18513));
  NOR2X1 G13011 (.A1(W15174), .A2(W20375), .ZN(W25789));
  NOR2X1 G13012 (.A1(W804), .A2(W44166), .ZN(O18503));
  NOR2X1 G13013 (.A1(W8397), .A2(W1781), .ZN(O18504));
  NOR2X1 G13014 (.A1(W5729), .A2(W46091), .ZN(O18505));
  NOR2X1 G13015 (.A1(W17316), .A2(W44393), .ZN(W49715));
  NOR2X1 G13016 (.A1(W17920), .A2(I1708), .ZN(W24906));
  NOR2X1 G13017 (.A1(W6393), .A2(W10238), .ZN(O18511));
  NOR2X1 G13018 (.A1(I839), .A2(W1991), .ZN(W24907));
  NOR2X1 G13019 (.A1(W21066), .A2(W19718), .ZN(W25802));
  NOR2X1 G13020 (.A1(I1163), .A2(W193), .ZN(W1285));
  NOR2X1 G13021 (.A1(W593), .A2(I1473), .ZN(W1284));
  NOR2X1 G13022 (.A1(W23983), .A2(W13617), .ZN(W24908));
  NOR2X1 G13023 (.A1(I1888), .A2(W642), .ZN(W1282));
  NOR2X1 G13024 (.A1(W14687), .A2(W8269), .ZN(O3239));
  NOR2X1 G13025 (.A1(W1111), .A2(I44), .ZN(W1280));
  NOR2X1 G13026 (.A1(I1997), .A2(I1519), .ZN(W1278));
  NOR2X1 G13027 (.A1(W38034), .A2(W39918), .ZN(O18431));
  NOR2X1 G13028 (.A1(W9596), .A2(W13593), .ZN(O3541));
  NOR2X1 G13029 (.A1(W21673), .A2(I1461), .ZN(W24876));
  NOR2X1 G13030 (.A1(W4235), .A2(W16558), .ZN(O3225));
  NOR2X1 G13031 (.A1(W1014), .A2(W13218), .ZN(O3540));
  NOR2X1 G13032 (.A1(W1322), .A2(W927), .ZN(W1382));
  NOR2X1 G13033 (.A1(W233), .A2(I700), .ZN(W1381));
  NOR2X1 G13034 (.A1(I79), .A2(W1276), .ZN(W1380));
  NOR2X1 G13035 (.A1(W10581), .A2(W23762), .ZN(W24881));
  NOR2X1 G13036 (.A1(I700), .A2(W48), .ZN(W1389));
  NOR2X1 G13037 (.A1(I316), .A2(W961), .ZN(W1377));
  NOR2X1 G13038 (.A1(W17212), .A2(W36095), .ZN(O18433));
  NOR2X1 G13039 (.A1(W32099), .A2(W15969), .ZN(O18434));
  NOR2X1 G13040 (.A1(W15220), .A2(W997), .ZN(O3539));
  NOR2X1 G13041 (.A1(W14982), .A2(W4623), .ZN(O18439));
  NOR2X1 G13042 (.A1(W434), .A2(I1250), .ZN(W1372));
  NOR2X1 G13043 (.A1(W16790), .A2(W9810), .ZN(W25815));
  NOR2X1 G13044 (.A1(W11681), .A2(W748), .ZN(O18442));
  NOR2X1 G13045 (.A1(W52), .A2(I1472), .ZN(W1399));
  NOR2X1 G13046 (.A1(W1040), .A2(I482), .ZN(O12));
  NOR2X1 G13047 (.A1(W6084), .A2(W4727), .ZN(O18402));
  NOR2X1 G13048 (.A1(W33231), .A2(W30070), .ZN(O18403));
  NOR2X1 G13049 (.A1(I766), .A2(I136), .ZN(W1404));
  NOR2X1 G13050 (.A1(W14046), .A2(W11021), .ZN(W25830));
  NOR2X1 G13051 (.A1(W29887), .A2(W267), .ZN(O18407));
  NOR2X1 G13052 (.A1(W13233), .A2(W21614), .ZN(O3543));
  NOR2X1 G13053 (.A1(W21765), .A2(W24660), .ZN(O3223));
  NOR2X1 G13054 (.A1(W38956), .A2(W21736), .ZN(O18444));
  NOR2X1 G13055 (.A1(W24051), .A2(W41401), .ZN(O18413));
  NOR2X1 G13056 (.A1(I587), .A2(I962), .ZN(W1397));
  NOR2X1 G13057 (.A1(W758), .A2(I1665), .ZN(W1396));
  NOR2X1 G13058 (.A1(I842), .A2(W500), .ZN(W1395));
  NOR2X1 G13059 (.A1(I137), .A2(I686), .ZN(W1393));
  NOR2X1 G13060 (.A1(W8554), .A2(W21898), .ZN(W25824));
  NOR2X1 G13061 (.A1(W19520), .A2(W105), .ZN(O18416));
  NOR2X1 G13062 (.A1(W431), .A2(I1872), .ZN(W1340));
  NOR2X1 G13063 (.A1(I1177), .A2(W1355), .ZN(W25809));
  NOR2X1 G13064 (.A1(W992), .A2(W1056), .ZN(W1348));
  NOR2X1 G13065 (.A1(W1145), .A2(W931), .ZN(W1347));
  NOR2X1 G13066 (.A1(W12899), .A2(W5931), .ZN(O18461));
  NOR2X1 G13067 (.A1(I1659), .A2(W251), .ZN(W1345));
  NOR2X1 G13068 (.A1(W24228), .A2(I1075), .ZN(W25807));
  NOR2X1 G13069 (.A1(I70), .A2(I1429), .ZN(W1342));
  NOR2X1 G13070 (.A1(W1578), .A2(W14814), .ZN(O3535));
  NOR2X1 G13071 (.A1(W21715), .A2(W5697), .ZN(W24889));
  NOR2X1 G13072 (.A1(I746), .A2(W1073), .ZN(W1339));
  NOR2X1 G13073 (.A1(W793), .A2(W1205), .ZN(W1338));
  NOR2X1 G13074 (.A1(W23265), .A2(W19527), .ZN(O18464));
  NOR2X1 G13075 (.A1(W9), .A2(W948), .ZN(W1336));
  NOR2X1 G13076 (.A1(W16165), .A2(W1790), .ZN(W25804));
  NOR2X1 G13077 (.A1(W716), .A2(I272), .ZN(W1333));
  NOR2X1 G13078 (.A1(W1172), .A2(W24998), .ZN(O18468));
  NOR2X1 G13079 (.A1(I452), .A2(W39313), .ZN(O18453));
  NOR2X1 G13080 (.A1(W23116), .A2(W2987), .ZN(O18445));
  NOR2X1 G13081 (.A1(W42454), .A2(W30980), .ZN(O18447));
  NOR2X1 G13082 (.A1(W5209), .A2(W15089), .ZN(W25814));
  NOR2X1 G13083 (.A1(W18576), .A2(W20362), .ZN(O18449));
  NOR2X1 G13084 (.A1(I524), .A2(W1202), .ZN(W1364));
  NOR2X1 G13085 (.A1(I319), .A2(W19413), .ZN(W25813));
  NOR2X1 G13086 (.A1(W10368), .A2(W23982), .ZN(O18451));
  NOR2X1 G13087 (.A1(I987), .A2(I1887), .ZN(W1360));
  NOR2X1 G13088 (.A1(W22950), .A2(W25454), .ZN(W25892));
  NOR2X1 G13089 (.A1(W24603), .A2(W7837), .ZN(O3230));
  NOR2X1 G13090 (.A1(W713), .A2(I923), .ZN(W1357));
  NOR2X1 G13091 (.A1(W91), .A2(W742), .ZN(W1356));
  NOR2X1 G13092 (.A1(W584), .A2(W8), .ZN(W1355));
  NOR2X1 G13093 (.A1(W358), .A2(I1282), .ZN(W1353));
  NOR2X1 G13094 (.A1(I613), .A2(W1012), .ZN(W1352));
  NOR2X1 G13095 (.A1(W32290), .A2(W26781), .ZN(O18456));
  NOR2X1 G13096 (.A1(W8317), .A2(W9104), .ZN(W24746));
  NOR2X1 G13097 (.A1(W21587), .A2(W8310), .ZN(W25971));
  NOR2X1 G13098 (.A1(W14232), .A2(W46119), .ZN(O18039));
  NOR2X1 G13099 (.A1(W4475), .A2(W2679), .ZN(O18042));
  NOR2X1 G13100 (.A1(W14255), .A2(W40001), .ZN(O18045));
  NOR2X1 G13101 (.A1(W457), .A2(I1075), .ZN(W1772));
  NOR2X1 G13102 (.A1(W2881), .A2(W46233), .ZN(O18047));
  NOR2X1 G13103 (.A1(W417), .A2(I46), .ZN(W1770));
  NOR2X1 G13104 (.A1(I895), .A2(W895), .ZN(W1769));
  NOR2X1 G13105 (.A1(W828), .A2(I1332), .ZN(W1777));
  NOR2X1 G13106 (.A1(I711), .A2(I1728), .ZN(W1767));
  NOR2X1 G13107 (.A1(W24376), .A2(W4826), .ZN(O3180));
  NOR2X1 G13108 (.A1(W731), .A2(W437), .ZN(W1765));
  NOR2X1 G13109 (.A1(I1415), .A2(W5832), .ZN(W24748));
  NOR2X1 G13110 (.A1(W18675), .A2(W4419), .ZN(W25970));
  NOR2X1 G13111 (.A1(W4966), .A2(I249), .ZN(W25969));
  NOR2X1 G13112 (.A1(W32276), .A2(W46931), .ZN(O18053));
  NOR2X1 G13113 (.A1(I1953), .A2(W1382), .ZN(W49237));
  NOR2X1 G13114 (.A1(W41877), .A2(W3214), .ZN(W49209));
  NOR2X1 G13115 (.A1(W2810), .A2(W24343), .ZN(O3176));
  NOR2X1 G13116 (.A1(W25222), .A2(W42823), .ZN(O18019));
  NOR2X1 G13117 (.A1(W39197), .A2(W23908), .ZN(W49199));
  NOR2X1 G13118 (.A1(W3462), .A2(W31041), .ZN(O18021));
  NOR2X1 G13119 (.A1(W1751), .A2(I1702), .ZN(W1794));
  NOR2X1 G13120 (.A1(W26390), .A2(W3618), .ZN(O18022));
  NOR2X1 G13121 (.A1(W6553), .A2(W13178), .ZN(O3591));
  NOR2X1 G13122 (.A1(W42367), .A2(W13077), .ZN(O18027));
  NOR2X1 G13123 (.A1(W1658), .A2(W1710), .ZN(W1759));
  NOR2X1 G13124 (.A1(W1021), .A2(W373), .ZN(W1787));
  NOR2X1 G13125 (.A1(W3346), .A2(W48936), .ZN(O18030));
  NOR2X1 G13126 (.A1(W650), .A2(I426), .ZN(W1784));
  NOR2X1 G13127 (.A1(W18399), .A2(W200), .ZN(W25974));
  NOR2X1 G13128 (.A1(W31426), .A2(W6169), .ZN(O18035));
  NOR2X1 G13129 (.A1(I29), .A2(W1216), .ZN(W1779));
  NOR2X1 G13130 (.A1(W66), .A2(W1176), .ZN(W1778));
  NOR2X1 G13131 (.A1(W15893), .A2(W314), .ZN(O18083));
  NOR2X1 G13132 (.A1(W1656), .A2(W898), .ZN(W1740));
  NOR2X1 G13133 (.A1(W474), .A2(I316), .ZN(W1738));
  NOR2X1 G13134 (.A1(W4493), .A2(W30771), .ZN(O18076));
  NOR2X1 G13135 (.A1(W5044), .A2(I334), .ZN(O18077));
  NOR2X1 G13136 (.A1(W21436), .A2(W2011), .ZN(O18080));
  NOR2X1 G13137 (.A1(I1532), .A2(W796), .ZN(W1733));
  NOR2X1 G13138 (.A1(W45776), .A2(W21498), .ZN(O18082));
  NOR2X1 G13139 (.A1(I1130), .A2(I1775), .ZN(W1731));
  NOR2X1 G13140 (.A1(I1243), .A2(I1053), .ZN(W1741));
  NOR2X1 G13141 (.A1(W1664), .A2(I1076), .ZN(W1729));
  NOR2X1 G13142 (.A1(W23383), .A2(W31877), .ZN(O18084));
  NOR2X1 G13143 (.A1(W472), .A2(I1459), .ZN(W1727));
  NOR2X1 G13144 (.A1(W4380), .A2(W31528), .ZN(O18090));
  NOR2X1 G13145 (.A1(I712), .A2(I658), .ZN(W1724));
  NOR2X1 G13146 (.A1(W21557), .A2(W19428), .ZN(W25956));
  NOR2X1 G13147 (.A1(W23810), .A2(W19950), .ZN(W25955));
  NOR2X1 G13148 (.A1(W11678), .A2(W12877), .ZN(W24753));
  NOR2X1 G13149 (.A1(W6516), .A2(W37042), .ZN(O18054));
  NOR2X1 G13150 (.A1(I1242), .A2(I1526), .ZN(W1757));
  NOR2X1 G13151 (.A1(W22566), .A2(W23117), .ZN(O18055));
  NOR2X1 G13152 (.A1(W14929), .A2(W12790), .ZN(W25968));
  NOR2X1 G13153 (.A1(I1654), .A2(I338), .ZN(W1753));
  NOR2X1 G13154 (.A1(W1035), .A2(W783), .ZN(W1752));
  NOR2X1 G13155 (.A1(I870), .A2(I1804), .ZN(W1751));
  NOR2X1 G13156 (.A1(W46443), .A2(W24134), .ZN(O18058));
  NOR2X1 G13157 (.A1(W10008), .A2(W7062), .ZN(O3175));
  NOR2X1 G13158 (.A1(W14327), .A2(W10519), .ZN(O18065));
  NOR2X1 G13159 (.A1(W27617), .A2(W6973), .ZN(O18069));
  NOR2X1 G13160 (.A1(W13392), .A2(I554), .ZN(O18071));
  NOR2X1 G13161 (.A1(W1139), .A2(W1207), .ZN(W1745));
  NOR2X1 G13162 (.A1(W25744), .A2(W17551), .ZN(O18072));
  NOR2X1 G13163 (.A1(I1306), .A2(W14027), .ZN(O3183));
  NOR2X1 G13164 (.A1(W4069), .A2(W18144), .ZN(O3589));
  NOR2X1 G13165 (.A1(I122), .A2(I156), .ZN(W1850));
  NOR2X1 G13166 (.A1(W20631), .A2(W9159), .ZN(O17955));
  NOR2X1 G13167 (.A1(W50), .A2(I969), .ZN(W1857));
  NOR2X1 G13168 (.A1(W38708), .A2(W42307), .ZN(O17957));
  NOR2X1 G13169 (.A1(W14877), .A2(W14544), .ZN(O3171));
  NOR2X1 G13170 (.A1(W21853), .A2(W40673), .ZN(O17959));
  NOR2X1 G13171 (.A1(W10757), .A2(W16874), .ZN(O3600));
  NOR2X1 G13172 (.A1(W11645), .A2(W9105), .ZN(W26005));
  NOR2X1 G13173 (.A1(I1452), .A2(W316), .ZN(W1851));
  NOR2X1 G13174 (.A1(I337), .A2(I630), .ZN(W1859));
  NOR2X1 G13175 (.A1(I1608), .A2(W1063), .ZN(W1849));
  NOR2X1 G13176 (.A1(W1113), .A2(W1327), .ZN(W1848));
  NOR2X1 G13177 (.A1(W32041), .A2(W16816), .ZN(O17964));
  NOR2X1 G13178 (.A1(W30333), .A2(W30752), .ZN(O17966));
  NOR2X1 G13179 (.A1(W34384), .A2(W9289), .ZN(O17967));
  NOR2X1 G13180 (.A1(I1824), .A2(W22073), .ZN(O17969));
  NOR2X1 G13181 (.A1(W42833), .A2(W283), .ZN(O17970));
  NOR2X1 G13182 (.A1(W1460), .A2(W462), .ZN(W1842));
  NOR2X1 G13183 (.A1(W25730), .A2(W24790), .ZN(O17945));
  NOR2X1 G13184 (.A1(W939), .A2(W500), .ZN(W1878));
  NOR2X1 G13185 (.A1(I824), .A2(I1875), .ZN(W1876));
  NOR2X1 G13186 (.A1(I993), .A2(I431), .ZN(W1875));
  NOR2X1 G13187 (.A1(W41829), .A2(W29087), .ZN(O17940));
  NOR2X1 G13188 (.A1(W48669), .A2(W10495), .ZN(W49116));
  NOR2X1 G13189 (.A1(I1506), .A2(I1505), .ZN(W1872));
  NOR2X1 G13190 (.A1(I446), .A2(W139), .ZN(W1871));
  NOR2X1 G13191 (.A1(W14848), .A2(W17763), .ZN(W24713));
  NOR2X1 G13192 (.A1(W651), .A2(W539), .ZN(W1841));
  NOR2X1 G13193 (.A1(I764), .A2(I1174), .ZN(W1868));
  NOR2X1 G13194 (.A1(W42578), .A2(W46422), .ZN(O17947));
  NOR2X1 G13195 (.A1(W6254), .A2(W17918), .ZN(O3602));
  NOR2X1 G13196 (.A1(I567), .A2(W746), .ZN(W1864));
  NOR2X1 G13197 (.A1(W25276), .A2(W17592), .ZN(O17951));
  NOR2X1 G13198 (.A1(W8274), .A2(W41671), .ZN(O17952));
  NOR2X1 G13199 (.A1(W14210), .A2(W18380), .ZN(W26008));
  NOR2X1 G13200 (.A1(W1005), .A2(W120), .ZN(W1808));
  NOR2X1 G13201 (.A1(W377), .A2(W45559), .ZN(W49174));
  NOR2X1 G13202 (.A1(W20961), .A2(W38351), .ZN(W49175));
  NOR2X1 G13203 (.A1(W19507), .A2(W24299), .ZN(W25987));
  NOR2X1 G13204 (.A1(W3740), .A2(W12290), .ZN(W49178));
  NOR2X1 G13205 (.A1(W801), .A2(W20795), .ZN(W24732));
  NOR2X1 G13206 (.A1(W994), .A2(I1163), .ZN(W1811));
  NOR2X1 G13207 (.A1(W624), .A2(W22), .ZN(W1810));
  NOR2X1 G13208 (.A1(W208), .A2(I1880), .ZN(W1809));
  NOR2X1 G13209 (.A1(W18633), .A2(W25369), .ZN(O3594));
  NOR2X1 G13210 (.A1(W1754), .A2(W1237), .ZN(W1807));
  NOR2X1 G13211 (.A1(I646), .A2(I1161), .ZN(W1806));
  NOR2X1 G13212 (.A1(W11774), .A2(W17785), .ZN(W25986));
  NOR2X1 G13213 (.A1(W14902), .A2(W41012), .ZN(O18010));
  NOR2X1 G13214 (.A1(I1695), .A2(I218), .ZN(W1803));
  NOR2X1 G13215 (.A1(W4658), .A2(W22071), .ZN(W24734));
  NOR2X1 G13216 (.A1(W396), .A2(W1189), .ZN(W1800));
  NOR2X1 G13217 (.A1(I690), .A2(W512), .ZN(W1829));
  NOR2X1 G13218 (.A1(W4121), .A2(W22601), .ZN(W24721));
  NOR2X1 G13219 (.A1(W12648), .A2(W28498), .ZN(O17973));
  NOR2X1 G13220 (.A1(W19279), .A2(W11237), .ZN(W26002));
  NOR2X1 G13221 (.A1(W197), .A2(I160), .ZN(W1837));
  NOR2X1 G13222 (.A1(W33489), .A2(W33774), .ZN(O17983));
  NOR2X1 G13223 (.A1(I1289), .A2(W804), .ZN(W1833));
  NOR2X1 G13224 (.A1(W41926), .A2(W26783), .ZN(O17985));
  NOR2X1 G13225 (.A1(W28723), .A2(W25810), .ZN(O17988));
  NOR2X1 G13226 (.A1(W5354), .A2(I1938), .ZN(O18094));
  NOR2X1 G13227 (.A1(W1155), .A2(W1), .ZN(W1828));
  NOR2X1 G13228 (.A1(W17923), .A2(W4667), .ZN(O17991));
  NOR2X1 G13229 (.A1(W706), .A2(W1287), .ZN(W1824));
  NOR2X1 G13230 (.A1(W534), .A2(I998), .ZN(W1823));
  NOR2X1 G13231 (.A1(W12086), .A2(W33281), .ZN(O17994));
  NOR2X1 G13232 (.A1(I32), .A2(W56), .ZN(W1819));
  NOR2X1 G13233 (.A1(W223), .A2(W1747), .ZN(W1818));
  NOR2X1 G13234 (.A1(W20321), .A2(W40529), .ZN(O18187));
  NOR2X1 G13235 (.A1(I376), .A2(I1755), .ZN(W1621));
  NOR2X1 G13236 (.A1(W8934), .A2(W6015), .ZN(O18181));
  NOR2X1 G13237 (.A1(I1544), .A2(I509), .ZN(W1619));
  NOR2X1 G13238 (.A1(W885), .A2(W193), .ZN(W1618));
  NOR2X1 G13239 (.A1(I1341), .A2(I1873), .ZN(W1617));
  NOR2X1 G13240 (.A1(W25682), .A2(W21860), .ZN(W25910));
  NOR2X1 G13241 (.A1(W2629), .A2(W39942), .ZN(O18185));
  NOR2X1 G13242 (.A1(W29936), .A2(W11108), .ZN(O18186));
  NOR2X1 G13243 (.A1(W689), .A2(W478), .ZN(W1622));
  NOR2X1 G13244 (.A1(W1149), .A2(W1539), .ZN(W1612));
  NOR2X1 G13245 (.A1(W826), .A2(W186), .ZN(W1609));
  NOR2X1 G13246 (.A1(I1245), .A2(I1795), .ZN(W1608));
  NOR2X1 G13247 (.A1(W3020), .A2(W35348), .ZN(O18190));
  NOR2X1 G13248 (.A1(W40339), .A2(W34237), .ZN(O18191));
  NOR2X1 G13249 (.A1(I1113), .A2(I1208), .ZN(W1602));
  NOR2X1 G13250 (.A1(W509), .A2(I1005), .ZN(W1601));
  NOR2X1 G13251 (.A1(W7424), .A2(W17854), .ZN(W25903));
  NOR2X1 G13252 (.A1(W13121), .A2(W26753), .ZN(O18176));
  NOR2X1 G13253 (.A1(W11691), .A2(I1932), .ZN(O18168));
  NOR2X1 G13254 (.A1(W44698), .A2(W24341), .ZN(O18169));
  NOR2X1 G13255 (.A1(W999), .A2(W1020), .ZN(W1639));
  NOR2X1 G13256 (.A1(I1281), .A2(I501), .ZN(W1638));
  NOR2X1 G13257 (.A1(I1123), .A2(I1665), .ZN(W1636));
  NOR2X1 G13258 (.A1(W7140), .A2(W4820), .ZN(W25915));
  NOR2X1 G13259 (.A1(I354), .A2(W16040), .ZN(W25913));
  NOR2X1 G13260 (.A1(I1979), .A2(I1980), .ZN(W1632));
  NOR2X1 G13261 (.A1(W40885), .A2(W9819), .ZN(O18197));
  NOR2X1 G13262 (.A1(I1649), .A2(W8531), .ZN(W24795));
  NOR2X1 G13263 (.A1(W960), .A2(I744), .ZN(W1628));
  NOR2X1 G13264 (.A1(W13009), .A2(W28530), .ZN(O18178));
  NOR2X1 G13265 (.A1(W34591), .A2(W3146), .ZN(O18179));
  NOR2X1 G13266 (.A1(W8607), .A2(W3859), .ZN(W24796));
  NOR2X1 G13267 (.A1(I51), .A2(W140), .ZN(W1624));
  NOR2X1 G13268 (.A1(I677), .A2(I236), .ZN(W1623));
  NOR2X1 G13269 (.A1(W1358), .A2(W6237), .ZN(W25893));
  NOR2X1 G13270 (.A1(W751), .A2(I1307), .ZN(W1580));
  NOR2X1 G13271 (.A1(W16967), .A2(W44993), .ZN(O18223));
  NOR2X1 G13272 (.A1(W26919), .A2(I335), .ZN(O18224));
  NOR2X1 G13273 (.A1(W185), .A2(W97), .ZN(W1577));
  NOR2X1 G13274 (.A1(W36666), .A2(W8458), .ZN(O18225));
  NOR2X1 G13275 (.A1(W15479), .A2(W48969), .ZN(O18227));
  NOR2X1 G13276 (.A1(W7743), .A2(W22490), .ZN(O18229));
  NOR2X1 G13277 (.A1(I243), .A2(W21380), .ZN(O3567));
  NOR2X1 G13278 (.A1(W33188), .A2(W10666), .ZN(O18222));
  NOR2X1 G13279 (.A1(W1440), .A2(I743), .ZN(W1571));
  NOR2X1 G13280 (.A1(W19262), .A2(I283), .ZN(W24813));
  NOR2X1 G13281 (.A1(W213), .A2(I1323), .ZN(W1569));
  NOR2X1 G13282 (.A1(I1333), .A2(W1119), .ZN(W1568));
  NOR2X1 G13283 (.A1(W43914), .A2(W16081), .ZN(W49426));
  NOR2X1 G13284 (.A1(W1518), .A2(W705), .ZN(W1566));
  NOR2X1 G13285 (.A1(W24536), .A2(W7751), .ZN(W24814));
  NOR2X1 G13286 (.A1(W10926), .A2(W3413), .ZN(W24808));
  NOR2X1 G13287 (.A1(I242), .A2(I1707), .ZN(W1598));
  NOR2X1 G13288 (.A1(W4900), .A2(W26126), .ZN(O18198));
  NOR2X1 G13289 (.A1(W37703), .A2(I1815), .ZN(O18199));
  NOR2X1 G13290 (.A1(W9961), .A2(W17106), .ZN(W24804));
  NOR2X1 G13291 (.A1(W24883), .A2(W6405), .ZN(W25901));
  NOR2X1 G13292 (.A1(W4324), .A2(W9263), .ZN(O3569));
  NOR2X1 G13293 (.A1(W24732), .A2(W12950), .ZN(W25899));
  NOR2X1 G13294 (.A1(W21650), .A2(W49199), .ZN(O18212));
  NOR2X1 G13295 (.A1(I1568), .A2(I544), .ZN(W1642));
  NOR2X1 G13296 (.A1(I1881), .A2(W692), .ZN(W1589));
  NOR2X1 G13297 (.A1(W14216), .A2(W10731), .ZN(O18215));
  NOR2X1 G13298 (.A1(W24473), .A2(W43104), .ZN(O18216));
  NOR2X1 G13299 (.A1(W43), .A2(W1365), .ZN(W1585));
  NOR2X1 G13300 (.A1(W14023), .A2(W20902), .ZN(W24810));
  NOR2X1 G13301 (.A1(W37408), .A2(W16956), .ZN(O18220));
  NOR2X1 G13302 (.A1(W38970), .A2(W22560), .ZN(O18221));
  NOR2X1 G13303 (.A1(W29440), .A2(W12290), .ZN(O18123));
  NOR2X1 G13304 (.A1(W1601), .A2(W375), .ZN(W1701));
  NOR2X1 G13305 (.A1(W440), .A2(W42), .ZN(W1700));
  NOR2X1 G13306 (.A1(W1159), .A2(W23740), .ZN(W25949));
  NOR2X1 G13307 (.A1(W13097), .A2(W40340), .ZN(O18116));
  NOR2X1 G13308 (.A1(W14845), .A2(W36016), .ZN(O18118));
  NOR2X1 G13309 (.A1(W3247), .A2(W20577), .ZN(W24766));
  NOR2X1 G13310 (.A1(W5838), .A2(W11873), .ZN(W24767));
  NOR2X1 G13311 (.A1(W529), .A2(I94), .ZN(W1693));
  NOR2X1 G13312 (.A1(I1774), .A2(W620), .ZN(W1703));
  NOR2X1 G13313 (.A1(W907), .A2(I531), .ZN(W1691));
  NOR2X1 G13314 (.A1(W22), .A2(I671), .ZN(W1690));
  NOR2X1 G13315 (.A1(W4589), .A2(W4658), .ZN(O18124));
  NOR2X1 G13316 (.A1(W444), .A2(I250), .ZN(W1688));
  NOR2X1 G13317 (.A1(W48739), .A2(W26340), .ZN(O18125));
  NOR2X1 G13318 (.A1(W8769), .A2(W8958), .ZN(W25947));
  NOR2X1 G13319 (.A1(W1764), .A2(W27480), .ZN(O18129));
  NOR2X1 G13320 (.A1(W4981), .A2(W16818), .ZN(O18130));
  NOR2X1 G13321 (.A1(W22836), .A2(W27608), .ZN(O18102));
  NOR2X1 G13322 (.A1(W27178), .A2(W36926), .ZN(O18095));
  NOR2X1 G13323 (.A1(W26577), .A2(W2258), .ZN(O18096));
  NOR2X1 G13324 (.A1(W30222), .A2(W6019), .ZN(O18097));
  NOR2X1 G13325 (.A1(I1743), .A2(I1684), .ZN(W1717));
  NOR2X1 G13326 (.A1(W1303), .A2(W1453), .ZN(W1716));
  NOR2X1 G13327 (.A1(W11843), .A2(I578), .ZN(O18100));
  NOR2X1 G13328 (.A1(W38384), .A2(W38767), .ZN(O18101));
  NOR2X1 G13329 (.A1(W248), .A2(I1306), .ZN(W1713));
  NOR2X1 G13330 (.A1(I980), .A2(I264), .ZN(W1682));
  NOR2X1 G13331 (.A1(I1588), .A2(I521), .ZN(W1711));
  NOR2X1 G13332 (.A1(W41497), .A2(W13520), .ZN(O18103));
  NOR2X1 G13333 (.A1(W663), .A2(I1844), .ZN(W1708));
  NOR2X1 G13334 (.A1(W13185), .A2(W2533), .ZN(W24762));
  NOR2X1 G13335 (.A1(I1593), .A2(W167), .ZN(W1706));
  NOR2X1 G13336 (.A1(W22431), .A2(W41612), .ZN(O18106));
  NOR2X1 G13337 (.A1(W16327), .A2(W229), .ZN(O18110));
  NOR2X1 G13338 (.A1(W1712), .A2(W11847), .ZN(O3581));
  NOR2X1 G13339 (.A1(W813), .A2(W718), .ZN(W1664));
  NOR2X1 G13340 (.A1(W4767), .A2(W25493), .ZN(W25937));
  NOR2X1 G13341 (.A1(I1326), .A2(W642), .ZN(W1662));
  NOR2X1 G13342 (.A1(W6516), .A2(W20609), .ZN(W24778));
  NOR2X1 G13343 (.A1(I1629), .A2(W56), .ZN(W1659));
  NOR2X1 G13344 (.A1(W12188), .A2(W11710), .ZN(W24779));
  NOR2X1 G13345 (.A1(W27232), .A2(W5506), .ZN(O18153));
  NOR2X1 G13346 (.A1(W8807), .A2(W24234), .ZN(O3582));
  NOR2X1 G13347 (.A1(W14543), .A2(W22318), .ZN(O3190));
  NOR2X1 G13348 (.A1(W989), .A2(I12), .ZN(W1652));
  NOR2X1 G13349 (.A1(W18704), .A2(W14184), .ZN(O18155));
  NOR2X1 G13350 (.A1(W44842), .A2(W3869), .ZN(O18156));
  NOR2X1 G13351 (.A1(W4853), .A2(I1036), .ZN(O3580));
  NOR2X1 G13352 (.A1(W1666), .A2(W14685), .ZN(W25925));
  NOR2X1 G13353 (.A1(I446), .A2(I866), .ZN(W1645));
  NOR2X1 G13354 (.A1(W6821), .A2(W7923), .ZN(W25920));
  NOR2X1 G13355 (.A1(I649), .A2(W1155), .ZN(W1673));
  NOR2X1 G13356 (.A1(W1477), .A2(W845), .ZN(W1681));
  NOR2X1 G13357 (.A1(W512), .A2(I1011), .ZN(W1680));
  NOR2X1 G13358 (.A1(W17707), .A2(W25676), .ZN(W25945));
  NOR2X1 G13359 (.A1(W16471), .A2(W25257), .ZN(W25942));
  NOR2X1 G13360 (.A1(W762), .A2(I176), .ZN(W1677));
  NOR2X1 G13361 (.A1(W40740), .A2(W20324), .ZN(O18134));
  NOR2X1 G13362 (.A1(I1672), .A2(I1121), .ZN(W1675));
  NOR2X1 G13363 (.A1(I1322), .A2(I467), .ZN(W1674));
  NOR2X1 G13364 (.A1(W3267), .A2(W2620), .ZN(W4451));
  NOR2X1 G13365 (.A1(W9808), .A2(W24598), .ZN(W25941));
  NOR2X1 G13366 (.A1(I746), .A2(W1421), .ZN(W1671));
  NOR2X1 G13367 (.A1(W10), .A2(W29294), .ZN(O18140));
  NOR2X1 G13368 (.A1(W13580), .A2(W4724), .ZN(W25940));
  NOR2X1 G13369 (.A1(I1648), .A2(I1777), .ZN(O18142));
  NOR2X1 G13370 (.A1(W750), .A2(W1377), .ZN(W1667));
  NOR2X1 G13371 (.A1(W2695), .A2(I274), .ZN(W25938));
  NOR2X1 G13372 (.A1(W23328), .A2(W19972), .ZN(W27846));
  NOR2X1 G13373 (.A1(W3679), .A2(W1177), .ZN(W7343));
  NOR2X1 G13374 (.A1(W489), .A2(W5917), .ZN(W7342));
  NOR2X1 G13375 (.A1(W670), .A2(W5458), .ZN(W7341));
  NOR2X1 G13376 (.A1(W4032), .A2(I1934), .ZN(W7340));
  NOR2X1 G13377 (.A1(W17414), .A2(W15866), .ZN(W22893));
  NOR2X1 G13378 (.A1(W27085), .A2(W11160), .ZN(W27848));
  NOR2X1 G13379 (.A1(W28467), .A2(W14112), .ZN(O13215));
  NOR2X1 G13380 (.A1(W14234), .A2(W37657), .ZN(O13216));
  NOR2X1 G13381 (.A1(W25919), .A2(W26087), .ZN(O4251));
  NOR2X1 G13382 (.A1(I1810), .A2(I512), .ZN(O178));
  NOR2X1 G13383 (.A1(I1478), .A2(I391), .ZN(W7333));
  NOR2X1 G13384 (.A1(W42106), .A2(W10571), .ZN(O13219));
  NOR2X1 G13385 (.A1(W3557), .A2(W2233), .ZN(O13221));
  NOR2X1 G13386 (.A1(W18125), .A2(W27129), .ZN(O4250));
  NOR2X1 G13387 (.A1(W40285), .A2(W31066), .ZN(W43568));
  NOR2X1 G13388 (.A1(W4458), .A2(W3758), .ZN(W7327));
  NOR2X1 G13389 (.A1(W2902), .A2(W5576), .ZN(W7352));
  NOR2X1 G13390 (.A1(W9811), .A2(W8523), .ZN(W22886));
  NOR2X1 G13391 (.A1(W1620), .A2(W3457), .ZN(W7363));
  NOR2X1 G13392 (.A1(I527), .A2(W71), .ZN(W7362));
  NOR2X1 G13393 (.A1(W842), .A2(W859), .ZN(W7361));
  NOR2X1 G13394 (.A1(W6118), .A2(I1681), .ZN(W7359));
  NOR2X1 G13395 (.A1(W8694), .A2(W17399), .ZN(O13202));
  NOR2X1 G13396 (.A1(W20326), .A2(W28879), .ZN(O13203));
  NOR2X1 G13397 (.A1(W8574), .A2(W20169), .ZN(O13204));
  NOR2X1 G13398 (.A1(W4414), .A2(W1369), .ZN(W7326));
  NOR2X1 G13399 (.A1(W11993), .A2(W42869), .ZN(W43547));
  NOR2X1 G13400 (.A1(W17817), .A2(W34335), .ZN(O13209));
  NOR2X1 G13401 (.A1(W2983), .A2(W2139), .ZN(W7349));
  NOR2X1 G13402 (.A1(I337), .A2(I57), .ZN(W7348));
  NOR2X1 G13403 (.A1(W39810), .A2(W718), .ZN(O13211));
  NOR2X1 G13404 (.A1(W17060), .A2(W20892), .ZN(W27850));
  NOR2X1 G13405 (.A1(W22601), .A2(W38010), .ZN(O13213));
  NOR2X1 G13406 (.A1(W14073), .A2(W11625), .ZN(O13246));
  NOR2X1 G13407 (.A1(W6298), .A2(I1076), .ZN(W7305));
  NOR2X1 G13408 (.A1(W2481), .A2(W27125), .ZN(O4244));
  NOR2X1 G13409 (.A1(W92), .A2(W3493), .ZN(W7303));
  NOR2X1 G13410 (.A1(W1534), .A2(I613), .ZN(W7302));
  NOR2X1 G13411 (.A1(W28541), .A2(W36723), .ZN(O13239));
  NOR2X1 G13412 (.A1(W249), .A2(W19314), .ZN(O13241));
  NOR2X1 G13413 (.A1(W26806), .A2(W6907), .ZN(W43593));
  NOR2X1 G13414 (.A1(W17986), .A2(W12830), .ZN(W27831));
  NOR2X1 G13415 (.A1(W4021), .A2(W1730), .ZN(W7306));
  NOR2X1 G13416 (.A1(W17173), .A2(W1040), .ZN(W43605));
  NOR2X1 G13417 (.A1(W2183), .A2(W7213), .ZN(W7293));
  NOR2X1 G13418 (.A1(W12836), .A2(W1672), .ZN(O13253));
  NOR2X1 G13419 (.A1(W14908), .A2(W20505), .ZN(O13254));
  NOR2X1 G13420 (.A1(W16173), .A2(W30613), .ZN(O13255));
  NOR2X1 G13421 (.A1(W1490), .A2(W1351), .ZN(O13256));
  NOR2X1 G13422 (.A1(W3189), .A2(W21560), .ZN(W27827));
  NOR2X1 G13423 (.A1(W2234), .A2(W6504), .ZN(W7316));
  NOR2X1 G13424 (.A1(I1806), .A2(W26375), .ZN(O13224));
  NOR2X1 G13425 (.A1(W5921), .A2(W2587), .ZN(W7324));
  NOR2X1 G13426 (.A1(W14303), .A2(W9433), .ZN(W22898));
  NOR2X1 G13427 (.A1(W39575), .A2(W3836), .ZN(O13227));
  NOR2X1 G13428 (.A1(W3286), .A2(W6120), .ZN(W7320));
  NOR2X1 G13429 (.A1(W33859), .A2(W38738), .ZN(W43575));
  NOR2X1 G13430 (.A1(W644), .A2(I1592), .ZN(W7318));
  NOR2X1 G13431 (.A1(W42699), .A2(W12646), .ZN(O13229));
  NOR2X1 G13432 (.A1(W4673), .A2(W22019), .ZN(W43536));
  NOR2X1 G13433 (.A1(W34806), .A2(W40108), .ZN(O13230));
  NOR2X1 G13434 (.A1(W6050), .A2(W2475), .ZN(W7314));
  NOR2X1 G13435 (.A1(W22005), .A2(W10638), .ZN(W43580));
  NOR2X1 G13436 (.A1(W6373), .A2(W782), .ZN(W7312));
  NOR2X1 G13437 (.A1(W2735), .A2(W8288), .ZN(O13232));
  NOR2X1 G13438 (.A1(I1712), .A2(W26177), .ZN(O4245));
  NOR2X1 G13439 (.A1(W5327), .A2(W5523), .ZN(W7307));
  NOR2X1 G13440 (.A1(W21399), .A2(W15741), .ZN(W22869));
  NOR2X1 G13441 (.A1(W25879), .A2(W20117), .ZN(W27868));
  NOR2X1 G13442 (.A1(W4663), .A2(W4951), .ZN(O13156));
  NOR2X1 G13443 (.A1(W22795), .A2(W34320), .ZN(O13157));
  NOR2X1 G13444 (.A1(W1859), .A2(W672), .ZN(W7416));
  NOR2X1 G13445 (.A1(I418), .A2(W19781), .ZN(W22867));
  NOR2X1 G13446 (.A1(W212), .A2(W7107), .ZN(W7413));
  NOR2X1 G13447 (.A1(W964), .A2(W3424), .ZN(W7411));
  NOR2X1 G13448 (.A1(W33570), .A2(W11363), .ZN(O13161));
  NOR2X1 G13449 (.A1(I1119), .A2(W4570), .ZN(W7420));
  NOR2X1 G13450 (.A1(W5294), .A2(I554), .ZN(W7408));
  NOR2X1 G13451 (.A1(W2066), .A2(W5552), .ZN(W7407));
  NOR2X1 G13452 (.A1(W3922), .A2(W20365), .ZN(W22870));
  NOR2X1 G13453 (.A1(W17752), .A2(W12573), .ZN(O13164));
  NOR2X1 G13454 (.A1(W6587), .A2(W5036), .ZN(W22871));
  NOR2X1 G13455 (.A1(W13701), .A2(W11124), .ZN(W22872));
  NOR2X1 G13456 (.A1(W6207), .A2(W5491), .ZN(W7402));
  NOR2X1 G13457 (.A1(W4719), .A2(W26954), .ZN(W27869));
  NOR2X1 G13458 (.A1(W6215), .A2(W2512), .ZN(W27872));
  NOR2X1 G13459 (.A1(W16306), .A2(W9386), .ZN(W43462));
  NOR2X1 G13460 (.A1(W5300), .A2(W2104), .ZN(W7435));
  NOR2X1 G13461 (.A1(W1386), .A2(W814), .ZN(W7434));
  NOR2X1 G13462 (.A1(W22076), .A2(W13427), .ZN(W22859));
  NOR2X1 G13463 (.A1(W6997), .A2(I1283), .ZN(W7432));
  NOR2X1 G13464 (.A1(W6997), .A2(I435), .ZN(W7431));
  NOR2X1 G13465 (.A1(W7321), .A2(I804), .ZN(W22861));
  NOR2X1 G13466 (.A1(W3610), .A2(W5837), .ZN(W7401));
  NOR2X1 G13467 (.A1(W1914), .A2(I1980), .ZN(W7427));
  NOR2X1 G13468 (.A1(W6515), .A2(W10658), .ZN(W22863));
  NOR2X1 G13469 (.A1(W14532), .A2(W12045), .ZN(O2623));
  NOR2X1 G13470 (.A1(W15124), .A2(W27355), .ZN(O13152));
  NOR2X1 G13471 (.A1(W7421), .A2(W25650), .ZN(O13153));
  NOR2X1 G13472 (.A1(W26859), .A2(W6874), .ZN(O13154));
  NOR2X1 G13473 (.A1(W2211), .A2(W2505), .ZN(W7421));
  NOR2X1 G13474 (.A1(W32514), .A2(W29444), .ZN(W43523));
  NOR2X1 G13475 (.A1(W25569), .A2(W31014), .ZN(O13180));
  NOR2X1 G13476 (.A1(I1065), .A2(W3341), .ZN(W7382));
  NOR2X1 G13477 (.A1(I887), .A2(W8237), .ZN(W22880));
  NOR2X1 G13478 (.A1(I549), .A2(W16487), .ZN(O2626));
  NOR2X1 G13479 (.A1(W7048), .A2(I258), .ZN(W7379));
  NOR2X1 G13480 (.A1(W16433), .A2(W21637), .ZN(W43513));
  NOR2X1 G13481 (.A1(W23340), .A2(W6000), .ZN(O13185));
  NOR2X1 G13482 (.A1(W37694), .A2(W528), .ZN(W43517));
  NOR2X1 G13483 (.A1(W227), .A2(W74), .ZN(O13179));
  NOR2X1 G13484 (.A1(W21752), .A2(W14271), .ZN(W27856));
  NOR2X1 G13485 (.A1(W453), .A2(W1348), .ZN(W22885));
  NOR2X1 G13486 (.A1(I626), .A2(I1308), .ZN(W7370));
  NOR2X1 G13487 (.A1(W1453), .A2(W14173), .ZN(W43532));
  NOR2X1 G13488 (.A1(W39516), .A2(W31613), .ZN(O13198));
  NOR2X1 G13489 (.A1(W39335), .A2(W11120), .ZN(W43535));
  NOR2X1 G13490 (.A1(W3167), .A2(W5752), .ZN(W7366));
  NOR2X1 G13491 (.A1(W5727), .A2(W1638), .ZN(W7287));
  NOR2X1 G13492 (.A1(W6247), .A2(W4062), .ZN(W7385));
  NOR2X1 G13493 (.A1(I313), .A2(W2892), .ZN(W22879));
  NOR2X1 G13494 (.A1(W1627), .A2(W3946), .ZN(W43504));
  NOR2X1 G13495 (.A1(I562), .A2(W11901), .ZN(W22878));
  NOR2X1 G13496 (.A1(W27036), .A2(W26030), .ZN(W27861));
  NOR2X1 G13497 (.A1(W4246), .A2(W17860), .ZN(W22875));
  NOR2X1 G13498 (.A1(I1168), .A2(W5687), .ZN(W7392));
  NOR2X1 G13499 (.A1(I965), .A2(I1030), .ZN(W7393));
  NOR2X1 G13500 (.A1(W6793), .A2(W4749), .ZN(W7394));
  NOR2X1 G13501 (.A1(W31622), .A2(I1622), .ZN(O13172));
  NOR2X1 G13502 (.A1(I1268), .A2(W29122), .ZN(O13170));
  NOR2X1 G13503 (.A1(W2738), .A2(W266), .ZN(W7397));
  NOR2X1 G13504 (.A1(W3686), .A2(W4391), .ZN(O4257));
  NOR2X1 G13505 (.A1(W24643), .A2(W23688), .ZN(O4258));
  NOR2X1 G13506 (.A1(I1366), .A2(W4179), .ZN(W7400));
  NOR2X1 G13507 (.A1(W912), .A2(W2621), .ZN(W7185));
  NOR2X1 G13508 (.A1(W23911), .A2(W19751), .ZN(O13314));
  NOR2X1 G13509 (.A1(W8176), .A2(W13600), .ZN(O13315));
  NOR2X1 G13510 (.A1(I1639), .A2(W1311), .ZN(W7192));
  NOR2X1 G13511 (.A1(W10052), .A2(W19582), .ZN(O13316));
  NOR2X1 G13512 (.A1(W5957), .A2(W817), .ZN(W7189));
  NOR2X1 G13513 (.A1(I1467), .A2(W16602), .ZN(O13318));
  NOR2X1 G13514 (.A1(W25581), .A2(W25599), .ZN(O13319));
  NOR2X1 G13515 (.A1(W8201), .A2(W8027), .ZN(O13323));
  NOR2X1 G13516 (.A1(W1197), .A2(W3640), .ZN(W27803));
  NOR2X1 G13517 (.A1(W16158), .A2(W9252), .ZN(W27800));
  NOR2X1 G13518 (.A1(W21298), .A2(W24251), .ZN(W27799));
  NOR2X1 G13519 (.A1(W5887), .A2(W20489), .ZN(O13325));
  NOR2X1 G13520 (.A1(W898), .A2(I1837), .ZN(O168));
  NOR2X1 G13521 (.A1(W37041), .A2(W37017), .ZN(O13326));
  NOR2X1 G13522 (.A1(I1875), .A2(W14881), .ZN(O13327));
  NOR2X1 G13523 (.A1(I1608), .A2(W14830), .ZN(W22937));
  NOR2X1 G13524 (.A1(W25959), .A2(W20135), .ZN(O4238));
  NOR2X1 G13525 (.A1(W32423), .A2(W21776), .ZN(W43679));
  NOR2X1 G13526 (.A1(I75), .A2(W5593), .ZN(W7212));
  NOR2X1 G13527 (.A1(W2545), .A2(W12723), .ZN(W43682));
  NOR2X1 G13528 (.A1(W22229), .A2(W38595), .ZN(W43683));
  NOR2X1 G13529 (.A1(W8090), .A2(W1394), .ZN(W22928));
  NOR2X1 G13530 (.A1(W1162), .A2(W2219), .ZN(W7207));
  NOR2X1 G13531 (.A1(W4240), .A2(W18098), .ZN(O2639));
  NOR2X1 G13532 (.A1(W4205), .A2(W1671), .ZN(W7205));
  NOR2X1 G13533 (.A1(I1004), .A2(W19855), .ZN(W22938));
  NOR2X1 G13534 (.A1(W10436), .A2(W383), .ZN(O4237));
  NOR2X1 G13535 (.A1(W788), .A2(W36015), .ZN(W43691));
  NOR2X1 G13536 (.A1(W609), .A2(W4800), .ZN(W7201));
  NOR2X1 G13537 (.A1(W15778), .A2(W26621), .ZN(W43692));
  NOR2X1 G13538 (.A1(W35848), .A2(W10746), .ZN(W43694));
  NOR2X1 G13539 (.A1(W43205), .A2(W4750), .ZN(W43695));
  NOR2X1 G13540 (.A1(W6654), .A2(W522), .ZN(W7197));
  NOR2X1 G13541 (.A1(W11802), .A2(W21775), .ZN(W22951));
  NOR2X1 G13542 (.A1(W13768), .A2(W398), .ZN(W22947));
  NOR2X1 G13543 (.A1(W6379), .A2(W2241), .ZN(W7157));
  NOR2X1 G13544 (.A1(W26725), .A2(W19330), .ZN(O4234));
  NOR2X1 G13545 (.A1(W36501), .A2(W29790), .ZN(O13351));
  NOR2X1 G13546 (.A1(W29209), .A2(W41926), .ZN(O13352));
  NOR2X1 G13547 (.A1(W7043), .A2(W4492), .ZN(W7153));
  NOR2X1 G13548 (.A1(W12897), .A2(W8166), .ZN(O4233));
  NOR2X1 G13549 (.A1(W2185), .A2(W6921), .ZN(O167));
  NOR2X1 G13550 (.A1(W2616), .A2(W2626), .ZN(W27792));
  NOR2X1 G13551 (.A1(I1608), .A2(W136), .ZN(W7147));
  NOR2X1 G13552 (.A1(W2391), .A2(W4113), .ZN(W7146));
  NOR2X1 G13553 (.A1(W8752), .A2(W22602), .ZN(O13357));
  NOR2X1 G13554 (.A1(W13775), .A2(W7135), .ZN(O13359));
  NOR2X1 G13555 (.A1(I1617), .A2(W4275), .ZN(W7141));
  NOR2X1 G13556 (.A1(W823), .A2(W4332), .ZN(W7140));
  NOR2X1 G13557 (.A1(W25334), .A2(W12991), .ZN(O13360));
  NOR2X1 G13558 (.A1(W11169), .A2(I146), .ZN(W27795));
  NOR2X1 G13559 (.A1(W17053), .A2(W9499), .ZN(W22939));
  NOR2X1 G13560 (.A1(W35225), .A2(W26575), .ZN(O13333));
  NOR2X1 G13561 (.A1(W30769), .A2(W36798), .ZN(O13334));
  NOR2X1 G13562 (.A1(W43129), .A2(W20947), .ZN(O13335));
  NOR2X1 G13563 (.A1(W22779), .A2(W10895), .ZN(O13337));
  NOR2X1 G13564 (.A1(W3742), .A2(W7040), .ZN(W7171));
  NOR2X1 G13565 (.A1(W20077), .A2(W2633), .ZN(W22940));
  NOR2X1 G13566 (.A1(W2475), .A2(W10532), .ZN(W22941));
  NOR2X1 G13567 (.A1(W12288), .A2(W24500), .ZN(W43678));
  NOR2X1 G13568 (.A1(W4317), .A2(W377), .ZN(W7166));
  NOR2X1 G13569 (.A1(W20436), .A2(W13452), .ZN(O4235));
  NOR2X1 G13570 (.A1(W9796), .A2(W1813), .ZN(O13344));
  NOR2X1 G13571 (.A1(W2600), .A2(W219), .ZN(W22945));
  NOR2X1 G13572 (.A1(W4979), .A2(I1538), .ZN(W7162));
  NOR2X1 G13573 (.A1(W4493), .A2(W5613), .ZN(W7161));
  NOR2X1 G13574 (.A1(W4275), .A2(W1847), .ZN(W7160));
  NOR2X1 G13575 (.A1(W12465), .A2(W4196), .ZN(W22915));
  NOR2X1 G13576 (.A1(W6794), .A2(W6461), .ZN(O174));
  NOR2X1 G13577 (.A1(W3194), .A2(W9557), .ZN(W22912));
  NOR2X1 G13578 (.A1(W6224), .A2(W2764), .ZN(W7266));
  NOR2X1 G13579 (.A1(W13816), .A2(W27664), .ZN(O13274));
  NOR2X1 G13580 (.A1(W5962), .A2(W5641), .ZN(W7264));
  NOR2X1 G13581 (.A1(W15774), .A2(W15322), .ZN(O4242));
  NOR2X1 G13582 (.A1(I1712), .A2(I446), .ZN(W7262));
  NOR2X1 G13583 (.A1(W2280), .A2(W75), .ZN(W7261));
  NOR2X1 G13584 (.A1(W826), .A2(W943), .ZN(W7270));
  NOR2X1 G13585 (.A1(W833), .A2(I297), .ZN(W7259));
  NOR2X1 G13586 (.A1(W25076), .A2(W40400), .ZN(O13276));
  NOR2X1 G13587 (.A1(W2850), .A2(W284), .ZN(W7257));
  NOR2X1 G13588 (.A1(W1125), .A2(W3633), .ZN(W7256));
  NOR2X1 G13589 (.A1(I1439), .A2(W6158), .ZN(W7255));
  NOR2X1 G13590 (.A1(W6411), .A2(I1698), .ZN(W7254));
  NOR2X1 G13591 (.A1(W2056), .A2(W5034), .ZN(W7253));
  NOR2X1 G13592 (.A1(W27778), .A2(W2815), .ZN(O13265));
  NOR2X1 G13593 (.A1(W27), .A2(W2284), .ZN(W7286));
  NOR2X1 G13594 (.A1(I710), .A2(W2937), .ZN(W7285));
  NOR2X1 G13595 (.A1(W20976), .A2(W10112), .ZN(W22908));
  NOR2X1 G13596 (.A1(W36503), .A2(W12062), .ZN(O13260));
  NOR2X1 G13597 (.A1(W21544), .A2(W29954), .ZN(O13262));
  NOR2X1 G13598 (.A1(W19099), .A2(W14520), .ZN(W22909));
  NOR2X1 G13599 (.A1(W4587), .A2(W401), .ZN(O13263));
  NOR2X1 G13600 (.A1(W5419), .A2(W20992), .ZN(O13264));
  NOR2X1 G13601 (.A1(W42164), .A2(W31963), .ZN(O13278));
  NOR2X1 G13602 (.A1(W4673), .A2(W5340), .ZN(W7277));
  NOR2X1 G13603 (.A1(W1839), .A2(W2229), .ZN(W7276));
  NOR2X1 G13604 (.A1(W19479), .A2(W7375), .ZN(W43622));
  NOR2X1 G13605 (.A1(W17455), .A2(W24053), .ZN(W27826));
  NOR2X1 G13606 (.A1(W12042), .A2(W27953), .ZN(O13267));
  NOR2X1 G13607 (.A1(W3148), .A2(W17630), .ZN(W27824));
  NOR2X1 G13608 (.A1(W14838), .A2(W3937), .ZN(O13272));
  NOR2X1 G13609 (.A1(W31649), .A2(W1104), .ZN(W43668));
  NOR2X1 G13610 (.A1(W9502), .A2(W4937), .ZN(W27812));
  NOR2X1 G13611 (.A1(W14786), .A2(W38609), .ZN(O13292));
  NOR2X1 G13612 (.A1(W7361), .A2(W12313), .ZN(W22925));
  NOR2X1 G13613 (.A1(W4052), .A2(W4478), .ZN(W7227));
  NOR2X1 G13614 (.A1(W260), .A2(W3883), .ZN(W7226));
  NOR2X1 G13615 (.A1(W16521), .A2(W27054), .ZN(W27811));
  NOR2X1 G13616 (.A1(W2693), .A2(W10325), .ZN(O13296));
  NOR2X1 G13617 (.A1(W4108), .A2(I1769), .ZN(W7223));
  NOR2X1 G13618 (.A1(W22937), .A2(W22397), .ZN(O4240));
  NOR2X1 G13619 (.A1(W34377), .A2(W14143), .ZN(W43669));
  NOR2X1 G13620 (.A1(W19964), .A2(W9570), .ZN(O13297));
  NOR2X1 G13621 (.A1(W27003), .A2(W11990), .ZN(W43672));
  NOR2X1 G13622 (.A1(I1732), .A2(W2874), .ZN(O171));
  NOR2X1 G13623 (.A1(W1374), .A2(W6119), .ZN(W7217));
  NOR2X1 G13624 (.A1(W4348), .A2(W11774), .ZN(O13302));
  NOR2X1 G13625 (.A1(W3828), .A2(W2742), .ZN(W7215));
  NOR2X1 G13626 (.A1(W20720), .A2(I995), .ZN(W43460));
  NOR2X1 G13627 (.A1(W797), .A2(W2185), .ZN(W7232));
  NOR2X1 G13628 (.A1(W6935), .A2(W3658), .ZN(O13289));
  NOR2X1 G13629 (.A1(W4707), .A2(W1224), .ZN(W7234));
  NOR2X1 G13630 (.A1(W5184), .A2(W5460), .ZN(W7236));
  NOR2X1 G13631 (.A1(W6264), .A2(W11955), .ZN(W43658));
  NOR2X1 G13632 (.A1(W39225), .A2(W2718), .ZN(W43657));
  NOR2X1 G13633 (.A1(W4156), .A2(W2755), .ZN(W7239));
  NOR2X1 G13634 (.A1(W1097), .A2(W4137), .ZN(W43654));
  NOR2X1 G13635 (.A1(W12608), .A2(W13489), .ZN(W27815));
  NOR2X1 G13636 (.A1(W38298), .A2(W30564), .ZN(O13284));
  NOR2X1 G13637 (.A1(W4996), .A2(W4822), .ZN(W7244));
  NOR2X1 G13638 (.A1(W40178), .A2(W41808), .ZN(W43646));
  NOR2X1 G13639 (.A1(W12917), .A2(W22540), .ZN(O2637));
  NOR2X1 G13640 (.A1(W3702), .A2(W37274), .ZN(O13279));
  NOR2X1 G13641 (.A1(W5277), .A2(W6381), .ZN(W7250));
  NOR2X1 G13642 (.A1(I1679), .A2(W2923), .ZN(W7638));
  NOR2X1 G13643 (.A1(W7645), .A2(W14747), .ZN(O12969));
  NOR2X1 G13644 (.A1(W4346), .A2(W1182), .ZN(W7645));
  NOR2X1 G13645 (.A1(W22295), .A2(I147), .ZN(O2614));
  NOR2X1 G13646 (.A1(W20779), .A2(W25621), .ZN(O4294));
  NOR2X1 G13647 (.A1(W14950), .A2(W21742), .ZN(W22784));
  NOR2X1 G13648 (.A1(W1521), .A2(W24805), .ZN(O12973));
  NOR2X1 G13649 (.A1(W5682), .A2(W7564), .ZN(W7640));
  NOR2X1 G13650 (.A1(I179), .A2(W5748), .ZN(W7639));
  NOR2X1 G13651 (.A1(W6649), .A2(W41006), .ZN(O12968));
  NOR2X1 G13652 (.A1(W13285), .A2(I326), .ZN(W22785));
  NOR2X1 G13653 (.A1(W1460), .A2(W41920), .ZN(O12975));
  NOR2X1 G13654 (.A1(W7003), .A2(W231), .ZN(W7635));
  NOR2X1 G13655 (.A1(W5029), .A2(W111), .ZN(W7634));
  NOR2X1 G13656 (.A1(W7014), .A2(W4802), .ZN(W7633));
  NOR2X1 G13657 (.A1(W17762), .A2(I346), .ZN(O12976));
  NOR2X1 G13658 (.A1(W38223), .A2(W35907), .ZN(O12977));
  NOR2X1 G13659 (.A1(W6600), .A2(I86), .ZN(O12959));
  NOR2X1 G13660 (.A1(W15644), .A2(W18600), .ZN(W27967));
  NOR2X1 G13661 (.A1(W5232), .A2(W2570), .ZN(W7665));
  NOR2X1 G13662 (.A1(W947), .A2(W5042), .ZN(W7663));
  NOR2X1 G13663 (.A1(W5691), .A2(W6447), .ZN(W7662));
  NOR2X1 G13664 (.A1(I1373), .A2(W1959), .ZN(W7661));
  NOR2X1 G13665 (.A1(W14448), .A2(W10341), .ZN(O12956));
  NOR2X1 G13666 (.A1(W16308), .A2(W6226), .ZN(W22777));
  NOR2X1 G13667 (.A1(W2636), .A2(W28252), .ZN(O12958));
  NOR2X1 G13668 (.A1(W955), .A2(W27173), .ZN(W43262));
  NOR2X1 G13669 (.A1(W25471), .A2(W17811), .ZN(W27962));
  NOR2X1 G13670 (.A1(W628), .A2(I362), .ZN(O4295));
  NOR2X1 G13671 (.A1(W3526), .A2(I752), .ZN(W7652));
  NOR2X1 G13672 (.A1(W13881), .A2(W8413), .ZN(W43244));
  NOR2X1 G13673 (.A1(W38587), .A2(W14036), .ZN(O12965));
  NOR2X1 G13674 (.A1(W15140), .A2(I572), .ZN(W27959));
  NOR2X1 G13675 (.A1(W1284), .A2(W4990), .ZN(W7648));
  NOR2X1 G13676 (.A1(W18908), .A2(W35311), .ZN(W43305));
  NOR2X1 G13677 (.A1(W235), .A2(W13680), .ZN(O13009));
  NOR2X1 G13678 (.A1(W15511), .A2(I780), .ZN(O13011));
  NOR2X1 G13679 (.A1(W10792), .A2(W19763), .ZN(W27938));
  NOR2X1 G13680 (.A1(W16085), .A2(W42345), .ZN(O13015));
  NOR2X1 G13681 (.A1(I608), .A2(W12853), .ZN(W43301));
  NOR2X1 G13682 (.A1(W30103), .A2(W9936), .ZN(O13016));
  NOR2X1 G13683 (.A1(W5451), .A2(W6956), .ZN(W7598));
  NOR2X1 G13684 (.A1(W11696), .A2(W34999), .ZN(O13018));
  NOR2X1 G13685 (.A1(W1465), .A2(W138), .ZN(W7606));
  NOR2X1 G13686 (.A1(W5492), .A2(I1809), .ZN(W7595));
  NOR2X1 G13687 (.A1(I1909), .A2(W5652), .ZN(W7594));
  NOR2X1 G13688 (.A1(W16049), .A2(W6399), .ZN(W22802));
  NOR2X1 G13689 (.A1(W15036), .A2(W784), .ZN(O13022));
  NOR2X1 G13690 (.A1(W6768), .A2(W267), .ZN(W7591));
  NOR2X1 G13691 (.A1(W6561), .A2(W16341), .ZN(O13024));
  NOR2X1 G13692 (.A1(W7004), .A2(I65), .ZN(W7589));
  NOR2X1 G13693 (.A1(W7076), .A2(I879), .ZN(W7619));
  NOR2X1 G13694 (.A1(W17417), .A2(W8658), .ZN(O2615));
  NOR2X1 G13695 (.A1(W1682), .A2(W12623), .ZN(W27956));
  NOR2X1 G13696 (.A1(W17633), .A2(W25263), .ZN(W27954));
  NOR2X1 G13697 (.A1(W16158), .A2(W2918), .ZN(W27953));
  NOR2X1 G13698 (.A1(W12902), .A2(W10664), .ZN(O12991));
  NOR2X1 G13699 (.A1(W35012), .A2(W20584), .ZN(O12992));
  NOR2X1 G13700 (.A1(W1823), .A2(W568), .ZN(W7621));
  NOR2X1 G13701 (.A1(W3917), .A2(W2614), .ZN(W7620));
  NOR2X1 G13702 (.A1(W19462), .A2(W8212), .ZN(O12954));
  NOR2X1 G13703 (.A1(W25678), .A2(I898), .ZN(O12999));
  NOR2X1 G13704 (.A1(W593), .A2(W11938), .ZN(W27944));
  NOR2X1 G13705 (.A1(W5672), .A2(W26636), .ZN(W27942));
  NOR2X1 G13706 (.A1(W5565), .A2(W4471), .ZN(W7611));
  NOR2X1 G13707 (.A1(W42860), .A2(W4320), .ZN(O13003));
  NOR2X1 G13708 (.A1(W1930), .A2(W10286), .ZN(O4290));
  NOR2X1 G13709 (.A1(W656), .A2(W5815), .ZN(W7608));
  NOR2X1 G13710 (.A1(W17061), .A2(W12689), .ZN(W22757));
  NOR2X1 G13711 (.A1(W8631), .A2(W9990), .ZN(W27996));
  NOR2X1 G13712 (.A1(W12540), .A2(W3074), .ZN(W22753));
  NOR2X1 G13713 (.A1(W7264), .A2(W6745), .ZN(W7720));
  NOR2X1 G13714 (.A1(W17182), .A2(W17015), .ZN(O4308));
  NOR2X1 G13715 (.A1(W10681), .A2(W609), .ZN(W27994));
  NOR2X1 G13716 (.A1(W40787), .A2(W15757), .ZN(O12906));
  NOR2X1 G13717 (.A1(W12385), .A2(W17540), .ZN(W27992));
  NOR2X1 G13718 (.A1(W15406), .A2(W18105), .ZN(W43173));
  NOR2X1 G13719 (.A1(W20405), .A2(W36880), .ZN(O12900));
  NOR2X1 G13720 (.A1(W1950), .A2(W33491), .ZN(O12914));
  NOR2X1 G13721 (.A1(W5234), .A2(W13529), .ZN(W27987));
  NOR2X1 G13722 (.A1(W4859), .A2(W4698), .ZN(W7710));
  NOR2X1 G13723 (.A1(W1025), .A2(W2343), .ZN(W7708));
  NOR2X1 G13724 (.A1(W8031), .A2(W2584), .ZN(W27983));
  NOR2X1 G13725 (.A1(W42305), .A2(W21047), .ZN(O12918));
  NOR2X1 G13726 (.A1(W26713), .A2(W23949), .ZN(W27982));
  NOR2X1 G13727 (.A1(I306), .A2(W1111), .ZN(W7731));
  NOR2X1 G13728 (.A1(W721), .A2(W2974), .ZN(W7740));
  NOR2X1 G13729 (.A1(W15151), .A2(W27108), .ZN(W43147));
  NOR2X1 G13730 (.A1(W16856), .A2(W12728), .ZN(W22748));
  NOR2X1 G13731 (.A1(W24940), .A2(W2523), .ZN(W43153));
  NOR2X1 G13732 (.A1(W2475), .A2(W6321), .ZN(W7736));
  NOR2X1 G13733 (.A1(W8497), .A2(W12498), .ZN(W43155));
  NOR2X1 G13734 (.A1(W21780), .A2(W12137), .ZN(O12891));
  NOR2X1 G13735 (.A1(W25826), .A2(W27105), .ZN(O12892));
  NOR2X1 G13736 (.A1(W38702), .A2(W12550), .ZN(O12921));
  NOR2X1 G13737 (.A1(W1488), .A2(W27764), .ZN(O12894));
  NOR2X1 G13738 (.A1(W9474), .A2(W1301), .ZN(W27998));
  NOR2X1 G13739 (.A1(W1973), .A2(W6946), .ZN(W7728));
  NOR2X1 G13740 (.A1(W26699), .A2(W31322), .ZN(O12896));
  NOR2X1 G13741 (.A1(W19532), .A2(W23812), .ZN(W27997));
  NOR2X1 G13742 (.A1(W25248), .A2(W23179), .ZN(O12899));
  NOR2X1 G13743 (.A1(I928), .A2(W4091), .ZN(W7724));
  NOR2X1 G13744 (.A1(W26607), .A2(W22772), .ZN(W43223));
  NOR2X1 G13745 (.A1(W6406), .A2(W125), .ZN(W7686));
  NOR2X1 G13746 (.A1(W16446), .A2(W12132), .ZN(O4302));
  NOR2X1 G13747 (.A1(W18300), .A2(W1320), .ZN(O4300));
  NOR2X1 G13748 (.A1(W7119), .A2(I1490), .ZN(O194));
  NOR2X1 G13749 (.A1(W508), .A2(W5309), .ZN(W7682));
  NOR2X1 G13750 (.A1(W38879), .A2(W13140), .ZN(O12946));
  NOR2X1 G13751 (.A1(W5153), .A2(I968), .ZN(W7679));
  NOR2X1 G13752 (.A1(W1075), .A2(W4992), .ZN(W7678));
  NOR2X1 G13753 (.A1(W7090), .A2(W7072), .ZN(O4303));
  NOR2X1 G13754 (.A1(I313), .A2(W7119), .ZN(W7675));
  NOR2X1 G13755 (.A1(W28551), .A2(W9432), .ZN(W43224));
  NOR2X1 G13756 (.A1(W8429), .A2(W35630), .ZN(O12948));
  NOR2X1 G13757 (.A1(W6062), .A2(W6818), .ZN(W7671));
  NOR2X1 G13758 (.A1(W34149), .A2(W41189), .ZN(O12951));
  NOR2X1 G13759 (.A1(W22550), .A2(I146), .ZN(O12952));
  NOR2X1 G13760 (.A1(W40848), .A2(W39354), .ZN(O12953));
  NOR2X1 G13761 (.A1(W4703), .A2(W5426), .ZN(W7588));
  NOR2X1 G13762 (.A1(W12721), .A2(W20865), .ZN(O12939));
  NOR2X1 G13763 (.A1(W2599), .A2(W7368), .ZN(W7689));
  NOR2X1 G13764 (.A1(W14890), .A2(W22878), .ZN(W27977));
  NOR2X1 G13765 (.A1(W5379), .A2(W14314), .ZN(O2606));
  NOR2X1 G13766 (.A1(W38354), .A2(W7302), .ZN(O12934));
  NOR2X1 G13767 (.A1(W115), .A2(W17221), .ZN(W22764));
  NOR2X1 G13768 (.A1(W6308), .A2(W7082), .ZN(W7695));
  NOR2X1 G13769 (.A1(W42898), .A2(W32921), .ZN(W43203));
  NOR2X1 G13770 (.A1(W6849), .A2(W9676), .ZN(O4305));
  NOR2X1 G13771 (.A1(W18961), .A2(W27367), .ZN(O12929));
  NOR2X1 G13772 (.A1(I1243), .A2(W29553), .ZN(O12926));
  NOR2X1 G13773 (.A1(W5593), .A2(W679), .ZN(W7700));
  NOR2X1 G13774 (.A1(W26179), .A2(W41775), .ZN(O12925));
  NOR2X1 G13775 (.A1(W7521), .A2(I1795), .ZN(W7702));
  NOR2X1 G13776 (.A1(W38922), .A2(W26001), .ZN(O12923));
  NOR2X1 G13777 (.A1(W981), .A2(I1959), .ZN(W7482));
  NOR2X1 G13778 (.A1(I920), .A2(W6892), .ZN(W7490));
  NOR2X1 G13779 (.A1(W191), .A2(W917), .ZN(W7489));
  NOR2X1 G13780 (.A1(W17980), .A2(W12281), .ZN(O13105));
  NOR2X1 G13781 (.A1(W14403), .A2(W33400), .ZN(O13106));
  NOR2X1 G13782 (.A1(W6361), .A2(W872), .ZN(W7486));
  NOR2X1 G13783 (.A1(W22539), .A2(W13755), .ZN(W27891));
  NOR2X1 G13784 (.A1(W7444), .A2(W2048), .ZN(O186));
  NOR2X1 G13785 (.A1(W5287), .A2(W20691), .ZN(W22846));
  NOR2X1 G13786 (.A1(W33890), .A2(W10608), .ZN(W43411));
  NOR2X1 G13787 (.A1(W841), .A2(W6871), .ZN(W7481));
  NOR2X1 G13788 (.A1(W42552), .A2(W22007), .ZN(O13108));
  NOR2X1 G13789 (.A1(W4559), .A2(I815), .ZN(W7479));
  NOR2X1 G13790 (.A1(W4622), .A2(W2001), .ZN(W7478));
  NOR2X1 G13791 (.A1(I1212), .A2(W7233), .ZN(W7477));
  NOR2X1 G13792 (.A1(W26748), .A2(W9401), .ZN(O13110));
  NOR2X1 G13793 (.A1(W32674), .A2(W20110), .ZN(W43420));
  NOR2X1 G13794 (.A1(W27504), .A2(W20538), .ZN(O13097));
  NOR2X1 G13795 (.A1(W5342), .A2(W19396), .ZN(O4268));
  NOR2X1 G13796 (.A1(W3716), .A2(W407), .ZN(W7508));
  NOR2X1 G13797 (.A1(W4239), .A2(W3274), .ZN(W7506));
  NOR2X1 G13798 (.A1(W3304), .A2(W3330), .ZN(W7505));
  NOR2X1 G13799 (.A1(W36736), .A2(W5001), .ZN(W43395));
  NOR2X1 G13800 (.A1(I1031), .A2(W1867), .ZN(W7502));
  NOR2X1 G13801 (.A1(W1986), .A2(W3527), .ZN(W22842));
  NOR2X1 G13802 (.A1(W4303), .A2(W847), .ZN(W27893));
  NOR2X1 G13803 (.A1(W21758), .A2(W12467), .ZN(O2621));
  NOR2X1 G13804 (.A1(W5992), .A2(W2027), .ZN(W7498));
  NOR2X1 G13805 (.A1(W29582), .A2(W13433), .ZN(W43402));
  NOR2X1 G13806 (.A1(W4755), .A2(W23779), .ZN(W27892));
  NOR2X1 G13807 (.A1(W34117), .A2(W43054), .ZN(O13099));
  NOR2X1 G13808 (.A1(W1914), .A2(W300), .ZN(W7494));
  NOR2X1 G13809 (.A1(W34248), .A2(W40412), .ZN(O13104));
  NOR2X1 G13810 (.A1(W487), .A2(W7107), .ZN(W7492));
  NOR2X1 G13811 (.A1(W1123), .A2(W9793), .ZN(W22857));
  NOR2X1 G13812 (.A1(W19866), .A2(I1937), .ZN(W43437));
  NOR2X1 G13813 (.A1(W13765), .A2(W4127), .ZN(O13124));
  NOR2X1 G13814 (.A1(W4842), .A2(I930), .ZN(W7454));
  NOR2X1 G13815 (.A1(W11831), .A2(W7806), .ZN(W27880));
  NOR2X1 G13816 (.A1(W34872), .A2(W9989), .ZN(W43440));
  NOR2X1 G13817 (.A1(W15416), .A2(W7878), .ZN(O13128));
  NOR2X1 G13818 (.A1(W4436), .A2(W27897), .ZN(O13131));
  NOR2X1 G13819 (.A1(W37510), .A2(I1459), .ZN(O13132));
  NOR2X1 G13820 (.A1(W2829), .A2(W5268), .ZN(O184));
  NOR2X1 G13821 (.A1(W35881), .A2(W40082), .ZN(O13136));
  NOR2X1 G13822 (.A1(W8176), .A2(W5869), .ZN(O13137));
  NOR2X1 G13823 (.A1(W1720), .A2(W3204), .ZN(W7443));
  NOR2X1 G13824 (.A1(W4147), .A2(W1528), .ZN(W7442));
  NOR2X1 G13825 (.A1(W39681), .A2(W38805), .ZN(O13139));
  NOR2X1 G13826 (.A1(W4250), .A2(W6985), .ZN(W7440));
  NOR2X1 G13827 (.A1(W39184), .A2(W37810), .ZN(W43459));
  NOR2X1 G13828 (.A1(W12356), .A2(W38669), .ZN(O13089));
  NOR2X1 G13829 (.A1(W2331), .A2(I1288), .ZN(W7458));
  NOR2X1 G13830 (.A1(W7958), .A2(W12320), .ZN(W22853));
  NOR2X1 G13831 (.A1(I192), .A2(W340), .ZN(O185));
  NOR2X1 G13832 (.A1(W4690), .A2(W706), .ZN(W7461));
  NOR2X1 G13833 (.A1(W21689), .A2(W42478), .ZN(O13121));
  NOR2X1 G13834 (.A1(W15842), .A2(W3516), .ZN(W27885));
  NOR2X1 G13835 (.A1(W7121), .A2(I1333), .ZN(W7465));
  NOR2X1 G13836 (.A1(W1697), .A2(W8138), .ZN(W22850));
  NOR2X1 G13837 (.A1(W27544), .A2(W36529), .ZN(O13117));
  NOR2X1 G13838 (.A1(W26686), .A2(W4491), .ZN(O13116));
  NOR2X1 G13839 (.A1(W30414), .A2(W18795), .ZN(O13115));
  NOR2X1 G13840 (.A1(W16956), .A2(W33055), .ZN(O13114));
  NOR2X1 G13841 (.A1(W18354), .A2(W5015), .ZN(W27889));
  NOR2X1 G13842 (.A1(W17342), .A2(W27421), .ZN(W43423));
  NOR2X1 G13843 (.A1(W1694), .A2(W23358), .ZN(W27890));
  NOR2X1 G13844 (.A1(W2150), .A2(I1246), .ZN(W7559));
  NOR2X1 G13845 (.A1(I1466), .A2(W17607), .ZN(O13037));
  NOR2X1 G13846 (.A1(W17271), .A2(I802), .ZN(W22807));
  NOR2X1 G13847 (.A1(W6327), .A2(W14757), .ZN(O4285));
  NOR2X1 G13848 (.A1(W8551), .A2(W22384), .ZN(W22809));
  NOR2X1 G13849 (.A1(W11789), .A2(W25951), .ZN(O13042));
  NOR2X1 G13850 (.A1(W826), .A2(W2630), .ZN(W7563));
  NOR2X1 G13851 (.A1(W19477), .A2(W27200), .ZN(O4283));
  NOR2X1 G13852 (.A1(W1313), .A2(W3305), .ZN(O189));
  NOR2X1 G13853 (.A1(I204), .A2(W4974), .ZN(W7570));
  NOR2X1 G13854 (.A1(W1893), .A2(W2719), .ZN(W7557));
  NOR2X1 G13855 (.A1(W2953), .A2(W10739), .ZN(O13049));
  NOR2X1 G13856 (.A1(W26843), .A2(W22242), .ZN(W27927));
  NOR2X1 G13857 (.A1(W26675), .A2(W5493), .ZN(O4281));
  NOR2X1 G13858 (.A1(W14607), .A2(W6958), .ZN(W22817));
  NOR2X1 G13859 (.A1(W17098), .A2(I1065), .ZN(W27924));
  NOR2X1 G13860 (.A1(W4222), .A2(W7289), .ZN(W7550));
  NOR2X1 G13861 (.A1(W3720), .A2(I521), .ZN(W7578));
  NOR2X1 G13862 (.A1(W388), .A2(W1354), .ZN(O13025));
  NOR2X1 G13863 (.A1(W4215), .A2(W31520), .ZN(O13026));
  NOR2X1 G13864 (.A1(W775), .A2(W103), .ZN(W7584));
  NOR2X1 G13865 (.A1(W3909), .A2(W6378), .ZN(W7583));
  NOR2X1 G13866 (.A1(W14022), .A2(W4342), .ZN(O13029));
  NOR2X1 G13867 (.A1(I1166), .A2(W33691), .ZN(O13030));
  NOR2X1 G13868 (.A1(W1453), .A2(I698), .ZN(W7580));
  NOR2X1 G13869 (.A1(W6731), .A2(W320), .ZN(O2617));
  NOR2X1 G13870 (.A1(W18819), .A2(W23852), .ZN(O13055));
  NOR2X1 G13871 (.A1(W18804), .A2(I1421), .ZN(W22805));
  NOR2X1 G13872 (.A1(W4655), .A2(W3162), .ZN(W7576));
  NOR2X1 G13873 (.A1(I1138), .A2(W2135), .ZN(W7575));
  NOR2X1 G13874 (.A1(W9679), .A2(W12415), .ZN(O13033));
  NOR2X1 G13875 (.A1(W36216), .A2(W12910), .ZN(O13034));
  NOR2X1 G13876 (.A1(W6376), .A2(W5893), .ZN(W7572));
  NOR2X1 G13877 (.A1(W12019), .A2(W22495), .ZN(W22806));
  NOR2X1 G13878 (.A1(W4077), .A2(W3694), .ZN(W7519));
  NOR2X1 G13879 (.A1(W1339), .A2(W1735), .ZN(W7529));
  NOR2X1 G13880 (.A1(W10619), .A2(W10889), .ZN(W27911));
  NOR2X1 G13881 (.A1(I1176), .A2(W1312), .ZN(W22831));
  NOR2X1 G13882 (.A1(W16122), .A2(W821), .ZN(W22832));
  NOR2X1 G13883 (.A1(W23533), .A2(W17981), .ZN(W27908));
  NOR2X1 G13884 (.A1(W16366), .A2(W5705), .ZN(W27905));
  NOR2X1 G13885 (.A1(W962), .A2(W5360), .ZN(W7521));
  NOR2X1 G13886 (.A1(W27339), .A2(W32351), .ZN(O13083));
  NOR2X1 G13887 (.A1(W14659), .A2(W5386), .ZN(O4276));
  NOR2X1 G13888 (.A1(W14486), .A2(W3422), .ZN(O4272));
  NOR2X1 G13889 (.A1(I625), .A2(I1338), .ZN(O187));
  NOR2X1 G13890 (.A1(W36631), .A2(W18726), .ZN(O13087));
  NOR2X1 G13891 (.A1(W4597), .A2(W6726), .ZN(W7515));
  NOR2X1 G13892 (.A1(I941), .A2(W6079), .ZN(W7514));
  NOR2X1 G13893 (.A1(W26994), .A2(W40688), .ZN(W43387));
  NOR2X1 G13894 (.A1(W22596), .A2(W29321), .ZN(O13088));
  NOR2X1 G13895 (.A1(W16087), .A2(W28526), .ZN(O13361));
  NOR2X1 G13896 (.A1(W6008), .A2(W5217), .ZN(W7531));
  NOR2X1 G13897 (.A1(W10610), .A2(W6166), .ZN(W27915));
  NOR2X1 G13898 (.A1(W20002), .A2(W18739), .ZN(O4277));
  NOR2X1 G13899 (.A1(W13283), .A2(W7999), .ZN(W27919));
  NOR2X1 G13900 (.A1(W2920), .A2(W2811), .ZN(W7535));
  NOR2X1 G13901 (.A1(W20029), .A2(W60), .ZN(W22825));
  NOR2X1 G13902 (.A1(W6771), .A2(W8832), .ZN(O13069));
  NOR2X1 G13903 (.A1(W30498), .A2(W39052), .ZN(W43361));
  NOR2X1 G13904 (.A1(W8419), .A2(W2833), .ZN(O2619));
  NOR2X1 G13905 (.A1(W39186), .A2(W14395), .ZN(O13065));
  NOR2X1 G13906 (.A1(W40234), .A2(W26626), .ZN(O13063));
  NOR2X1 G13907 (.A1(W24448), .A2(W5827), .ZN(O4279));
  NOR2X1 G13908 (.A1(W19005), .A2(W20319), .ZN(W22820));
  NOR2X1 G13909 (.A1(W6506), .A2(W1019), .ZN(W7546));
  NOR2X1 G13910 (.A1(I554), .A2(W35781), .ZN(O13060));
  NOR2X1 G13911 (.A1(W30945), .A2(W27969), .ZN(O13700));
  NOR2X1 G13912 (.A1(W5347), .A2(W5101), .ZN(W6725));
  NOR2X1 G13913 (.A1(W2055), .A2(W10065), .ZN(O13695));
  NOR2X1 G13914 (.A1(W36298), .A2(W12943), .ZN(W44187));
  NOR2X1 G13915 (.A1(W40565), .A2(W32537), .ZN(O13698));
  NOR2X1 G13916 (.A1(I1911), .A2(I628), .ZN(W6719));
  NOR2X1 G13917 (.A1(W212), .A2(W38161), .ZN(W44192));
  NOR2X1 G13918 (.A1(W399), .A2(W5288), .ZN(O146));
  NOR2X1 G13919 (.A1(W9094), .A2(W20198), .ZN(W23100));
  NOR2X1 G13920 (.A1(W1909), .A2(W6227), .ZN(W6727));
  NOR2X1 G13921 (.A1(W17771), .A2(W11120), .ZN(W23101));
  NOR2X1 G13922 (.A1(I1514), .A2(W7349), .ZN(W23102));
  NOR2X1 G13923 (.A1(W4802), .A2(W3588), .ZN(W6711));
  NOR2X1 G13924 (.A1(W118), .A2(W5501), .ZN(W6710));
  NOR2X1 G13925 (.A1(W3426), .A2(W1590), .ZN(W6709));
  NOR2X1 G13926 (.A1(I890), .A2(W17447), .ZN(O2677));
  NOR2X1 G13927 (.A1(W8285), .A2(W4647), .ZN(W27623));
  NOR2X1 G13928 (.A1(W2858), .A2(W1185), .ZN(W6737));
  NOR2X1 G13929 (.A1(I588), .A2(W10311), .ZN(W44158));
  NOR2X1 G13930 (.A1(W28675), .A2(W40392), .ZN(O13678));
  NOR2X1 G13931 (.A1(W4832), .A2(W18968), .ZN(W44161));
  NOR2X1 G13932 (.A1(W33972), .A2(W27379), .ZN(W44162));
  NOR2X1 G13933 (.A1(W15979), .A2(W1953), .ZN(W23092));
  NOR2X1 G13934 (.A1(W15014), .A2(W10306), .ZN(O2675));
  NOR2X1 G13935 (.A1(W3689), .A2(W2415), .ZN(O149));
  NOR2X1 G13936 (.A1(W17103), .A2(W2138), .ZN(O13682));
  NOR2X1 G13937 (.A1(W998), .A2(W15336), .ZN(W27622));
  NOR2X1 G13938 (.A1(W22027), .A2(W867), .ZN(O13686));
  NOR2X1 G13939 (.A1(W26603), .A2(W18581), .ZN(W27638));
  NOR2X1 G13940 (.A1(W6099), .A2(I1688), .ZN(W6732));
  NOR2X1 G13941 (.A1(W4439), .A2(W1610), .ZN(W6731));
  NOR2X1 G13942 (.A1(W12532), .A2(W9733), .ZN(O13693));
  NOR2X1 G13943 (.A1(W6579), .A2(W6117), .ZN(W6729));
  NOR2X1 G13944 (.A1(W31704), .A2(W6499), .ZN(W44181));
  NOR2X1 G13945 (.A1(W40758), .A2(W18036), .ZN(W44247));
  NOR2X1 G13946 (.A1(W20965), .A2(W2945), .ZN(W27607));
  NOR2X1 G13947 (.A1(W23694), .A2(W41839), .ZN(O13735));
  NOR2X1 G13948 (.A1(W1560), .A2(W5571), .ZN(W6679));
  NOR2X1 G13949 (.A1(W1782), .A2(W5423), .ZN(W6678));
  NOR2X1 G13950 (.A1(W7689), .A2(W2709), .ZN(O13739));
  NOR2X1 G13951 (.A1(W25116), .A2(W36670), .ZN(O13740));
  NOR2X1 G13952 (.A1(W19774), .A2(W18214), .ZN(O13742));
  NOR2X1 G13953 (.A1(W6546), .A2(W35207), .ZN(O13743));
  NOR2X1 G13954 (.A1(W22628), .A2(W19805), .ZN(W23120));
  NOR2X1 G13955 (.A1(W37046), .A2(W20107), .ZN(W44255));
  NOR2X1 G13956 (.A1(W1331), .A2(W3175), .ZN(W6669));
  NOR2X1 G13957 (.A1(W16188), .A2(W41475), .ZN(O13753));
  NOR2X1 G13958 (.A1(W11938), .A2(W15396), .ZN(O13755));
  NOR2X1 G13959 (.A1(W6569), .A2(I1270), .ZN(W6666));
  NOR2X1 G13960 (.A1(W33773), .A2(W5054), .ZN(O13756));
  NOR2X1 G13961 (.A1(W21067), .A2(W37573), .ZN(W44263));
  NOR2X1 G13962 (.A1(W482), .A2(W22148), .ZN(O13725));
  NOR2X1 G13963 (.A1(W12333), .A2(W6305), .ZN(O13713));
  NOR2X1 G13964 (.A1(W10700), .A2(I498), .ZN(O4169));
  NOR2X1 G13965 (.A1(W5531), .A2(W8017), .ZN(O13717));
  NOR2X1 G13966 (.A1(W1670), .A2(I576), .ZN(W6696));
  NOR2X1 G13967 (.A1(W2148), .A2(W6406), .ZN(W6695));
  NOR2X1 G13968 (.A1(W5313), .A2(W1472), .ZN(O142));
  NOR2X1 G13969 (.A1(W22794), .A2(W5258), .ZN(W27615));
  NOR2X1 G13970 (.A1(W20701), .A2(W3659), .ZN(O2680));
  NOR2X1 G13971 (.A1(W15160), .A2(W32116), .ZN(O13676));
  NOR2X1 G13972 (.A1(W6801), .A2(W27537), .ZN(O13726));
  NOR2X1 G13973 (.A1(I114), .A2(W3653), .ZN(W6689));
  NOR2X1 G13974 (.A1(W13833), .A2(W13251), .ZN(W23116));
  NOR2X1 G13975 (.A1(I239), .A2(W5432), .ZN(W6687));
  NOR2X1 G13976 (.A1(W2608), .A2(W15864), .ZN(O4167));
  NOR2X1 G13977 (.A1(W10743), .A2(W133), .ZN(W27611));
  NOR2X1 G13978 (.A1(W20496), .A2(W1143), .ZN(O13731));
  NOR2X1 G13979 (.A1(W10516), .A2(W29210), .ZN(O13647));
  NOR2X1 G13980 (.A1(W924), .A2(W4177), .ZN(W6801));
  NOR2X1 G13981 (.A1(W35295), .A2(W9879), .ZN(O13637));
  NOR2X1 G13982 (.A1(W23381), .A2(W15689), .ZN(W27655));
  NOR2X1 G13983 (.A1(W26866), .A2(W18028), .ZN(O4177));
  NOR2X1 G13984 (.A1(W4343), .A2(W1353), .ZN(W6797));
  NOR2X1 G13985 (.A1(W42029), .A2(W20634), .ZN(O13644));
  NOR2X1 G13986 (.A1(W3963), .A2(W2640), .ZN(W6795));
  NOR2X1 G13987 (.A1(W3554), .A2(I1686), .ZN(W6794));
  NOR2X1 G13988 (.A1(W30476), .A2(W42510), .ZN(O13634));
  NOR2X1 G13989 (.A1(W22578), .A2(W26880), .ZN(O13648));
  NOR2X1 G13990 (.A1(W6640), .A2(W3727), .ZN(W6791));
  NOR2X1 G13991 (.A1(W12951), .A2(W13451), .ZN(O13649));
  NOR2X1 G13992 (.A1(W12868), .A2(W16549), .ZN(W27652));
  NOR2X1 G13993 (.A1(I1986), .A2(W4899), .ZN(O151));
  NOR2X1 G13994 (.A1(W10087), .A2(W19923), .ZN(W27650));
  NOR2X1 G13995 (.A1(W25650), .A2(W3790), .ZN(O13653));
  NOR2X1 G13996 (.A1(W8123), .A2(W43288), .ZN(O13627));
  NOR2X1 G13997 (.A1(I1475), .A2(W18215), .ZN(W23067));
  NOR2X1 G13998 (.A1(W16895), .A2(W56), .ZN(O13621));
  NOR2X1 G13999 (.A1(W9056), .A2(W6574), .ZN(O4184));
  NOR2X1 G14000 (.A1(W5667), .A2(W2857), .ZN(W6821));
  NOR2X1 G14001 (.A1(W41545), .A2(W18668), .ZN(O13623));
  NOR2X1 G14002 (.A1(W6579), .A2(W5042), .ZN(W6817));
  NOR2X1 G14003 (.A1(W15820), .A2(W22707), .ZN(W23071));
  NOR2X1 G14004 (.A1(W17013), .A2(W10565), .ZN(W23073));
  NOR2X1 G14005 (.A1(W19852), .A2(W15266), .ZN(W27648));
  NOR2X1 G14006 (.A1(I389), .A2(W35686), .ZN(O13628));
  NOR2X1 G14007 (.A1(W3406), .A2(W22955), .ZN(W27656));
  NOR2X1 G14008 (.A1(W26896), .A2(W34328), .ZN(O13632));
  NOR2X1 G14009 (.A1(W6585), .A2(W2051), .ZN(W6806));
  NOR2X1 G14010 (.A1(I1189), .A2(W1889), .ZN(W6805));
  NOR2X1 G14011 (.A1(W3727), .A2(W221), .ZN(W6804));
  NOR2X1 G14012 (.A1(W40128), .A2(W32823), .ZN(O13633));
  NOR2X1 G14013 (.A1(W4988), .A2(W2531), .ZN(W6756));
  NOR2X1 G14014 (.A1(W22191), .A2(W41792), .ZN(O13665));
  NOR2X1 G14015 (.A1(W5353), .A2(I1022), .ZN(W6765));
  NOR2X1 G14016 (.A1(W4215), .A2(W1065), .ZN(W6764));
  NOR2X1 G14017 (.A1(W31696), .A2(W629), .ZN(O13666));
  NOR2X1 G14018 (.A1(W10311), .A2(W25110), .ZN(W27643));
  NOR2X1 G14019 (.A1(W3190), .A2(W4361), .ZN(W6760));
  NOR2X1 G14020 (.A1(W1829), .A2(W22883), .ZN(O13668));
  NOR2X1 G14021 (.A1(W6938), .A2(W21253), .ZN(W23088));
  NOR2X1 G14022 (.A1(W27258), .A2(W5263), .ZN(O13664));
  NOR2X1 G14023 (.A1(W27387), .A2(W11240), .ZN(W44150));
  NOR2X1 G14024 (.A1(W1916), .A2(W6573), .ZN(W6753));
  NOR2X1 G14025 (.A1(W4294), .A2(I464), .ZN(W6752));
  NOR2X1 G14026 (.A1(W27028), .A2(W9417), .ZN(O13675));
  NOR2X1 G14027 (.A1(W1020), .A2(W1594), .ZN(W6750));
  NOR2X1 G14028 (.A1(W5542), .A2(W3517), .ZN(W6749));
  NOR2X1 G14029 (.A1(I237), .A2(W163), .ZN(W6748));
  NOR2X1 G14030 (.A1(W27157), .A2(W15396), .ZN(O4163));
  NOR2X1 G14031 (.A1(W39352), .A2(W25520), .ZN(O13662));
  NOR2X1 G14032 (.A1(I1563), .A2(W5213), .ZN(W6769));
  NOR2X1 G14033 (.A1(W2814), .A2(I1912), .ZN(W23084));
  NOR2X1 G14034 (.A1(W1260), .A2(I1437), .ZN(W6772));
  NOR2X1 G14035 (.A1(I124), .A2(W5689), .ZN(W6773));
  NOR2X1 G14036 (.A1(W23519), .A2(W18691), .ZN(O13660));
  NOR2X1 G14037 (.A1(W43633), .A2(W38845), .ZN(W44131));
  NOR2X1 G14038 (.A1(W13697), .A2(W30623), .ZN(O13659));
  NOR2X1 G14039 (.A1(W32477), .A2(W41531), .ZN(O13658));
  NOR2X1 G14040 (.A1(W2671), .A2(W4761), .ZN(W6779));
  NOR2X1 G14041 (.A1(I1460), .A2(W319), .ZN(W6780));
  NOR2X1 G14042 (.A1(W29474), .A2(W11129), .ZN(O13656));
  NOR2X1 G14043 (.A1(W3204), .A2(W3599), .ZN(W6782));
  NOR2X1 G14044 (.A1(W2881), .A2(W454), .ZN(O150));
  NOR2X1 G14045 (.A1(W1428), .A2(I1265), .ZN(W6784));
  NOR2X1 G14046 (.A1(W2585), .A2(I1434), .ZN(W6563));
  NOR2X1 G14047 (.A1(W15535), .A2(W17129), .ZN(W23153));
  NOR2X1 G14048 (.A1(W34612), .A2(W33958), .ZN(W44358));
  NOR2X1 G14049 (.A1(I478), .A2(I695), .ZN(W6569));
  NOR2X1 G14050 (.A1(W11513), .A2(W40945), .ZN(O13839));
  NOR2X1 G14051 (.A1(W9847), .A2(W15933), .ZN(W23154));
  NOR2X1 G14052 (.A1(W4782), .A2(W14536), .ZN(W27584));
  NOR2X1 G14053 (.A1(W38535), .A2(W26115), .ZN(W44364));
  NOR2X1 G14054 (.A1(W2831), .A2(W2214), .ZN(O136));
  NOR2X1 G14055 (.A1(I352), .A2(W18258), .ZN(W23152));
  NOR2X1 G14056 (.A1(W4900), .A2(W2120), .ZN(W6560));
  NOR2X1 G14057 (.A1(I762), .A2(W855), .ZN(W6559));
  NOR2X1 G14058 (.A1(W9137), .A2(I1254), .ZN(W27579));
  NOR2X1 G14059 (.A1(W3450), .A2(W3927), .ZN(W6557));
  NOR2X1 G14060 (.A1(W17739), .A2(W19364), .ZN(O13848));
  NOR2X1 G14061 (.A1(W3372), .A2(W4707), .ZN(O13850));
  NOR2X1 G14062 (.A1(W4855), .A2(W4647), .ZN(W6554));
  NOR2X1 G14063 (.A1(W18144), .A2(W1050), .ZN(O4156));
  NOR2X1 G14064 (.A1(W2184), .A2(W975), .ZN(W6589));
  NOR2X1 G14065 (.A1(W39288), .A2(W4959), .ZN(O13822));
  NOR2X1 G14066 (.A1(I30), .A2(W42352), .ZN(O13823));
  NOR2X1 G14067 (.A1(W20321), .A2(W3589), .ZN(O4157));
  NOR2X1 G14068 (.A1(W3665), .A2(W2320), .ZN(O2691));
  NOR2X1 G14069 (.A1(W20057), .A2(I1892), .ZN(W23147));
  NOR2X1 G14070 (.A1(W2936), .A2(W10531), .ZN(W27589));
  NOR2X1 G14071 (.A1(W33), .A2(W4625), .ZN(W6582));
  NOR2X1 G14072 (.A1(W3189), .A2(I372), .ZN(W27578));
  NOR2X1 G14073 (.A1(W6389), .A2(W2102), .ZN(O137));
  NOR2X1 G14074 (.A1(W43513), .A2(W434), .ZN(O13831));
  NOR2X1 G14075 (.A1(W5465), .A2(W5669), .ZN(W6578));
  NOR2X1 G14076 (.A1(W706), .A2(W267), .ZN(W6577));
  NOR2X1 G14077 (.A1(W4362), .A2(W4567), .ZN(O4155));
  NOR2X1 G14078 (.A1(W13483), .A2(W18977), .ZN(W44352));
  NOR2X1 G14079 (.A1(W849), .A2(W687), .ZN(W6573));
  NOR2X1 G14080 (.A1(W40078), .A2(W33989), .ZN(O13862));
  NOR2X1 G14081 (.A1(W5793), .A2(W5396), .ZN(W6534));
  NOR2X1 G14082 (.A1(W2529), .A2(W3756), .ZN(W6533));
  NOR2X1 G14083 (.A1(W4732), .A2(W3101), .ZN(W6532));
  NOR2X1 G14084 (.A1(W24345), .A2(W13830), .ZN(W27574));
  NOR2X1 G14085 (.A1(W5198), .A2(W1169), .ZN(W6530));
  NOR2X1 G14086 (.A1(W549), .A2(I1162), .ZN(W6529));
  NOR2X1 G14087 (.A1(W37148), .A2(W15631), .ZN(O13861));
  NOR2X1 G14088 (.A1(W12483), .A2(W10388), .ZN(W44388));
  NOR2X1 G14089 (.A1(I5), .A2(W3937), .ZN(O135));
  NOR2X1 G14090 (.A1(W14557), .A2(W4643), .ZN(W23168));
  NOR2X1 G14091 (.A1(W5842), .A2(W51), .ZN(W6521));
  NOR2X1 G14092 (.A1(W24434), .A2(W5094), .ZN(W44393));
  NOR2X1 G14093 (.A1(W18680), .A2(W38209), .ZN(O13865));
  NOR2X1 G14094 (.A1(W17535), .A2(W20177), .ZN(W27564));
  NOR2X1 G14095 (.A1(W22246), .A2(W40664), .ZN(W44397));
  NOR2X1 G14096 (.A1(W19268), .A2(W4043), .ZN(W23171));
  NOR2X1 G14097 (.A1(W445), .A2(W6484), .ZN(W6544));
  NOR2X1 G14098 (.A1(I981), .A2(W18816), .ZN(O4152));
  NOR2X1 G14099 (.A1(I612), .A2(W3042), .ZN(W6551));
  NOR2X1 G14100 (.A1(W24086), .A2(W16524), .ZN(W44375));
  NOR2X1 G14101 (.A1(W3060), .A2(W1449), .ZN(W6549));
  NOR2X1 G14102 (.A1(W4153), .A2(W4971), .ZN(W6548));
  NOR2X1 G14103 (.A1(W29184), .A2(W42490), .ZN(O13853));
  NOR2X1 G14104 (.A1(W670), .A2(W18781), .ZN(W23161));
  NOR2X1 G14105 (.A1(W5771), .A2(W27810), .ZN(O13855));
  NOR2X1 G14106 (.A1(W6394), .A2(W21036), .ZN(W23144));
  NOR2X1 G14107 (.A1(W4764), .A2(W4951), .ZN(W6543));
  NOR2X1 G14108 (.A1(W2816), .A2(W5063), .ZN(W6542));
  NOR2X1 G14109 (.A1(W3812), .A2(W5219), .ZN(W6541));
  NOR2X1 G14110 (.A1(W21303), .A2(W6878), .ZN(O2694));
  NOR2X1 G14111 (.A1(W2334), .A2(W1395), .ZN(W6539));
  NOR2X1 G14112 (.A1(W2316), .A2(W2418), .ZN(W6538));
  NOR2X1 G14113 (.A1(W5462), .A2(W5464), .ZN(W6537));
  NOR2X1 G14114 (.A1(W738), .A2(W1694), .ZN(W6636));
  NOR2X1 G14115 (.A1(W29723), .A2(W26696), .ZN(O13780));
  NOR2X1 G14116 (.A1(W6225), .A2(W697), .ZN(W6644));
  NOR2X1 G14117 (.A1(W980), .A2(W1888), .ZN(W44289));
  NOR2X1 G14118 (.A1(W1679), .A2(W1508), .ZN(W6642));
  NOR2X1 G14119 (.A1(W16032), .A2(W7619), .ZN(O13783));
  NOR2X1 G14120 (.A1(I1339), .A2(W42570), .ZN(O13785));
  NOR2X1 G14121 (.A1(W904), .A2(I1664), .ZN(W6638));
  NOR2X1 G14122 (.A1(W620), .A2(W3962), .ZN(W6637));
  NOR2X1 G14123 (.A1(W3480), .A2(W6292), .ZN(W6646));
  NOR2X1 G14124 (.A1(W2809), .A2(W5678), .ZN(W6635));
  NOR2X1 G14125 (.A1(W1112), .A2(I338), .ZN(W6634));
  NOR2X1 G14126 (.A1(W2201), .A2(W5778), .ZN(W6633));
  NOR2X1 G14127 (.A1(W3216), .A2(W1022), .ZN(W6632));
  NOR2X1 G14128 (.A1(W1574), .A2(W10064), .ZN(O2683));
  NOR2X1 G14129 (.A1(W449), .A2(W5724), .ZN(W6630));
  NOR2X1 G14130 (.A1(W43022), .A2(W9565), .ZN(O13788));
  NOR2X1 G14131 (.A1(W11940), .A2(W36201), .ZN(O13772));
  NOR2X1 G14132 (.A1(W34066), .A2(W5614), .ZN(O13760));
  NOR2X1 G14133 (.A1(W5526), .A2(W769), .ZN(W6661));
  NOR2X1 G14134 (.A1(W2605), .A2(W26823), .ZN(O13762));
  NOR2X1 G14135 (.A1(W8325), .A2(W419), .ZN(W23125));
  NOR2X1 G14136 (.A1(W2467), .A2(W10268), .ZN(W23126));
  NOR2X1 G14137 (.A1(W13212), .A2(W7787), .ZN(W23127));
  NOR2X1 G14138 (.A1(W4140), .A2(W1713), .ZN(W23128));
  NOR2X1 G14139 (.A1(W25964), .A2(W31793), .ZN(O13771));
  NOR2X1 G14140 (.A1(W6584), .A2(W3372), .ZN(W6628));
  NOR2X1 G14141 (.A1(W586), .A2(W4094), .ZN(W6653));
  NOR2X1 G14142 (.A1(W5730), .A2(W2168), .ZN(W6652));
  NOR2X1 G14143 (.A1(W11595), .A2(W19867), .ZN(O13775));
  NOR2X1 G14144 (.A1(W12423), .A2(W21231), .ZN(W23129));
  NOR2X1 G14145 (.A1(W4622), .A2(W1250), .ZN(W6649));
  NOR2X1 G14146 (.A1(W15962), .A2(W42594), .ZN(O13779));
  NOR2X1 G14147 (.A1(I1158), .A2(W719), .ZN(W6647));
  NOR2X1 G14148 (.A1(W24442), .A2(W28428), .ZN(O13813));
  NOR2X1 G14149 (.A1(W635), .A2(W3680), .ZN(W6608));
  NOR2X1 G14150 (.A1(W22642), .A2(W17858), .ZN(O2685));
  NOR2X1 G14151 (.A1(W42872), .A2(W21487), .ZN(W44326));
  NOR2X1 G14152 (.A1(W1029), .A2(W12063), .ZN(O2686));
  NOR2X1 G14153 (.A1(I612), .A2(W4310), .ZN(W6604));
  NOR2X1 G14154 (.A1(I1501), .A2(W5635), .ZN(W6603));
  NOR2X1 G14155 (.A1(I839), .A2(W646), .ZN(W6602));
  NOR2X1 G14156 (.A1(I481), .A2(W4241), .ZN(W6601));
  NOR2X1 G14157 (.A1(W6156), .A2(W26716), .ZN(O13805));
  NOR2X1 G14158 (.A1(W6081), .A2(W13595), .ZN(W27596));
  NOR2X1 G14159 (.A1(W826), .A2(I6), .ZN(O2688));
  NOR2X1 G14160 (.A1(W2850), .A2(W1703), .ZN(W23141));
  NOR2X1 G14161 (.A1(W13718), .A2(W25489), .ZN(O13818));
  NOR2X1 G14162 (.A1(W1074), .A2(W1656), .ZN(W6594));
  NOR2X1 G14163 (.A1(W1340), .A2(W2823), .ZN(W6592));
  NOR2X1 G14164 (.A1(W33525), .A2(W26501), .ZN(W44337));
  NOR2X1 G14165 (.A1(W35617), .A2(W41196), .ZN(O13619));
  NOR2X1 G14166 (.A1(W16729), .A2(W4395), .ZN(O4161));
  NOR2X1 G14167 (.A1(W24376), .A2(W14610), .ZN(O13799));
  NOR2X1 G14168 (.A1(W2380), .A2(W2951), .ZN(W6614));
  NOR2X1 G14169 (.A1(W2872), .A2(W1387), .ZN(W6615));
  NOR2X1 G14170 (.A1(W4183), .A2(I1495), .ZN(W6616));
  NOR2X1 G14171 (.A1(I51), .A2(W7870), .ZN(W23133));
  NOR2X1 G14172 (.A1(W4543), .A2(W5658), .ZN(W6618));
  NOR2X1 G14173 (.A1(W11777), .A2(W23327), .ZN(O13798));
  NOR2X1 G14174 (.A1(W2190), .A2(W4465), .ZN(O13797));
  NOR2X1 G14175 (.A1(W1346), .A2(W5457), .ZN(W6622));
  NOR2X1 G14176 (.A1(W6512), .A2(I1463), .ZN(W6623));
  NOR2X1 G14177 (.A1(W40709), .A2(W44091), .ZN(W44307));
  NOR2X1 G14178 (.A1(W2779), .A2(W21493), .ZN(W44305));
  NOR2X1 G14179 (.A1(W3831), .A2(W1181), .ZN(W6626));
  NOR2X1 G14180 (.A1(W22232), .A2(W28540), .ZN(O13793));
  NOR2X1 G14181 (.A1(W30652), .A2(W35850), .ZN(W43864));
  NOR2X1 G14182 (.A1(W6058), .A2(W3234), .ZN(W7037));
  NOR2X1 G14183 (.A1(W24175), .A2(W5160), .ZN(O4217));
  NOR2X1 G14184 (.A1(W3531), .A2(W835), .ZN(W7033));
  NOR2X1 G14185 (.A1(W6288), .A2(W5799), .ZN(W7031));
  NOR2X1 G14186 (.A1(W4246), .A2(W16690), .ZN(O2654));
  NOR2X1 G14187 (.A1(W252), .A2(I1893), .ZN(W7029));
  NOR2X1 G14188 (.A1(W1490), .A2(W19274), .ZN(O2656));
  NOR2X1 G14189 (.A1(W28914), .A2(W6993), .ZN(O13444));
  NOR2X1 G14190 (.A1(W12384), .A2(W15279), .ZN(W43848));
  NOR2X1 G14191 (.A1(W19472), .A2(W36402), .ZN(O13445));
  NOR2X1 G14192 (.A1(I1355), .A2(W2876), .ZN(W7023));
  NOR2X1 G14193 (.A1(I1003), .A2(W25803), .ZN(O13446));
  NOR2X1 G14194 (.A1(W13276), .A2(W7927), .ZN(O13447));
  NOR2X1 G14195 (.A1(W5914), .A2(W1519), .ZN(W7020));
  NOR2X1 G14196 (.A1(W4351), .A2(W3738), .ZN(W7018));
  NOR2X1 G14197 (.A1(W12182), .A2(W22106), .ZN(O13450));
  NOR2X1 G14198 (.A1(W33613), .A2(W32469), .ZN(O13425));
  NOR2X1 G14199 (.A1(W37388), .A2(W20345), .ZN(O13420));
  NOR2X1 G14200 (.A1(W2182), .A2(W5698), .ZN(W7057));
  NOR2X1 G14201 (.A1(W2376), .A2(I1729), .ZN(W7056));
  NOR2X1 G14202 (.A1(W18243), .A2(W1917), .ZN(W27754));
  NOR2X1 G14203 (.A1(W38213), .A2(W34625), .ZN(O13422));
  NOR2X1 G14204 (.A1(W1258), .A2(W5783), .ZN(W7052));
  NOR2X1 G14205 (.A1(W36858), .A2(I1772), .ZN(O13423));
  NOR2X1 G14206 (.A1(W2715), .A2(W4198), .ZN(W7049));
  NOR2X1 G14207 (.A1(I1958), .A2(I1629), .ZN(O159));
  NOR2X1 G14208 (.A1(W22975), .A2(W23648), .ZN(O13426));
  NOR2X1 G14209 (.A1(W826), .A2(W22684), .ZN(W43843));
  NOR2X1 G14210 (.A1(W5933), .A2(W22769), .ZN(O13428));
  NOR2X1 G14211 (.A1(W7115), .A2(W32497), .ZN(O13429));
  NOR2X1 G14212 (.A1(W3927), .A2(W6919), .ZN(W7041));
  NOR2X1 G14213 (.A1(W601), .A2(W1651), .ZN(W7040));
  NOR2X1 G14214 (.A1(W16927), .A2(W32637), .ZN(O13430));
  NOR2X1 G14215 (.A1(W409), .A2(W12908), .ZN(W23008));
  NOR2X1 G14216 (.A1(W21114), .A2(W7156), .ZN(O13471));
  NOR2X1 G14217 (.A1(W297), .A2(W17925), .ZN(O13472));
  NOR2X1 G14218 (.A1(W35129), .A2(W35747), .ZN(O13475));
  NOR2X1 G14219 (.A1(W30150), .A2(W11051), .ZN(O13476));
  NOR2X1 G14220 (.A1(W43556), .A2(W8451), .ZN(O13477));
  NOR2X1 G14221 (.A1(W11217), .A2(W5483), .ZN(O4214));
  NOR2X1 G14222 (.A1(W24534), .A2(W41833), .ZN(O13479));
  NOR2X1 G14223 (.A1(W4105), .A2(W4545), .ZN(W6990));
  NOR2X1 G14224 (.A1(W1187), .A2(W3850), .ZN(W6998));
  NOR2X1 G14225 (.A1(W1809), .A2(W3910), .ZN(W6987));
  NOR2X1 G14226 (.A1(W1067), .A2(W1306), .ZN(W6986));
  NOR2X1 G14227 (.A1(W35624), .A2(W7155), .ZN(O13486));
  NOR2X1 G14228 (.A1(W26435), .A2(W40154), .ZN(O13487));
  NOR2X1 G14229 (.A1(W11180), .A2(W19230), .ZN(W23010));
  NOR2X1 G14230 (.A1(W28451), .A2(W24437), .ZN(O13489));
  NOR2X1 G14231 (.A1(W14928), .A2(W21833), .ZN(W23011));
  NOR2X1 G14232 (.A1(W17148), .A2(W4324), .ZN(O2657));
  NOR2X1 G14233 (.A1(W5920), .A2(W18615), .ZN(O13452));
  NOR2X1 G14234 (.A1(W32656), .A2(W34552), .ZN(O13454));
  NOR2X1 G14235 (.A1(I926), .A2(W3870), .ZN(W7012));
  NOR2X1 G14236 (.A1(W42630), .A2(W31844), .ZN(O13457));
  NOR2X1 G14237 (.A1(W14000), .A2(W13033), .ZN(O4215));
  NOR2X1 G14238 (.A1(W4792), .A2(W3369), .ZN(W7009));
  NOR2X1 G14239 (.A1(W21421), .A2(W6114), .ZN(W23003));
  NOR2X1 G14240 (.A1(W5791), .A2(W35625), .ZN(O13462));
  NOR2X1 G14241 (.A1(W9664), .A2(W19306), .ZN(O13418));
  NOR2X1 G14242 (.A1(W30713), .A2(W43208), .ZN(W43885));
  NOR2X1 G14243 (.A1(W22253), .A2(W17890), .ZN(O13463));
  NOR2X1 G14244 (.A1(W17100), .A2(W5284), .ZN(W43889));
  NOR2X1 G14245 (.A1(W1334), .A2(W4880), .ZN(W7002));
  NOR2X1 G14246 (.A1(W30686), .A2(W38088), .ZN(O15148));
  NOR2X1 G14247 (.A1(W10528), .A2(W17169), .ZN(O2658));
  NOR2X1 G14248 (.A1(W3851), .A2(W23675), .ZN(W27740));
  NOR2X1 G14249 (.A1(W1917), .A2(W2255), .ZN(W7105));
  NOR2X1 G14250 (.A1(W1729), .A2(W983), .ZN(W7113));
  NOR2X1 G14251 (.A1(W4466), .A2(W1892), .ZN(W7112));
  NOR2X1 G14252 (.A1(W2957), .A2(W1885), .ZN(W7111));
  NOR2X1 G14253 (.A1(W7228), .A2(W21641), .ZN(O4223));
  NOR2X1 G14254 (.A1(I1739), .A2(W1519), .ZN(W7109));
  NOR2X1 G14255 (.A1(W21081), .A2(W14415), .ZN(O13384));
  NOR2X1 G14256 (.A1(I1726), .A2(W4087), .ZN(O13385));
  NOR2X1 G14257 (.A1(W3667), .A2(W4605), .ZN(W7106));
  NOR2X1 G14258 (.A1(W3155), .A2(W2103), .ZN(W7114));
  NOR2X1 G14259 (.A1(W4244), .A2(W981), .ZN(W7103));
  NOR2X1 G14260 (.A1(W8256), .A2(W40833), .ZN(O13387));
  NOR2X1 G14261 (.A1(W9108), .A2(W23542), .ZN(O13389));
  NOR2X1 G14262 (.A1(W2902), .A2(W1760), .ZN(W7100));
  NOR2X1 G14263 (.A1(W18047), .A2(W21742), .ZN(W22969));
  NOR2X1 G14264 (.A1(W22108), .A2(W17581), .ZN(W27765));
  NOR2X1 G14265 (.A1(W13751), .A2(W29996), .ZN(O13392));
  NOR2X1 G14266 (.A1(I1600), .A2(I1273), .ZN(W7125));
  NOR2X1 G14267 (.A1(W2824), .A2(W6494), .ZN(W7136));
  NOR2X1 G14268 (.A1(W7898), .A2(W37301), .ZN(W43756));
  NOR2X1 G14269 (.A1(W5809), .A2(W666), .ZN(W7133));
  NOR2X1 G14270 (.A1(W8859), .A2(W20590), .ZN(W43759));
  NOR2X1 G14271 (.A1(I1164), .A2(W6164), .ZN(O4230));
  NOR2X1 G14272 (.A1(W30222), .A2(W998), .ZN(O13365));
  NOR2X1 G14273 (.A1(I1804), .A2(W3859), .ZN(W7129));
  NOR2X1 G14274 (.A1(W20677), .A2(W8816), .ZN(O13366));
  NOR2X1 G14275 (.A1(W6620), .A2(W2856), .ZN(W7096));
  NOR2X1 G14276 (.A1(W16861), .A2(W2532), .ZN(O4225));
  NOR2X1 G14277 (.A1(W35989), .A2(W38466), .ZN(O13370));
  NOR2X1 G14278 (.A1(W14360), .A2(W85), .ZN(W27771));
  NOR2X1 G14279 (.A1(W3969), .A2(I635), .ZN(W7120));
  NOR2X1 G14280 (.A1(I824), .A2(W2296), .ZN(W7119));
  NOR2X1 G14281 (.A1(W9550), .A2(W17616), .ZN(W22964));
  NOR2X1 G14282 (.A1(W7498), .A2(W22639), .ZN(O2646));
  NOR2X1 G14283 (.A1(I563), .A2(W1463), .ZN(W7067));
  NOR2X1 G14284 (.A1(W15045), .A2(W19789), .ZN(W22981));
  NOR2X1 G14285 (.A1(I320), .A2(W2073), .ZN(W7075));
  NOR2X1 G14286 (.A1(W5913), .A2(W5230), .ZN(W7074));
  NOR2X1 G14287 (.A1(W3146), .A2(W18886), .ZN(W27757));
  NOR2X1 G14288 (.A1(W3065), .A2(W6040), .ZN(W7072));
  NOR2X1 G14289 (.A1(W21979), .A2(I861), .ZN(O13409));
  NOR2X1 G14290 (.A1(W4204), .A2(I1622), .ZN(W7069));
  NOR2X1 G14291 (.A1(W20329), .A2(W11313), .ZN(O4220));
  NOR2X1 G14292 (.A1(W31157), .A2(W27944), .ZN(O13406));
  NOR2X1 G14293 (.A1(W8344), .A2(W2963), .ZN(W22985));
  NOR2X1 G14294 (.A1(W1017), .A2(W6532), .ZN(W7065));
  NOR2X1 G14295 (.A1(W2666), .A2(W6981), .ZN(W22986));
  NOR2X1 G14296 (.A1(W12054), .A2(W17174), .ZN(O13415));
  NOR2X1 G14297 (.A1(W8), .A2(I1140), .ZN(W7062));
  NOR2X1 G14298 (.A1(W2922), .A2(W17328), .ZN(O2651));
  NOR2X1 G14299 (.A1(W21677), .A2(W34676), .ZN(O13417));
  NOR2X1 G14300 (.A1(W12176), .A2(W10171), .ZN(W23013));
  NOR2X1 G14301 (.A1(W20046), .A2(W2609), .ZN(W22978));
  NOR2X1 G14302 (.A1(W6821), .A2(I203), .ZN(W7081));
  NOR2X1 G14303 (.A1(W1196), .A2(W2326), .ZN(W43808));
  NOR2X1 G14304 (.A1(W1926), .A2(I252), .ZN(W7083));
  NOR2X1 G14305 (.A1(W1258), .A2(W3421), .ZN(W7084));
  NOR2X1 G14306 (.A1(W13435), .A2(W40378), .ZN(O13403));
  NOR2X1 G14307 (.A1(W8366), .A2(I1028), .ZN(W22977));
  NOR2X1 G14308 (.A1(W6365), .A2(W14052), .ZN(O4221));
  NOR2X1 G14309 (.A1(W20899), .A2(W20771), .ZN(W22975));
  NOR2X1 G14310 (.A1(W1471), .A2(W22759), .ZN(O13398));
  NOR2X1 G14311 (.A1(I1407), .A2(W2649), .ZN(W7090));
  NOR2X1 G14312 (.A1(W4680), .A2(W20324), .ZN(W27761));
  NOR2X1 G14313 (.A1(W9259), .A2(W369), .ZN(O4222));
  NOR2X1 G14314 (.A1(W38381), .A2(W21850), .ZN(O13395));
  NOR2X1 G14315 (.A1(W10100), .A2(W6200), .ZN(O2648));
  NOR2X1 G14316 (.A1(W16953), .A2(W16994), .ZN(O13577));
  NOR2X1 G14317 (.A1(I1806), .A2(W16408), .ZN(W44029));
  NOR2X1 G14318 (.A1(W2824), .A2(W1280), .ZN(W6880));
  NOR2X1 G14319 (.A1(W15449), .A2(W34843), .ZN(O13575));
  NOR2X1 G14320 (.A1(W32013), .A2(W40566), .ZN(W44031));
  NOR2X1 G14321 (.A1(W4644), .A2(W3350), .ZN(W6877));
  NOR2X1 G14322 (.A1(W21315), .A2(W41266), .ZN(O13576));
  NOR2X1 G14323 (.A1(W1516), .A2(W2951), .ZN(W6875));
  NOR2X1 G14324 (.A1(W1014), .A2(W3272), .ZN(W6874));
  NOR2X1 G14325 (.A1(W39890), .A2(W41990), .ZN(O13574));
  NOR2X1 G14326 (.A1(W1865), .A2(I122), .ZN(O4195));
  NOR2X1 G14327 (.A1(W33944), .A2(W19642), .ZN(W44035));
  NOR2X1 G14328 (.A1(W40747), .A2(W6504), .ZN(O13578));
  NOR2X1 G14329 (.A1(W11910), .A2(W22194), .ZN(W23049));
  NOR2X1 G14330 (.A1(W5791), .A2(W20892), .ZN(W23050));
  NOR2X1 G14331 (.A1(W5598), .A2(I210), .ZN(W6867));
  NOR2X1 G14332 (.A1(W13026), .A2(W10713), .ZN(O4194));
  NOR2X1 G14333 (.A1(W37582), .A2(W17687), .ZN(W44018));
  NOR2X1 G14334 (.A1(W22961), .A2(W17714), .ZN(O4198));
  NOR2X1 G14335 (.A1(W1328), .A2(W1977), .ZN(W23043));
  NOR2X1 G14336 (.A1(W17827), .A2(W7441), .ZN(W27695));
  NOR2X1 G14337 (.A1(W6446), .A2(W2562), .ZN(W6895));
  NOR2X1 G14338 (.A1(W27204), .A2(W42681), .ZN(O13563));
  NOR2X1 G14339 (.A1(W5470), .A2(W21824), .ZN(W27694));
  NOR2X1 G14340 (.A1(W2730), .A2(W6072), .ZN(W6892));
  NOR2X1 G14341 (.A1(W11325), .A2(I462), .ZN(W23046));
  NOR2X1 G14342 (.A1(W4478), .A2(I811), .ZN(W6865));
  NOR2X1 G14343 (.A1(W11655), .A2(W7616), .ZN(O13569));
  NOR2X1 G14344 (.A1(W6090), .A2(W6398), .ZN(W6888));
  NOR2X1 G14345 (.A1(W615), .A2(W3656), .ZN(W6887));
  NOR2X1 G14346 (.A1(W39276), .A2(W9425), .ZN(O13571));
  NOR2X1 G14347 (.A1(W7731), .A2(W18173), .ZN(O4196));
  NOR2X1 G14348 (.A1(W27160), .A2(W1317), .ZN(O13573));
  NOR2X1 G14349 (.A1(W2729), .A2(I324), .ZN(O154));
  NOR2X1 G14350 (.A1(W1105), .A2(W7693), .ZN(O13604));
  NOR2X1 G14351 (.A1(W4240), .A2(W1875), .ZN(W6847));
  NOR2X1 G14352 (.A1(W17135), .A2(W20824), .ZN(W27683));
  NOR2X1 G14353 (.A1(W1116), .A2(I1470), .ZN(W6845));
  NOR2X1 G14354 (.A1(W1118), .A2(W8184), .ZN(W27678));
  NOR2X1 G14355 (.A1(W6685), .A2(W1702), .ZN(W6842));
  NOR2X1 G14356 (.A1(W42003), .A2(W4759), .ZN(O13602));
  NOR2X1 G14357 (.A1(W922), .A2(W2363), .ZN(W6840));
  NOR2X1 G14358 (.A1(I459), .A2(W6321), .ZN(W6838));
  NOR2X1 G14359 (.A1(W5546), .A2(W6291), .ZN(W6848));
  NOR2X1 G14360 (.A1(W2396), .A2(W1702), .ZN(W6836));
  NOR2X1 G14361 (.A1(W3915), .A2(W1773), .ZN(O13606));
  NOR2X1 G14362 (.A1(W40470), .A2(W5033), .ZN(O13607));
  NOR2X1 G14363 (.A1(W11586), .A2(W22806), .ZN(O2671));
  NOR2X1 G14364 (.A1(W9202), .A2(I1986), .ZN(O4185));
  NOR2X1 G14365 (.A1(W389), .A2(W2201), .ZN(W23065));
  NOR2X1 G14366 (.A1(W7945), .A2(W41221), .ZN(O13618));
  NOR2X1 G14367 (.A1(W4877), .A2(W4212), .ZN(W6899));
  NOR2X1 G14368 (.A1(W21967), .A2(W5802), .ZN(W23055));
  NOR2X1 G14369 (.A1(W6142), .A2(W3350), .ZN(W6850));
  NOR2X1 G14370 (.A1(I908), .A2(W5090), .ZN(W6851));
  NOR2X1 G14371 (.A1(W6700), .A2(W1795), .ZN(W6853));
  NOR2X1 G14372 (.A1(W17859), .A2(W12032), .ZN(O13593));
  NOR2X1 G14373 (.A1(W4490), .A2(I237), .ZN(W6855));
  NOR2X1 G14374 (.A1(W17653), .A2(W23667), .ZN(O13592));
  NOR2X1 G14375 (.A1(W2211), .A2(I1271), .ZN(W6857));
  NOR2X1 G14376 (.A1(W3714), .A2(W384), .ZN(W27686));
  NOR2X1 G14377 (.A1(W27410), .A2(W6849), .ZN(O4192));
  NOR2X1 G14378 (.A1(W14686), .A2(W23248), .ZN(O13587));
  NOR2X1 G14379 (.A1(W38270), .A2(W31982), .ZN(O13585));
  NOR2X1 G14380 (.A1(W271), .A2(W41613), .ZN(O13584));
  NOR2X1 G14381 (.A1(W4213), .A2(W2079), .ZN(W6863));
  NOR2X1 G14382 (.A1(W13834), .A2(W12963), .ZN(W44041));
  NOR2X1 G14383 (.A1(W37122), .A2(W17789), .ZN(O13526));
  NOR2X1 G14384 (.A1(W11611), .A2(W19563), .ZN(W27717));
  NOR2X1 G14385 (.A1(W25213), .A2(W22262), .ZN(O4207));
  NOR2X1 G14386 (.A1(W12170), .A2(W1123), .ZN(O13523));
  NOR2X1 G14387 (.A1(W13873), .A2(W11558), .ZN(O4206));
  NOR2X1 G14388 (.A1(W3231), .A2(I1924), .ZN(W6947));
  NOR2X1 G14389 (.A1(W1693), .A2(W3447), .ZN(W6946));
  NOR2X1 G14390 (.A1(W27787), .A2(W7375), .ZN(O13525));
  NOR2X1 G14391 (.A1(W35063), .A2(W466), .ZN(W43967));
  NOR2X1 G14392 (.A1(W2876), .A2(W32791), .ZN(O13516));
  NOR2X1 G14393 (.A1(W37702), .A2(W9172), .ZN(O13527));
  NOR2X1 G14394 (.A1(W3339), .A2(W936), .ZN(W6941));
  NOR2X1 G14395 (.A1(W12442), .A2(W15451), .ZN(O4205));
  NOR2X1 G14396 (.A1(I368), .A2(W5877), .ZN(W6939));
  NOR2X1 G14397 (.A1(W22720), .A2(W6951), .ZN(O13529));
  NOR2X1 G14398 (.A1(W5189), .A2(W18497), .ZN(W27709));
  NOR2X1 G14399 (.A1(W911), .A2(W226), .ZN(W6936));
  NOR2X1 G14400 (.A1(W244), .A2(I1256), .ZN(W6965));
  NOR2X1 G14401 (.A1(W6001), .A2(W340), .ZN(W6978));
  NOR2X1 G14402 (.A1(W25280), .A2(W14577), .ZN(W27733));
  NOR2X1 G14403 (.A1(W6939), .A2(W6032), .ZN(W6974));
  NOR2X1 G14404 (.A1(W2927), .A2(W257), .ZN(W6971));
  NOR2X1 G14405 (.A1(I917), .A2(W5825), .ZN(W6970));
  NOR2X1 G14406 (.A1(W3629), .A2(I960), .ZN(W6969));
  NOR2X1 G14407 (.A1(I1420), .A2(W20443), .ZN(O13498));
  NOR2X1 G14408 (.A1(W851), .A2(W7966), .ZN(O13501));
  NOR2X1 G14409 (.A1(W14771), .A2(W37681), .ZN(O13531));
  NOR2X1 G14410 (.A1(W3607), .A2(W31274), .ZN(W43937));
  NOR2X1 G14411 (.A1(W33643), .A2(W25469), .ZN(O13505));
  NOR2X1 G14412 (.A1(W33681), .A2(W11375), .ZN(W43942));
  NOR2X1 G14413 (.A1(I1055), .A2(W6736), .ZN(W6959));
  NOR2X1 G14414 (.A1(W20858), .A2(W26449), .ZN(O13508));
  NOR2X1 G14415 (.A1(W26173), .A2(W41734), .ZN(O13511));
  NOR2X1 G14416 (.A1(W3262), .A2(W639), .ZN(O4211));
  NOR2X1 G14417 (.A1(W9397), .A2(W917), .ZN(W27699));
  NOR2X1 G14418 (.A1(W21405), .A2(W27410), .ZN(O13546));
  NOR2X1 G14419 (.A1(W43439), .A2(W26077), .ZN(O13547));
  NOR2X1 G14420 (.A1(W3774), .A2(W2325), .ZN(O156));
  NOR2X1 G14421 (.A1(I1763), .A2(W37027), .ZN(O13549));
  NOR2X1 G14422 (.A1(I1361), .A2(W6955), .ZN(W23036));
  NOR2X1 G14423 (.A1(W21615), .A2(I1590), .ZN(O2666));
  NOR2X1 G14424 (.A1(I185), .A2(I1579), .ZN(W6910));
  NOR2X1 G14425 (.A1(W780), .A2(W2594), .ZN(W6908));
  NOR2X1 G14426 (.A1(I1480), .A2(I1489), .ZN(W6917));
  NOR2X1 G14427 (.A1(W7250), .A2(W20058), .ZN(O13556));
  NOR2X1 G14428 (.A1(W33252), .A2(W27599), .ZN(O13557));
  NOR2X1 G14429 (.A1(W1027), .A2(W289), .ZN(W6904));
  NOR2X1 G14430 (.A1(W15496), .A2(W1317), .ZN(O4200));
  NOR2X1 G14431 (.A1(W14771), .A2(W23474), .ZN(O4199));
  NOR2X1 G14432 (.A1(I737), .A2(W1014), .ZN(W6901));
  NOR2X1 G14433 (.A1(W30151), .A2(W29700), .ZN(O13559));
  NOR2X1 G14434 (.A1(W2402), .A2(W2651), .ZN(W7742));
  NOR2X1 G14435 (.A1(W5586), .A2(W6793), .ZN(W6918));
  NOR2X1 G14436 (.A1(W2803), .A2(W676), .ZN(W6919));
  NOR2X1 G14437 (.A1(W29710), .A2(W13631), .ZN(O13542));
  NOR2X1 G14438 (.A1(W2092), .A2(W8869), .ZN(O13541));
  NOR2X1 G14439 (.A1(W2851), .A2(W5455), .ZN(W6923));
  NOR2X1 G14440 (.A1(W2239), .A2(W3085), .ZN(W6924));
  NOR2X1 G14441 (.A1(W3210), .A2(W6938), .ZN(W43986));
  NOR2X1 G14442 (.A1(I112), .A2(W41589), .ZN(O13538));
  NOR2X1 G14443 (.A1(W22626), .A2(W13141), .ZN(W23033));
  NOR2X1 G14444 (.A1(W7895), .A2(W226), .ZN(W23032));
  NOR2X1 G14445 (.A1(W6406), .A2(W7972), .ZN(W27706));
  NOR2X1 G14446 (.A1(W33876), .A2(W24407), .ZN(O13536));
  NOR2X1 G14447 (.A1(W35486), .A2(W30554), .ZN(O13535));
  NOR2X1 G14448 (.A1(W22241), .A2(W14509), .ZN(O13533));
  NOR2X1 G14449 (.A1(W3085), .A2(W214), .ZN(W6934));
  NOR2X1 G14450 (.A1(W24453), .A2(W12185), .ZN(W28255));
  NOR2X1 G14451 (.A1(W5049), .A2(W19394), .ZN(W22477));
  NOR2X1 G14452 (.A1(W2994), .A2(W5630), .ZN(W8538));
  NOR2X1 G14453 (.A1(I1366), .A2(I356), .ZN(W8536));
  NOR2X1 G14454 (.A1(I1133), .A2(W8440), .ZN(W8534));
  NOR2X1 G14455 (.A1(W7588), .A2(I266), .ZN(W8533));
  NOR2X1 G14456 (.A1(W2845), .A2(W1615), .ZN(O2528));
  NOR2X1 G14457 (.A1(W38757), .A2(W41523), .ZN(O12282));
  NOR2X1 G14458 (.A1(W2094), .A2(W20837), .ZN(W22481));
  NOR2X1 G14459 (.A1(W3196), .A2(W562), .ZN(W8540));
  NOR2X1 G14460 (.A1(W13198), .A2(W13129), .ZN(W28254));
  NOR2X1 G14461 (.A1(W5218), .A2(W4438), .ZN(O234));
  NOR2X1 G14462 (.A1(W33391), .A2(W11929), .ZN(W42364));
  NOR2X1 G14463 (.A1(W1025), .A2(W928), .ZN(W8525));
  NOR2X1 G14464 (.A1(I1698), .A2(W3129), .ZN(W8524));
  NOR2X1 G14465 (.A1(W7423), .A2(W2147), .ZN(W8523));
  NOR2X1 G14466 (.A1(W4487), .A2(I1750), .ZN(W8522));
  NOR2X1 G14467 (.A1(I1367), .A2(W20044), .ZN(O2524));
  NOR2X1 G14468 (.A1(I1167), .A2(I294), .ZN(W8556));
  NOR2X1 G14469 (.A1(W40045), .A2(W14976), .ZN(O12270));
  NOR2X1 G14470 (.A1(I13), .A2(W8008), .ZN(W8554));
  NOR2X1 G14471 (.A1(I1606), .A2(W6323), .ZN(O12271));
  NOR2X1 G14472 (.A1(W11785), .A2(W13724), .ZN(O2523));
  NOR2X1 G14473 (.A1(W6233), .A2(W4372), .ZN(W8551));
  NOR2X1 G14474 (.A1(W81), .A2(W3224), .ZN(W8550));
  NOR2X1 G14475 (.A1(W1337), .A2(W6046), .ZN(W8549));
  NOR2X1 G14476 (.A1(W5233), .A2(W2541), .ZN(W8521));
  NOR2X1 G14477 (.A1(I1020), .A2(W32201), .ZN(W42344));
  NOR2X1 G14478 (.A1(W8412), .A2(I72), .ZN(W8546));
  NOR2X1 G14479 (.A1(W4903), .A2(W8248), .ZN(W8545));
  NOR2X1 G14480 (.A1(W4518), .A2(W7531), .ZN(W8544));
  NOR2X1 G14481 (.A1(W22271), .A2(W6933), .ZN(O2525));
  NOR2X1 G14482 (.A1(W1893), .A2(W34812), .ZN(O12276));
  NOR2X1 G14483 (.A1(W5794), .A2(W2822), .ZN(O2526));
  NOR2X1 G14484 (.A1(W7524), .A2(W4922), .ZN(W8493));
  NOR2X1 G14485 (.A1(W4552), .A2(W11095), .ZN(O12294));
  NOR2X1 G14486 (.A1(W6929), .A2(W3028), .ZN(W8501));
  NOR2X1 G14487 (.A1(W13474), .A2(W18061), .ZN(W22490));
  NOR2X1 G14488 (.A1(W29548), .A2(W26863), .ZN(W42385));
  NOR2X1 G14489 (.A1(W6099), .A2(W5204), .ZN(W8498));
  NOR2X1 G14490 (.A1(W15265), .A2(W2049), .ZN(O2531));
  NOR2X1 G14491 (.A1(W7923), .A2(W27183), .ZN(O12300));
  NOR2X1 G14492 (.A1(W19537), .A2(W33323), .ZN(O12301));
  NOR2X1 G14493 (.A1(W21400), .A2(W10854), .ZN(W22489));
  NOR2X1 G14494 (.A1(W10789), .A2(W16231), .ZN(O12303));
  NOR2X1 G14495 (.A1(W1406), .A2(W532), .ZN(W8491));
  NOR2X1 G14496 (.A1(W7017), .A2(W3728), .ZN(W8490));
  NOR2X1 G14497 (.A1(W9028), .A2(W10881), .ZN(O12305));
  NOR2X1 G14498 (.A1(W6130), .A2(W6740), .ZN(W8487));
  NOR2X1 G14499 (.A1(W7114), .A2(W5441), .ZN(W8486));
  NOR2X1 G14500 (.A1(W7103), .A2(I1621), .ZN(W8485));
  NOR2X1 G14501 (.A1(W2203), .A2(W8427), .ZN(W28253));
  NOR2X1 G14502 (.A1(I117), .A2(W28599), .ZN(O12283));
  NOR2X1 G14503 (.A1(W4959), .A2(W2530), .ZN(W8519));
  NOR2X1 G14504 (.A1(W586), .A2(I1435), .ZN(W8518));
  NOR2X1 G14505 (.A1(W39765), .A2(W28518), .ZN(O12284));
  NOR2X1 G14506 (.A1(W26790), .A2(W1521), .ZN(O12285));
  NOR2X1 G14507 (.A1(W570), .A2(W4276), .ZN(W8515));
  NOR2X1 G14508 (.A1(I32), .A2(I1045), .ZN(W8514));
  NOR2X1 G14509 (.A1(I1749), .A2(I604), .ZN(W8513));
  NOR2X1 G14510 (.A1(I163), .A2(W20852), .ZN(W22472));
  NOR2X1 G14511 (.A1(W20963), .A2(W22133), .ZN(W42372));
  NOR2X1 G14512 (.A1(W2728), .A2(W4051), .ZN(W8510));
  NOR2X1 G14513 (.A1(W36900), .A2(W18372), .ZN(O12287));
  NOR2X1 G14514 (.A1(W5364), .A2(W31976), .ZN(O12288));
  NOR2X1 G14515 (.A1(W27869), .A2(W9460), .ZN(W28251));
  NOR2X1 G14516 (.A1(W13910), .A2(W17655), .ZN(O4417));
  NOR2X1 G14517 (.A1(I1159), .A2(I1118), .ZN(O4416));
  NOR2X1 G14518 (.A1(W2807), .A2(W6598), .ZN(W22456));
  NOR2X1 G14519 (.A1(W1653), .A2(W8257), .ZN(W8613));
  NOR2X1 G14520 (.A1(I1844), .A2(I492), .ZN(W8612));
  NOR2X1 G14521 (.A1(I1834), .A2(W20471), .ZN(W22453));
  NOR2X1 G14522 (.A1(W16787), .A2(W38078), .ZN(O12229));
  NOR2X1 G14523 (.A1(W3680), .A2(W8208), .ZN(W8609));
  NOR2X1 G14524 (.A1(W2320), .A2(W11565), .ZN(O12230));
  NOR2X1 G14525 (.A1(W12648), .A2(W18159), .ZN(O4424));
  NOR2X1 G14526 (.A1(W10595), .A2(W13339), .ZN(O12233));
  NOR2X1 G14527 (.A1(W29455), .A2(W19504), .ZN(O12227));
  NOR2X1 G14528 (.A1(W5207), .A2(W6446), .ZN(W8603));
  NOR2X1 G14529 (.A1(W5383), .A2(W6157), .ZN(W8602));
  NOR2X1 G14530 (.A1(W1089), .A2(W5186), .ZN(W8601));
  NOR2X1 G14531 (.A1(W34013), .A2(W22619), .ZN(O12236));
  NOR2X1 G14532 (.A1(I936), .A2(W3482), .ZN(W8599));
  NOR2X1 G14533 (.A1(W983), .A2(W26754), .ZN(W28270));
  NOR2X1 G14534 (.A1(W3652), .A2(I1950), .ZN(W8597));
  NOR2X1 G14535 (.A1(W4421), .A2(W5702), .ZN(W8625));
  NOR2X1 G14536 (.A1(W29892), .A2(W3250), .ZN(O12212));
  NOR2X1 G14537 (.A1(W31629), .A2(W11164), .ZN(O12215));
  NOR2X1 G14538 (.A1(W1969), .A2(I1110), .ZN(W8631));
  NOR2X1 G14539 (.A1(I297), .A2(W5294), .ZN(O239));
  NOR2X1 G14540 (.A1(W887), .A2(W13513), .ZN(W22446));
  NOR2X1 G14541 (.A1(W6135), .A2(W7769), .ZN(W8628));
  NOR2X1 G14542 (.A1(W40160), .A2(W23975), .ZN(W42267));
  NOR2X1 G14543 (.A1(W2953), .A2(W1570), .ZN(W8626));
  NOR2X1 G14544 (.A1(W335), .A2(I1474), .ZN(W8596));
  NOR2X1 G14545 (.A1(W10745), .A2(W12947), .ZN(O12219));
  NOR2X1 G14546 (.A1(W16048), .A2(W3213), .ZN(O4426));
  NOR2X1 G14547 (.A1(W37210), .A2(W41182), .ZN(W42274));
  NOR2X1 G14548 (.A1(W18719), .A2(W3858), .ZN(W22450));
  NOR2X1 G14549 (.A1(W121), .A2(W2418), .ZN(W8618));
  NOR2X1 G14550 (.A1(W1835), .A2(W12000), .ZN(W22451));
  NOR2X1 G14551 (.A1(I1052), .A2(W1786), .ZN(W8615));
  NOR2X1 G14552 (.A1(W5497), .A2(I1514), .ZN(W8567));
  NOR2X1 G14553 (.A1(W32495), .A2(W28092), .ZN(O12248));
  NOR2X1 G14554 (.A1(W14969), .A2(W3967), .ZN(O12249));
  NOR2X1 G14555 (.A1(W647), .A2(I934), .ZN(W8576));
  NOR2X1 G14556 (.A1(I1648), .A2(I1638), .ZN(W8573));
  NOR2X1 G14557 (.A1(W13164), .A2(W19895), .ZN(O12257));
  NOR2X1 G14558 (.A1(W1633), .A2(I292), .ZN(W8571));
  NOR2X1 G14559 (.A1(W12928), .A2(W22177), .ZN(W42324));
  NOR2X1 G14560 (.A1(W3537), .A2(W4313), .ZN(W8568));
  NOR2X1 G14561 (.A1(I1718), .A2(I310), .ZN(W8579));
  NOR2X1 G14562 (.A1(W1520), .A2(W8238), .ZN(W8566));
  NOR2X1 G14563 (.A1(W5659), .A2(W1434), .ZN(O236));
  NOR2X1 G14564 (.A1(W41506), .A2(W4267), .ZN(O12264));
  NOR2X1 G14565 (.A1(W18622), .A2(W33435), .ZN(O12265));
  NOR2X1 G14566 (.A1(W12743), .A2(W32405), .ZN(W42334));
  NOR2X1 G14567 (.A1(W1410), .A2(I194), .ZN(W8560));
  NOR2X1 G14568 (.A1(W11566), .A2(W14067), .ZN(W22471));
  NOR2X1 G14569 (.A1(W23072), .A2(W16706), .ZN(O12310));
  NOR2X1 G14570 (.A1(W536), .A2(W3942), .ZN(W8580));
  NOR2X1 G14571 (.A1(W1301), .A2(W5489), .ZN(W8581));
  NOR2X1 G14572 (.A1(I850), .A2(W7830), .ZN(W8582));
  NOR2X1 G14573 (.A1(W3554), .A2(W2774), .ZN(W8583));
  NOR2X1 G14574 (.A1(I1701), .A2(W5206), .ZN(W8585));
  NOR2X1 G14575 (.A1(W6253), .A2(W228), .ZN(W22464));
  NOR2X1 G14576 (.A1(W17526), .A2(W4794), .ZN(W22463));
  NOR2X1 G14577 (.A1(W17307), .A2(W17926), .ZN(O12244));
  NOR2X1 G14578 (.A1(W1705), .A2(W3802), .ZN(W8589));
  NOR2X1 G14579 (.A1(W24636), .A2(W687), .ZN(W28268));
  NOR2X1 G14580 (.A1(W22908), .A2(W1532), .ZN(O4422));
  NOR2X1 G14581 (.A1(W7033), .A2(W21800), .ZN(O2519));
  NOR2X1 G14582 (.A1(W28007), .A2(W40950), .ZN(W42299));
  NOR2X1 G14583 (.A1(I543), .A2(I532), .ZN(W22459));
  NOR2X1 G14584 (.A1(W2195), .A2(W13098), .ZN(W22458));
  NOR2X1 G14585 (.A1(W33278), .A2(W1144), .ZN(O12405));
  NOR2X1 G14586 (.A1(W23189), .A2(W18692), .ZN(W42499));
  NOR2X1 G14587 (.A1(W33215), .A2(W37822), .ZN(O12394));
  NOR2X1 G14588 (.A1(W19209), .A2(W19625), .ZN(O12396));
  NOR2X1 G14589 (.A1(W34796), .A2(W28484), .ZN(O12399));
  NOR2X1 G14590 (.A1(W18263), .A2(W24882), .ZN(W42510));
  NOR2X1 G14591 (.A1(W2264), .A2(W10233), .ZN(O4405));
  NOR2X1 G14592 (.A1(W7761), .A2(W5291), .ZN(W8386));
  NOR2X1 G14593 (.A1(I1419), .A2(W1643), .ZN(W8385));
  NOR2X1 G14594 (.A1(W14392), .A2(W12513), .ZN(O12392));
  NOR2X1 G14595 (.A1(W16858), .A2(W39426), .ZN(O12406));
  NOR2X1 G14596 (.A1(W7487), .A2(W6384), .ZN(W8381));
  NOR2X1 G14597 (.A1(W26844), .A2(W29550), .ZN(O12408));
  NOR2X1 G14598 (.A1(W5181), .A2(W4754), .ZN(W8379));
  NOR2X1 G14599 (.A1(I502), .A2(W8165), .ZN(O225));
  NOR2X1 G14600 (.A1(W3486), .A2(W20784), .ZN(W22523));
  NOR2X1 G14601 (.A1(W23048), .A2(W19722), .ZN(W42522));
  NOR2X1 G14602 (.A1(W4777), .A2(W294), .ZN(W8403));
  NOR2X1 G14603 (.A1(W2363), .A2(W8029), .ZN(W8412));
  NOR2X1 G14604 (.A1(W27056), .A2(W17265), .ZN(O4408));
  NOR2X1 G14605 (.A1(W20551), .A2(I1150), .ZN(O12380));
  NOR2X1 G14606 (.A1(W2161), .A2(W6855), .ZN(W8409));
  NOR2X1 G14607 (.A1(W1103), .A2(I524), .ZN(W8407));
  NOR2X1 G14608 (.A1(W4968), .A2(I665), .ZN(W8406));
  NOR2X1 G14609 (.A1(W4436), .A2(W2202), .ZN(W8405));
  NOR2X1 G14610 (.A1(W7166), .A2(W17771), .ZN(O4407));
  NOR2X1 G14611 (.A1(W5458), .A2(W3644), .ZN(W8375));
  NOR2X1 G14612 (.A1(W490), .A2(I1054), .ZN(W8402));
  NOR2X1 G14613 (.A1(W1336), .A2(W15672), .ZN(W22517));
  NOR2X1 G14614 (.A1(W6370), .A2(W1181), .ZN(O12386));
  NOR2X1 G14615 (.A1(W39948), .A2(W5861), .ZN(O12387));
  NOR2X1 G14616 (.A1(W16630), .A2(W41363), .ZN(O12390));
  NOR2X1 G14617 (.A1(W1061), .A2(W12599), .ZN(W22518));
  NOR2X1 G14618 (.A1(W4803), .A2(I1478), .ZN(W8396));
  NOR2X1 G14619 (.A1(W31763), .A2(W39581), .ZN(O12427));
  NOR2X1 G14620 (.A1(W1889), .A2(I557), .ZN(W8356));
  NOR2X1 G14621 (.A1(I109), .A2(W5513), .ZN(W8355));
  NOR2X1 G14622 (.A1(W1655), .A2(W3777), .ZN(W8354));
  NOR2X1 G14623 (.A1(W5263), .A2(W4993), .ZN(W8353));
  NOR2X1 G14624 (.A1(W5284), .A2(W12609), .ZN(W22530));
  NOR2X1 G14625 (.A1(I796), .A2(I1616), .ZN(W8351));
  NOR2X1 G14626 (.A1(W20960), .A2(W101), .ZN(O4403));
  NOR2X1 G14627 (.A1(W22944), .A2(W777), .ZN(O12425));
  NOR2X1 G14628 (.A1(W18955), .A2(W18466), .ZN(W22529));
  NOR2X1 G14629 (.A1(W1634), .A2(W5019), .ZN(W8347));
  NOR2X1 G14630 (.A1(W3812), .A2(W955), .ZN(W8345));
  NOR2X1 G14631 (.A1(I90), .A2(W17978), .ZN(W42552));
  NOR2X1 G14632 (.A1(I1508), .A2(W1619), .ZN(W8343));
  NOR2X1 G14633 (.A1(W7900), .A2(W2374), .ZN(O224));
  NOR2X1 G14634 (.A1(W7839), .A2(W7210), .ZN(W8341));
  NOR2X1 G14635 (.A1(W8003), .A2(I48), .ZN(W8340));
  NOR2X1 G14636 (.A1(W38123), .A2(W14379), .ZN(O12416));
  NOR2X1 G14637 (.A1(W6075), .A2(W6330), .ZN(W22524));
  NOR2X1 G14638 (.A1(W35793), .A2(W7416), .ZN(O12410));
  NOR2X1 G14639 (.A1(W3860), .A2(I1436), .ZN(W8372));
  NOR2X1 G14640 (.A1(W2561), .A2(W3226), .ZN(W8371));
  NOR2X1 G14641 (.A1(W31375), .A2(W5573), .ZN(O12411));
  NOR2X1 G14642 (.A1(W2050), .A2(W5126), .ZN(W8368));
  NOR2X1 G14643 (.A1(I1917), .A2(I764), .ZN(W22526));
  NOR2X1 G14644 (.A1(W14160), .A2(W7815), .ZN(O12415));
  NOR2X1 G14645 (.A1(W9322), .A2(W10572), .ZN(W22513));
  NOR2X1 G14646 (.A1(W889), .A2(W33605), .ZN(W42534));
  NOR2X1 G14647 (.A1(W6663), .A2(W7469), .ZN(W8363));
  NOR2X1 G14648 (.A1(W7391), .A2(W3847), .ZN(W8362));
  NOR2X1 G14649 (.A1(I115), .A2(W28886), .ZN(W42536));
  NOR2X1 G14650 (.A1(W16515), .A2(W12915), .ZN(W22527));
  NOR2X1 G14651 (.A1(W3319), .A2(W14595), .ZN(O2542));
  NOR2X1 G14652 (.A1(W4293), .A2(W455), .ZN(W8358));
  NOR2X1 G14653 (.A1(W7530), .A2(W447), .ZN(W42423));
  NOR2X1 G14654 (.A1(W15858), .A2(W27396), .ZN(O12324));
  NOR2X1 G14655 (.A1(W18049), .A2(W5817), .ZN(O2533));
  NOR2X1 G14656 (.A1(W3321), .A2(W7122), .ZN(O4412));
  NOR2X1 G14657 (.A1(W2080), .A2(W7737), .ZN(O230));
  NOR2X1 G14658 (.A1(W8016), .A2(W4108), .ZN(W8462));
  NOR2X1 G14659 (.A1(W4201), .A2(W27383), .ZN(W42421));
  NOR2X1 G14660 (.A1(W21791), .A2(I182), .ZN(O12329));
  NOR2X1 G14661 (.A1(W1694), .A2(W2282), .ZN(W8459));
  NOR2X1 G14662 (.A1(W16360), .A2(W11048), .ZN(O2532));
  NOR2X1 G14663 (.A1(W6560), .A2(W24719), .ZN(O12330));
  NOR2X1 G14664 (.A1(W1125), .A2(I289), .ZN(W8456));
  NOR2X1 G14665 (.A1(W7034), .A2(W1203), .ZN(W8455));
  NOR2X1 G14666 (.A1(I198), .A2(W31423), .ZN(O12334));
  NOR2X1 G14667 (.A1(W38961), .A2(W22723), .ZN(O12335));
  NOR2X1 G14668 (.A1(I547), .A2(W17342), .ZN(W42430));
  NOR2X1 G14669 (.A1(W18041), .A2(W23064), .ZN(W42432));
  NOR2X1 G14670 (.A1(W108), .A2(W27815), .ZN(O12319));
  NOR2X1 G14671 (.A1(W7118), .A2(W840), .ZN(W8483));
  NOR2X1 G14672 (.A1(W28019), .A2(W39281), .ZN(O12312));
  NOR2X1 G14673 (.A1(I304), .A2(W8748), .ZN(O12313));
  NOR2X1 G14674 (.A1(W1081), .A2(I350), .ZN(W8480));
  NOR2X1 G14675 (.A1(I114), .A2(W7023), .ZN(W8479));
  NOR2X1 G14676 (.A1(I1953), .A2(W1757), .ZN(O12314));
  NOR2X1 G14677 (.A1(W3190), .A2(W6666), .ZN(W8477));
  NOR2X1 G14678 (.A1(W24178), .A2(W23880), .ZN(W28239));
  NOR2X1 G14679 (.A1(I110), .A2(W8425), .ZN(W8449));
  NOR2X1 G14680 (.A1(W7759), .A2(W9327), .ZN(O12320));
  NOR2X1 G14681 (.A1(I980), .A2(I435), .ZN(W8473));
  NOR2X1 G14682 (.A1(W21025), .A2(W9061), .ZN(W22495));
  NOR2X1 G14683 (.A1(W18683), .A2(W8373), .ZN(O4413));
  NOR2X1 G14684 (.A1(W4610), .A2(I1310), .ZN(W8470));
  NOR2X1 G14685 (.A1(W2013), .A2(W7015), .ZN(W8469));
  NOR2X1 G14686 (.A1(W1267), .A2(W7373), .ZN(W8468));
  NOR2X1 G14687 (.A1(W4511), .A2(W3209), .ZN(W8421));
  NOR2X1 G14688 (.A1(W41712), .A2(W26137), .ZN(O12353));
  NOR2X1 G14689 (.A1(W11196), .A2(W37434), .ZN(O12354));
  NOR2X1 G14690 (.A1(I927), .A2(I1520), .ZN(W8428));
  NOR2X1 G14691 (.A1(I1152), .A2(W7237), .ZN(W8427));
  NOR2X1 G14692 (.A1(W660), .A2(W3697), .ZN(W8426));
  NOR2X1 G14693 (.A1(W14777), .A2(W16627), .ZN(W22510));
  NOR2X1 G14694 (.A1(W10245), .A2(W7779), .ZN(W22511));
  NOR2X1 G14695 (.A1(W1585), .A2(W4541), .ZN(W8423));
  NOR2X1 G14696 (.A1(W8648), .A2(W18436), .ZN(W22509));
  NOR2X1 G14697 (.A1(W17109), .A2(W22330), .ZN(O12363));
  NOR2X1 G14698 (.A1(W6032), .A2(W19494), .ZN(O12364));
  NOR2X1 G14699 (.A1(W31763), .A2(W15398), .ZN(O12365));
  NOR2X1 G14700 (.A1(W41704), .A2(W2728), .ZN(O12366));
  NOR2X1 G14701 (.A1(W33722), .A2(W30142), .ZN(O12367));
  NOR2X1 G14702 (.A1(W41294), .A2(W2185), .ZN(O12369));
  NOR2X1 G14703 (.A1(W20009), .A2(W40757), .ZN(O12370));
  NOR2X1 G14704 (.A1(W6893), .A2(W39934), .ZN(O12211));
  NOR2X1 G14705 (.A1(W11227), .A2(W3073), .ZN(W22508));
  NOR2X1 G14706 (.A1(I393), .A2(W25272), .ZN(O12351));
  NOR2X1 G14707 (.A1(W1529), .A2(I1689), .ZN(W8434));
  NOR2X1 G14708 (.A1(W2219), .A2(W1220), .ZN(W8435));
  NOR2X1 G14709 (.A1(W34373), .A2(W7409), .ZN(O12350));
  NOR2X1 G14710 (.A1(W40675), .A2(W41125), .ZN(O12346));
  NOR2X1 G14711 (.A1(W891), .A2(W3707), .ZN(W8439));
  NOR2X1 G14712 (.A1(W12679), .A2(W2183), .ZN(W22506));
  NOR2X1 G14713 (.A1(W2429), .A2(W5664), .ZN(W8441));
  NOR2X1 G14714 (.A1(W23619), .A2(W12332), .ZN(W28231));
  NOR2X1 G14715 (.A1(W3534), .A2(W6749), .ZN(O2537));
  NOR2X1 G14716 (.A1(W1456), .A2(I243), .ZN(W22503));
  NOR2X1 G14717 (.A1(W14543), .A2(W2801), .ZN(O2536));
  NOR2X1 G14718 (.A1(W5889), .A2(W23950), .ZN(O12340));
  NOR2X1 G14719 (.A1(W23695), .A2(W34326), .ZN(O12339));
  NOR2X1 G14720 (.A1(I228), .A2(W4190), .ZN(W8838));
  NOR2X1 G14721 (.A1(W4444), .A2(W5920), .ZN(O12064));
  NOR2X1 G14722 (.A1(W8199), .A2(W18330), .ZN(O12065));
  NOR2X1 G14723 (.A1(W41236), .A2(W30765), .ZN(O12066));
  NOR2X1 G14724 (.A1(W3114), .A2(W2361), .ZN(W8845));
  NOR2X1 G14725 (.A1(W1391), .A2(W6603), .ZN(W8842));
  NOR2X1 G14726 (.A1(W6757), .A2(W6382), .ZN(O250));
  NOR2X1 G14727 (.A1(W9637), .A2(W26851), .ZN(W42074));
  NOR2X1 G14728 (.A1(W4220), .A2(W6340), .ZN(W8839));
  NOR2X1 G14729 (.A1(W5883), .A2(W3637), .ZN(W8850));
  NOR2X1 G14730 (.A1(W58), .A2(I1876), .ZN(W8837));
  NOR2X1 G14731 (.A1(W6194), .A2(W9011), .ZN(W28373));
  NOR2X1 G14732 (.A1(W13470), .A2(W10305), .ZN(O12073));
  NOR2X1 G14733 (.A1(W28472), .A2(W41650), .ZN(O12074));
  NOR2X1 G14734 (.A1(W274), .A2(W24319), .ZN(O12075));
  NOR2X1 G14735 (.A1(W1270), .A2(W23242), .ZN(O12077));
  NOR2X1 G14736 (.A1(W2903), .A2(W5773), .ZN(O12078));
  NOR2X1 G14737 (.A1(W5311), .A2(W4434), .ZN(W8858));
  NOR2X1 G14738 (.A1(W8764), .A2(W9112), .ZN(W22366));
  NOR2X1 G14739 (.A1(W25099), .A2(W28708), .ZN(O12048));
  NOR2X1 G14740 (.A1(W16378), .A2(W18775), .ZN(W28387));
  NOR2X1 G14741 (.A1(W5330), .A2(W8619), .ZN(W8864));
  NOR2X1 G14742 (.A1(W16785), .A2(W10531), .ZN(O12050));
  NOR2X1 G14743 (.A1(W26556), .A2(W27766), .ZN(O12051));
  NOR2X1 G14744 (.A1(W17291), .A2(W22357), .ZN(W22369));
  NOR2X1 G14745 (.A1(W5358), .A2(W600), .ZN(W8859));
  NOR2X1 G14746 (.A1(W1543), .A2(I233), .ZN(O248));
  NOR2X1 G14747 (.A1(W6544), .A2(W7648), .ZN(W8857));
  NOR2X1 G14748 (.A1(W9092), .A2(I1956), .ZN(W22370));
  NOR2X1 G14749 (.A1(W5353), .A2(W16478), .ZN(W42056));
  NOR2X1 G14750 (.A1(I259), .A2(W18572), .ZN(W42058));
  NOR2X1 G14751 (.A1(W18460), .A2(W2119), .ZN(O12058));
  NOR2X1 G14752 (.A1(W18359), .A2(W23704), .ZN(O4474));
  NOR2X1 G14753 (.A1(W33213), .A2(W39157), .ZN(O12063));
  NOR2X1 G14754 (.A1(W8379), .A2(W4009), .ZN(O12096));
  NOR2X1 G14755 (.A1(I438), .A2(I1008), .ZN(W8808));
  NOR2X1 G14756 (.A1(W13516), .A2(W7107), .ZN(O12092));
  NOR2X1 G14757 (.A1(W19891), .A2(W2469), .ZN(O12093));
  NOR2X1 G14758 (.A1(I1714), .A2(W3465), .ZN(O4467));
  NOR2X1 G14759 (.A1(W4509), .A2(W1145), .ZN(W8803));
  NOR2X1 G14760 (.A1(W27198), .A2(W36433), .ZN(W42107));
  NOR2X1 G14761 (.A1(W9361), .A2(W9869), .ZN(W28360));
  NOR2X1 G14762 (.A1(I538), .A2(W20488), .ZN(W42109));
  NOR2X1 G14763 (.A1(W7091), .A2(W2450), .ZN(W8809));
  NOR2X1 G14764 (.A1(W1717), .A2(W6574), .ZN(O2495));
  NOR2X1 G14765 (.A1(W4301), .A2(W1140), .ZN(W8797));
  NOR2X1 G14766 (.A1(W13300), .A2(W11007), .ZN(W28359));
  NOR2X1 G14767 (.A1(W13851), .A2(W10154), .ZN(O12101));
  NOR2X1 G14768 (.A1(W6645), .A2(I1033), .ZN(W8794));
  NOR2X1 G14769 (.A1(W4811), .A2(W2398), .ZN(W8793));
  NOR2X1 G14770 (.A1(W22624), .A2(W13061), .ZN(W28358));
  NOR2X1 G14771 (.A1(W24872), .A2(W198), .ZN(W42092));
  NOR2X1 G14772 (.A1(W38959), .A2(W41575), .ZN(O12079));
  NOR2X1 G14773 (.A1(W6839), .A2(W6861), .ZN(W8827));
  NOR2X1 G14774 (.A1(W8273), .A2(W3960), .ZN(W8826));
  NOR2X1 G14775 (.A1(W126), .A2(W986), .ZN(W8824));
  NOR2X1 G14776 (.A1(W3676), .A2(W8741), .ZN(W8822));
  NOR2X1 G14777 (.A1(W3068), .A2(I1844), .ZN(W8821));
  NOR2X1 G14778 (.A1(W4039), .A2(W15854), .ZN(W28369));
  NOR2X1 G14779 (.A1(W7710), .A2(I1822), .ZN(W8819));
  NOR2X1 G14780 (.A1(W17704), .A2(W29861), .ZN(O12046));
  NOR2X1 G14781 (.A1(W3209), .A2(I255), .ZN(W8817));
  NOR2X1 G14782 (.A1(W37951), .A2(W15086), .ZN(O12085));
  NOR2X1 G14783 (.A1(W356), .A2(W8545), .ZN(W28368));
  NOR2X1 G14784 (.A1(W6988), .A2(W34336), .ZN(O12089));
  NOR2X1 G14785 (.A1(W8085), .A2(W2284), .ZN(W42099));
  NOR2X1 G14786 (.A1(W2424), .A2(W983), .ZN(W8811));
  NOR2X1 G14787 (.A1(W25713), .A2(W2388), .ZN(O12090));
  NOR2X1 G14788 (.A1(W5866), .A2(W26720), .ZN(W28406));
  NOR2X1 G14789 (.A1(W4822), .A2(W26407), .ZN(W28411));
  NOR2X1 G14790 (.A1(W6174), .A2(W23877), .ZN(W28408));
  NOR2X1 G14791 (.A1(W8365), .A2(W1634), .ZN(O254));
  NOR2X1 G14792 (.A1(W8499), .A2(W1522), .ZN(W8922));
  NOR2X1 G14793 (.A1(W6975), .A2(W4380), .ZN(W8920));
  NOR2X1 G14794 (.A1(W35209), .A2(W35117), .ZN(W41988));
  NOR2X1 G14795 (.A1(W5414), .A2(W5401), .ZN(W8918));
  NOR2X1 G14796 (.A1(W7295), .A2(W6115), .ZN(W8917));
  NOR2X1 G14797 (.A1(W12348), .A2(W38949), .ZN(O11999));
  NOR2X1 G14798 (.A1(W2827), .A2(W2002), .ZN(W8915));
  NOR2X1 G14799 (.A1(W5976), .A2(W3663), .ZN(W8914));
  NOR2X1 G14800 (.A1(I1939), .A2(W2126), .ZN(W8913));
  NOR2X1 G14801 (.A1(W29442), .A2(W16804), .ZN(O12006));
  NOR2X1 G14802 (.A1(W186), .A2(W5481), .ZN(W8911));
  NOR2X1 G14803 (.A1(W21059), .A2(W19217), .ZN(O4485));
  NOR2X1 G14804 (.A1(W13665), .A2(W13981), .ZN(W22353));
  NOR2X1 G14805 (.A1(W377), .A2(W7300), .ZN(O257));
  NOR2X1 G14806 (.A1(W22), .A2(W18708), .ZN(O2483));
  NOR2X1 G14807 (.A1(W17331), .A2(W12177), .ZN(O4492));
  NOR2X1 G14808 (.A1(W18156), .A2(W17835), .ZN(O4491));
  NOR2X1 G14809 (.A1(W33803), .A2(W30479), .ZN(O11988));
  NOR2X1 G14810 (.A1(W30817), .A2(W37738), .ZN(O11989));
  NOR2X1 G14811 (.A1(W14601), .A2(I1724), .ZN(W22338));
  NOR2X1 G14812 (.A1(W25616), .A2(I1121), .ZN(O11991));
  NOR2X1 G14813 (.A1(W26691), .A2(W2190), .ZN(O11992));
  NOR2X1 G14814 (.A1(W22135), .A2(W19190), .ZN(W22354));
  NOR2X1 G14815 (.A1(W18568), .A2(W23918), .ZN(W28417));
  NOR2X1 G14816 (.A1(W35950), .A2(W17197), .ZN(O11995));
  NOR2X1 G14817 (.A1(W2141), .A2(W8375), .ZN(O255));
  NOR2X1 G14818 (.A1(W7363), .A2(I594), .ZN(W8932));
  NOR2X1 G14819 (.A1(W15567), .A2(W18901), .ZN(W28412));
  NOR2X1 G14820 (.A1(W27827), .A2(W40240), .ZN(O11997));
  NOR2X1 G14821 (.A1(W2044), .A2(W8644), .ZN(O2484));
  NOR2X1 G14822 (.A1(W3156), .A2(W4464), .ZN(W8878));
  NOR2X1 G14823 (.A1(W20296), .A2(I1546), .ZN(O12028));
  NOR2X1 G14824 (.A1(W263), .A2(W2090), .ZN(W8885));
  NOR2X1 G14825 (.A1(W6602), .A2(W2960), .ZN(W8884));
  NOR2X1 G14826 (.A1(I570), .A2(W39267), .ZN(O12029));
  NOR2X1 G14827 (.A1(W16333), .A2(W9195), .ZN(O12031));
  NOR2X1 G14828 (.A1(W10177), .A2(W22723), .ZN(O12036));
  NOR2X1 G14829 (.A1(W4963), .A2(W2809), .ZN(O252));
  NOR2X1 G14830 (.A1(W2756), .A2(W17784), .ZN(W22359));
  NOR2X1 G14831 (.A1(W6038), .A2(W6703), .ZN(W8887));
  NOR2X1 G14832 (.A1(W3611), .A2(W4367), .ZN(W8877));
  NOR2X1 G14833 (.A1(W9675), .A2(W16187), .ZN(W22360));
  NOR2X1 G14834 (.A1(W11979), .A2(W41620), .ZN(W42032));
  NOR2X1 G14835 (.A1(I1384), .A2(W4172), .ZN(W28392));
  NOR2X1 G14836 (.A1(W21069), .A2(I750), .ZN(O2489));
  NOR2X1 G14837 (.A1(W2722), .A2(W1742), .ZN(W8870));
  NOR2X1 G14838 (.A1(W3112), .A2(W19435), .ZN(W22365));
  NOR2X1 G14839 (.A1(W10078), .A2(W18656), .ZN(O12103));
  NOR2X1 G14840 (.A1(W697), .A2(W5070), .ZN(W8888));
  NOR2X1 G14841 (.A1(W30941), .A2(I62), .ZN(W42019));
  NOR2X1 G14842 (.A1(W2318), .A2(W1914), .ZN(W8890));
  NOR2X1 G14843 (.A1(W7035), .A2(W1321), .ZN(W8892));
  NOR2X1 G14844 (.A1(W22870), .A2(W28633), .ZN(O12025));
  NOR2X1 G14845 (.A1(W31563), .A2(W37825), .ZN(O12022));
  NOR2X1 G14846 (.A1(W4054), .A2(W7076), .ZN(W8895));
  NOR2X1 G14847 (.A1(W2133), .A2(W6263), .ZN(W8898));
  NOR2X1 G14848 (.A1(I1660), .A2(W6582), .ZN(O253));
  NOR2X1 G14849 (.A1(W29328), .A2(W17567), .ZN(O12017));
  NOR2X1 G14850 (.A1(W6221), .A2(W24723), .ZN(O12016));
  NOR2X1 G14851 (.A1(W5726), .A2(W35448), .ZN(O12015));
  NOR2X1 G14852 (.A1(W12466), .A2(W15944), .ZN(O12014));
  NOR2X1 G14853 (.A1(W41054), .A2(W22315), .ZN(W42003));
  NOR2X1 G14854 (.A1(W13011), .A2(W23709), .ZN(W28399));
  NOR2X1 G14855 (.A1(W27818), .A2(W26852), .ZN(W28307));
  NOR2X1 G14856 (.A1(W1587), .A2(W5035), .ZN(O241));
  NOR2X1 G14857 (.A1(W6340), .A2(W7957), .ZN(W8689));
  NOR2X1 G14858 (.A1(W7673), .A2(W2146), .ZN(W8688));
  NOR2X1 G14859 (.A1(W834), .A2(W1828), .ZN(W8687));
  NOR2X1 G14860 (.A1(W2709), .A2(W304), .ZN(W8686));
  NOR2X1 G14861 (.A1(W34974), .A2(W6241), .ZN(O12179));
  NOR2X1 G14862 (.A1(W11149), .A2(W4362), .ZN(W42221));
  NOR2X1 G14863 (.A1(W7816), .A2(W3596), .ZN(W8681));
  NOR2X1 G14864 (.A1(W5244), .A2(W3911), .ZN(W8691));
  NOR2X1 G14865 (.A1(W5491), .A2(W6065), .ZN(W8678));
  NOR2X1 G14866 (.A1(W15885), .A2(W3736), .ZN(O2511));
  NOR2X1 G14867 (.A1(W7006), .A2(W15995), .ZN(W28305));
  NOR2X1 G14868 (.A1(W7970), .A2(W23082), .ZN(W28302));
  NOR2X1 G14869 (.A1(W1183), .A2(W38205), .ZN(O12191));
  NOR2X1 G14870 (.A1(W7917), .A2(W38251), .ZN(O12192));
  NOR2X1 G14871 (.A1(W4293), .A2(W2155), .ZN(W8670));
  NOR2X1 G14872 (.A1(I55), .A2(W7634), .ZN(W8699));
  NOR2X1 G14873 (.A1(W36778), .A2(W27397), .ZN(W42200));
  NOR2X1 G14874 (.A1(W9505), .A2(W4975), .ZN(W22422));
  NOR2X1 G14875 (.A1(W137), .A2(W2275), .ZN(W8706));
  NOR2X1 G14876 (.A1(W3989), .A2(I158), .ZN(W8705));
  NOR2X1 G14877 (.A1(W10330), .A2(W7353), .ZN(W28313));
  NOR2X1 G14878 (.A1(W2028), .A2(W19902), .ZN(O12169));
  NOR2X1 G14879 (.A1(W1356), .A2(W288), .ZN(W8702));
  NOR2X1 G14880 (.A1(W4111), .A2(W3155), .ZN(W8701));
  NOR2X1 G14881 (.A1(W1293), .A2(W1499), .ZN(W8669));
  NOR2X1 G14882 (.A1(W4040), .A2(W7330), .ZN(W8698));
  NOR2X1 G14883 (.A1(W33395), .A2(W269), .ZN(O12173));
  NOR2X1 G14884 (.A1(W22040), .A2(I1945), .ZN(O12174));
  NOR2X1 G14885 (.A1(W18414), .A2(W17047), .ZN(O12177));
  NOR2X1 G14886 (.A1(W12796), .A2(W4949), .ZN(O12178));
  NOR2X1 G14887 (.A1(W1225), .A2(W315), .ZN(W8693));
  NOR2X1 G14888 (.A1(I1364), .A2(W6166), .ZN(W8692));
  NOR2X1 G14889 (.A1(W4216), .A2(W14102), .ZN(W22443));
  NOR2X1 G14890 (.A1(I1393), .A2(W1772), .ZN(O12201));
  NOR2X1 G14891 (.A1(I436), .A2(W11620), .ZN(O12202));
  NOR2X1 G14892 (.A1(W38191), .A2(W12676), .ZN(O12203));
  NOR2X1 G14893 (.A1(W15176), .A2(W2542), .ZN(W22440));
  NOR2X1 G14894 (.A1(W41568), .A2(W35597), .ZN(W42252));
  NOR2X1 G14895 (.A1(W5503), .A2(W4195), .ZN(W8645));
  NOR2X1 G14896 (.A1(I1545), .A2(W5403), .ZN(O2515));
  NOR2X1 G14897 (.A1(W18335), .A2(W23202), .ZN(W28281));
  NOR2X1 G14898 (.A1(I690), .A2(W14002), .ZN(W28286));
  NOR2X1 G14899 (.A1(W15016), .A2(W7543), .ZN(O12207));
  NOR2X1 G14900 (.A1(W1701), .A2(W8470), .ZN(W8640));
  NOR2X1 G14901 (.A1(W2246), .A2(W22170), .ZN(O2516));
  NOR2X1 G14902 (.A1(W24648), .A2(W7783), .ZN(W28279));
  NOR2X1 G14903 (.A1(W7455), .A2(W2215), .ZN(W8637));
  NOR2X1 G14904 (.A1(W1322), .A2(W7087), .ZN(W8636));
  NOR2X1 G14905 (.A1(W31416), .A2(W7276), .ZN(O12210));
  NOR2X1 G14906 (.A1(W5468), .A2(W2369), .ZN(O243));
  NOR2X1 G14907 (.A1(W7475), .A2(I1616), .ZN(W8652));
  NOR2X1 G14908 (.A1(W1935), .A2(W6969), .ZN(W8653));
  NOR2X1 G14909 (.A1(W2381), .A2(W7338), .ZN(W8654));
  NOR2X1 G14910 (.A1(W2695), .A2(W6949), .ZN(W8655));
  NOR2X1 G14911 (.A1(W22843), .A2(W26751), .ZN(O4432));
  NOR2X1 G14912 (.A1(W20906), .A2(W16307), .ZN(W22437));
  NOR2X1 G14913 (.A1(W348), .A2(W3138), .ZN(W8658));
  NOR2X1 G14914 (.A1(W7238), .A2(W24583), .ZN(O12197));
  NOR2X1 G14915 (.A1(W39157), .A2(W39871), .ZN(O12196));
  NOR2X1 G14916 (.A1(W6133), .A2(W5166), .ZN(W8662));
  NOR2X1 G14917 (.A1(W1524), .A2(W4119), .ZN(W8663));
  NOR2X1 G14918 (.A1(W23629), .A2(W14602), .ZN(O12195));
  NOR2X1 G14919 (.A1(I1835), .A2(W2447), .ZN(W8665));
  NOR2X1 G14920 (.A1(W22701), .A2(W1906), .ZN(O12194));
  NOR2X1 G14921 (.A1(W17167), .A2(W23623), .ZN(O4434));
  NOR2X1 G14922 (.A1(W5401), .A2(I814), .ZN(O245));
  NOR2X1 G14923 (.A1(W7146), .A2(I927), .ZN(W8766));
  NOR2X1 G14924 (.A1(W6646), .A2(W6077), .ZN(W8765));
  NOR2X1 G14925 (.A1(W10220), .A2(W23961), .ZN(W28335));
  NOR2X1 G14926 (.A1(I1726), .A2(W7300), .ZN(W8763));
  NOR2X1 G14927 (.A1(W41342), .A2(W17833), .ZN(O12125));
  NOR2X1 G14928 (.A1(W3429), .A2(W71), .ZN(W8761));
  NOR2X1 G14929 (.A1(W6868), .A2(W738), .ZN(W8760));
  NOR2X1 G14930 (.A1(W40308), .A2(W33068), .ZN(W42144));
  NOR2X1 G14931 (.A1(W5408), .A2(W6590), .ZN(W8767));
  NOR2X1 G14932 (.A1(W15371), .A2(W23313), .ZN(W42145));
  NOR2X1 G14933 (.A1(W6906), .A2(W2154), .ZN(W42146));
  NOR2X1 G14934 (.A1(W2278), .A2(W3770), .ZN(W8755));
  NOR2X1 G14935 (.A1(W24393), .A2(W18711), .ZN(O12129));
  NOR2X1 G14936 (.A1(W29267), .A2(W22330), .ZN(O12130));
  NOR2X1 G14937 (.A1(W3712), .A2(W2813), .ZN(W8752));
  NOR2X1 G14938 (.A1(W5912), .A2(W18754), .ZN(W28331));
  NOR2X1 G14939 (.A1(W8677), .A2(W6146), .ZN(O4462));
  NOR2X1 G14940 (.A1(I1732), .A2(W19435), .ZN(W22388));
  NOR2X1 G14941 (.A1(W8467), .A2(W477), .ZN(O4464));
  NOR2X1 G14942 (.A1(W11533), .A2(W31957), .ZN(W42122));
  NOR2X1 G14943 (.A1(I66), .A2(W8681), .ZN(W8787));
  NOR2X1 G14944 (.A1(W21173), .A2(W19989), .ZN(W22390));
  NOR2X1 G14945 (.A1(W18701), .A2(W12928), .ZN(O4463));
  NOR2X1 G14946 (.A1(W7490), .A2(W4675), .ZN(W8784));
  NOR2X1 G14947 (.A1(W8657), .A2(I1393), .ZN(W8783));
  NOR2X1 G14948 (.A1(W8084), .A2(W10075), .ZN(W28328));
  NOR2X1 G14949 (.A1(W10152), .A2(W1508), .ZN(O12111));
  NOR2X1 G14950 (.A1(W1233), .A2(W9477), .ZN(W28345));
  NOR2X1 G14951 (.A1(W8694), .A2(W3149), .ZN(W8776));
  NOR2X1 G14952 (.A1(W624), .A2(W37028), .ZN(O12117));
  NOR2X1 G14953 (.A1(I1955), .A2(I495), .ZN(W8771));
  NOR2X1 G14954 (.A1(W8846), .A2(W14458), .ZN(W28336));
  NOR2X1 G14955 (.A1(W15919), .A2(W10862), .ZN(W22402));
  NOR2X1 G14956 (.A1(W21482), .A2(W12181), .ZN(W22419));
  NOR2X1 G14957 (.A1(W7458), .A2(W12108), .ZN(O12151));
  NOR2X1 G14958 (.A1(W8447), .A2(W7485), .ZN(W8728));
  NOR2X1 G14959 (.A1(I360), .A2(W5413), .ZN(W8726));
  NOR2X1 G14960 (.A1(W4491), .A2(I1334), .ZN(W22415));
  NOR2X1 G14961 (.A1(W5487), .A2(W14012), .ZN(W42187));
  NOR2X1 G14962 (.A1(I821), .A2(W7654), .ZN(O4443));
  NOR2X1 G14963 (.A1(W2428), .A2(I1282), .ZN(W8721));
  NOR2X1 G14964 (.A1(W4034), .A2(W2572), .ZN(W22418));
  NOR2X1 G14965 (.A1(W21663), .A2(W2940), .ZN(O4445));
  NOR2X1 G14966 (.A1(W1460), .A2(W6206), .ZN(W8718));
  NOR2X1 G14967 (.A1(W4833), .A2(W6593), .ZN(W8717));
  NOR2X1 G14968 (.A1(W2166), .A2(W17166), .ZN(O12163));
  NOR2X1 G14969 (.A1(W4114), .A2(W314), .ZN(W8715));
  NOR2X1 G14970 (.A1(W1509), .A2(W5915), .ZN(W8714));
  NOR2X1 G14971 (.A1(W7097), .A2(W4653), .ZN(W8713));
  NOR2X1 G14972 (.A1(W40991), .A2(W17392), .ZN(O12164));
  NOR2X1 G14973 (.A1(W3891), .A2(W3733), .ZN(W8339));
  NOR2X1 G14974 (.A1(W2658), .A2(W4157), .ZN(W8731));
  NOR2X1 G14975 (.A1(W20275), .A2(W15806), .ZN(O12146));
  NOR2X1 G14976 (.A1(W8996), .A2(W22257), .ZN(W22411));
  NOR2X1 G14977 (.A1(W4534), .A2(W1964), .ZN(W22410));
  NOR2X1 G14978 (.A1(W7018), .A2(W5334), .ZN(W8736));
  NOR2X1 G14979 (.A1(W6004), .A2(W8435), .ZN(W8737));
  NOR2X1 G14980 (.A1(W14639), .A2(W535), .ZN(O12145));
  NOR2X1 G14981 (.A1(W4077), .A2(I1864), .ZN(W8739));
  NOR2X1 G14982 (.A1(W12404), .A2(W27452), .ZN(O12141));
  NOR2X1 G14983 (.A1(W39328), .A2(W1741), .ZN(O12140));
  NOR2X1 G14984 (.A1(W4517), .A2(W17055), .ZN(O12139));
  NOR2X1 G14985 (.A1(W17615), .A2(W31813), .ZN(O12137));
  NOR2X1 G14986 (.A1(W8526), .A2(W3799), .ZN(W8746));
  NOR2X1 G14987 (.A1(I219), .A2(W2361), .ZN(W8747));
  NOR2X1 G14988 (.A1(W3813), .A2(W11091), .ZN(W28327));
  NOR2X1 G14989 (.A1(I276), .A2(W20615), .ZN(O4332));
  NOR2X1 G14990 (.A1(W17355), .A2(W14257), .ZN(W22679));
  NOR2X1 G14991 (.A1(W6590), .A2(I113), .ZN(W7941));
  NOR2X1 G14992 (.A1(W13764), .A2(W2794), .ZN(W22680));
  NOR2X1 G14993 (.A1(W645), .A2(I943), .ZN(W7939));
  NOR2X1 G14994 (.A1(I1882), .A2(W7788), .ZN(W7938));
  NOR2X1 G14995 (.A1(W18459), .A2(W23511), .ZN(W42955));
  NOR2X1 G14996 (.A1(W2633), .A2(W20530), .ZN(O4333));
  NOR2X1 G14997 (.A1(W18136), .A2(W19805), .ZN(W28058));
  NOR2X1 G14998 (.A1(W7289), .A2(I1011), .ZN(W7943));
  NOR2X1 G14999 (.A1(W35131), .A2(W33893), .ZN(W42964));
  NOR2X1 G15000 (.A1(W911), .A2(W381), .ZN(W7930));
  NOR2X1 G15001 (.A1(I1653), .A2(W906), .ZN(W7929));
  NOR2X1 G15002 (.A1(W30534), .A2(W37262), .ZN(O12747));
  NOR2X1 G15003 (.A1(W5478), .A2(W2601), .ZN(W7927));
  NOR2X1 G15004 (.A1(W15073), .A2(W8998), .ZN(W42967));
  NOR2X1 G15005 (.A1(I1175), .A2(I894), .ZN(W7925));
  NOR2X1 G15006 (.A1(W7381), .A2(I1246), .ZN(W7951));
  NOR2X1 G15007 (.A1(W13248), .A2(W26278), .ZN(O12724));
  NOR2X1 G15008 (.A1(W4589), .A2(W7210), .ZN(W7960));
  NOR2X1 G15009 (.A1(I1455), .A2(W4112), .ZN(W7958));
  NOR2X1 G15010 (.A1(W6237), .A2(W19992), .ZN(O12726));
  NOR2X1 G15011 (.A1(W1877), .A2(W25889), .ZN(W28065));
  NOR2X1 G15012 (.A1(W17723), .A2(W22523), .ZN(O12731));
  NOR2X1 G15013 (.A1(W17318), .A2(W33785), .ZN(W42946));
  NOR2X1 G15014 (.A1(W18391), .A2(W12086), .ZN(O12732));
  NOR2X1 G15015 (.A1(W16766), .A2(W15217), .ZN(O12749));
  NOR2X1 G15016 (.A1(I1953), .A2(W6477), .ZN(W7950));
  NOR2X1 G15017 (.A1(W677), .A2(I206), .ZN(W7949));
  NOR2X1 G15018 (.A1(W1803), .A2(W4795), .ZN(W7948));
  NOR2X1 G15019 (.A1(I732), .A2(W3132), .ZN(W7947));
  NOR2X1 G15020 (.A1(W23277), .A2(W18927), .ZN(W28063));
  NOR2X1 G15021 (.A1(W1859), .A2(W6764), .ZN(W7945));
  NOR2X1 G15022 (.A1(W14267), .A2(W24234), .ZN(O12734));
  NOR2X1 G15023 (.A1(W3545), .A2(W7521), .ZN(W7897));
  NOR2X1 G15024 (.A1(I825), .A2(W14258), .ZN(W22691));
  NOR2X1 G15025 (.A1(W23337), .A2(W3998), .ZN(O12765));
  NOR2X1 G15026 (.A1(W19757), .A2(W13632), .ZN(O2583));
  NOR2X1 G15027 (.A1(I886), .A2(W7167), .ZN(W7902));
  NOR2X1 G15028 (.A1(W3946), .A2(W4368), .ZN(W7901));
  NOR2X1 G15029 (.A1(W23875), .A2(W25732), .ZN(W28049));
  NOR2X1 G15030 (.A1(W3946), .A2(W2654), .ZN(W7899));
  NOR2X1 G15031 (.A1(W20580), .A2(W12883), .ZN(W22694));
  NOR2X1 G15032 (.A1(W6262), .A2(W38475), .ZN(W42989));
  NOR2X1 G15033 (.A1(W9395), .A2(W3179), .ZN(O4326));
  NOR2X1 G15034 (.A1(I388), .A2(I1948), .ZN(W7895));
  NOR2X1 G15035 (.A1(W19290), .A2(W9829), .ZN(W22696));
  NOR2X1 G15036 (.A1(W2986), .A2(W3730), .ZN(W7893));
  NOR2X1 G15037 (.A1(W38962), .A2(W33009), .ZN(O12772));
  NOR2X1 G15038 (.A1(W2194), .A2(I1040), .ZN(W7891));
  NOR2X1 G15039 (.A1(W10191), .A2(W24723), .ZN(O12773));
  NOR2X1 G15040 (.A1(W4187), .A2(W22531), .ZN(W22687));
  NOR2X1 G15041 (.A1(I512), .A2(W10619), .ZN(W42972));
  NOR2X1 G15042 (.A1(I324), .A2(W2814), .ZN(W22686));
  NOR2X1 G15043 (.A1(I1282), .A2(W714), .ZN(W7921));
  NOR2X1 G15044 (.A1(W5787), .A2(I588), .ZN(W7920));
  NOR2X1 G15045 (.A1(I1819), .A2(W6308), .ZN(W7919));
  NOR2X1 G15046 (.A1(I1034), .A2(W4952), .ZN(W7918));
  NOR2X1 G15047 (.A1(W362), .A2(W5311), .ZN(W7917));
  NOR2X1 G15048 (.A1(W5557), .A2(W27567), .ZN(O12756));
  NOR2X1 G15049 (.A1(W5519), .A2(W4259), .ZN(W7962));
  NOR2X1 G15050 (.A1(W3792), .A2(W6480), .ZN(W7914));
  NOR2X1 G15051 (.A1(W24559), .A2(I885), .ZN(O12757));
  NOR2X1 G15052 (.A1(I153), .A2(I1005), .ZN(W28052));
  NOR2X1 G15053 (.A1(W22865), .A2(W3839), .ZN(W28050));
  NOR2X1 G15054 (.A1(W9519), .A2(W13212), .ZN(O12759));
  NOR2X1 G15055 (.A1(W6855), .A2(W5106), .ZN(O12760));
  NOR2X1 G15056 (.A1(W10282), .A2(W1997), .ZN(O12761));
  NOR2X1 G15057 (.A1(W21095), .A2(W17565), .ZN(O2570));
  NOR2X1 G15058 (.A1(I1163), .A2(W340), .ZN(W8018));
  NOR2X1 G15059 (.A1(W7609), .A2(W1523), .ZN(W8017));
  NOR2X1 G15060 (.A1(W2879), .A2(W9536), .ZN(O2567));
  NOR2X1 G15061 (.A1(W5060), .A2(W22860), .ZN(O12679));
  NOR2X1 G15062 (.A1(W2594), .A2(I1550), .ZN(W22651));
  NOR2X1 G15063 (.A1(W6243), .A2(W6379), .ZN(W8013));
  NOR2X1 G15064 (.A1(W130), .A2(I1492), .ZN(W8012));
  NOR2X1 G15065 (.A1(W19713), .A2(W28935), .ZN(O12681));
  NOR2X1 G15066 (.A1(W25569), .A2(W14551), .ZN(W42872));
  NOR2X1 G15067 (.A1(W13818), .A2(W2567), .ZN(W28082));
  NOR2X1 G15068 (.A1(W26540), .A2(W24941), .ZN(O4340));
  NOR2X1 G15069 (.A1(W1021), .A2(W31920), .ZN(O12690));
  NOR2X1 G15070 (.A1(W20475), .A2(W22545), .ZN(O2574));
  NOR2X1 G15071 (.A1(W39353), .A2(W41774), .ZN(O12691));
  NOR2X1 G15072 (.A1(W6047), .A2(W20486), .ZN(O2575));
  NOR2X1 G15073 (.A1(W10094), .A2(W7152), .ZN(W22663));
  NOR2X1 G15074 (.A1(W8472), .A2(W4803), .ZN(W28089));
  NOR2X1 G15075 (.A1(W11163), .A2(W5486), .ZN(W28090));
  NOR2X1 G15076 (.A1(I1038), .A2(W21638), .ZN(W22645));
  NOR2X1 G15077 (.A1(W7196), .A2(W3085), .ZN(W8033));
  NOR2X1 G15078 (.A1(W9063), .A2(W16393), .ZN(O2564));
  NOR2X1 G15079 (.A1(W21988), .A2(W16973), .ZN(W22647));
  NOR2X1 G15080 (.A1(W41675), .A2(W24193), .ZN(O12666));
  NOR2X1 G15081 (.A1(W26453), .A2(W14346), .ZN(O12669));
  NOR2X1 G15082 (.A1(W25465), .A2(W30892), .ZN(W42864));
  NOR2X1 G15083 (.A1(W2997), .A2(W1472), .ZN(W7996));
  NOR2X1 G15084 (.A1(W7938), .A2(W3058), .ZN(W8026));
  NOR2X1 G15085 (.A1(W3651), .A2(W37404), .ZN(O12671));
  NOR2X1 G15086 (.A1(W6410), .A2(W107), .ZN(W8024));
  NOR2X1 G15087 (.A1(W19627), .A2(W7492), .ZN(W28088));
  NOR2X1 G15088 (.A1(W26065), .A2(W21345), .ZN(O12675));
  NOR2X1 G15089 (.A1(W6480), .A2(W5758), .ZN(W8021));
  NOR2X1 G15090 (.A1(W3253), .A2(W832), .ZN(W8020));
  NOR2X1 G15091 (.A1(I238), .A2(W6586), .ZN(W7971));
  NOR2X1 G15092 (.A1(W18940), .A2(W2061), .ZN(O12704));
  NOR2X1 G15093 (.A1(W21235), .A2(W12791), .ZN(O12705));
  NOR2X1 G15094 (.A1(I732), .A2(W4070), .ZN(W7977));
  NOR2X1 G15095 (.A1(W31562), .A2(W30406), .ZN(O12707));
  NOR2X1 G15096 (.A1(W24831), .A2(W36284), .ZN(O12711));
  NOR2X1 G15097 (.A1(W1340), .A2(W1493), .ZN(O12712));
  NOR2X1 G15098 (.A1(W17669), .A2(W18482), .ZN(W28072));
  NOR2X1 G15099 (.A1(W16011), .A2(W18934), .ZN(O12714));
  NOR2X1 G15100 (.A1(W18003), .A2(W15728), .ZN(O2577));
  NOR2X1 G15101 (.A1(W5883), .A2(W19602), .ZN(W28071));
  NOR2X1 G15102 (.A1(W9991), .A2(W22263), .ZN(W42926));
  NOR2X1 G15103 (.A1(W40371), .A2(W4177), .ZN(W42927));
  NOR2X1 G15104 (.A1(W6102), .A2(W406), .ZN(W7967));
  NOR2X1 G15105 (.A1(W20805), .A2(W15378), .ZN(O2580));
  NOR2X1 G15106 (.A1(W15011), .A2(W9489), .ZN(W22673));
  NOR2X1 G15107 (.A1(W23211), .A2(W23630), .ZN(O12722));
  NOR2X1 G15108 (.A1(W2985), .A2(W3894), .ZN(W7889));
  NOR2X1 G15109 (.A1(W10704), .A2(W8929), .ZN(W22668));
  NOR2X1 G15110 (.A1(I306), .A2(W477), .ZN(W7982));
  NOR2X1 G15111 (.A1(W26017), .A2(W9615), .ZN(O12701));
  NOR2X1 G15112 (.A1(W8137), .A2(W20412), .ZN(W22667));
  NOR2X1 G15113 (.A1(W2827), .A2(W7705), .ZN(O207));
  NOR2X1 G15114 (.A1(W6414), .A2(W25003), .ZN(O12699));
  NOR2X1 G15115 (.A1(W6235), .A2(W4426), .ZN(O12698));
  NOR2X1 G15116 (.A1(W6229), .A2(W3493), .ZN(W7988));
  NOR2X1 G15117 (.A1(I978), .A2(W5218), .ZN(W22666));
  NOR2X1 G15118 (.A1(W112), .A2(I1431), .ZN(W28073));
  NOR2X1 G15119 (.A1(W1268), .A2(W8319), .ZN(W28076));
  NOR2X1 G15120 (.A1(W39028), .A2(W18669), .ZN(O12695));
  NOR2X1 G15121 (.A1(I1079), .A2(W7553), .ZN(W7993));
  NOR2X1 G15122 (.A1(W7876), .A2(W32), .ZN(W7994));
  NOR2X1 G15123 (.A1(W7749), .A2(W6662), .ZN(W7995));
  NOR2X1 G15124 (.A1(W18798), .A2(W39503), .ZN(O12853));
  NOR2X1 G15125 (.A1(W11973), .A2(W10908), .ZN(O4313));
  NOR2X1 G15126 (.A1(W33862), .A2(W24270), .ZN(W43093));
  NOR2X1 G15127 (.A1(W2911), .A2(W26529), .ZN(O12849));
  NOR2X1 G15128 (.A1(W31775), .A2(W12181), .ZN(O12850));
  NOR2X1 G15129 (.A1(W4216), .A2(W4884), .ZN(W7793));
  NOR2X1 G15130 (.A1(W12513), .A2(W28481), .ZN(O12852));
  NOR2X1 G15131 (.A1(W9750), .A2(W19926), .ZN(W22732));
  NOR2X1 G15132 (.A1(W3281), .A2(W416), .ZN(W7790));
  NOR2X1 G15133 (.A1(W26357), .A2(W8234), .ZN(W28018));
  NOR2X1 G15134 (.A1(W6364), .A2(W38076), .ZN(O12854));
  NOR2X1 G15135 (.A1(W2271), .A2(W474), .ZN(W7787));
  NOR2X1 G15136 (.A1(W3796), .A2(W20630), .ZN(W28016));
  NOR2X1 G15137 (.A1(W32949), .A2(W965), .ZN(W43104));
  NOR2X1 G15138 (.A1(W2312), .A2(W22721), .ZN(O2594));
  NOR2X1 G15139 (.A1(W5467), .A2(W973), .ZN(W7783));
  NOR2X1 G15140 (.A1(W2396), .A2(W15226), .ZN(W28012));
  NOR2X1 G15141 (.A1(W4077), .A2(W10945), .ZN(W22726));
  NOR2X1 G15142 (.A1(W8088), .A2(W2651), .ZN(O12829));
  NOR2X1 G15143 (.A1(W25119), .A2(W42731), .ZN(O12830));
  NOR2X1 G15144 (.A1(W20376), .A2(W1518), .ZN(O2592));
  NOR2X1 G15145 (.A1(W5374), .A2(I443), .ZN(W7814));
  NOR2X1 G15146 (.A1(W7685), .A2(W909), .ZN(W7813));
  NOR2X1 G15147 (.A1(W3630), .A2(W751), .ZN(O202));
  NOR2X1 G15148 (.A1(W19993), .A2(W22376), .ZN(O4318));
  NOR2X1 G15149 (.A1(I356), .A2(W15131), .ZN(O12835));
  NOR2X1 G15150 (.A1(I1234), .A2(W19121), .ZN(O12858));
  NOR2X1 G15151 (.A1(W33857), .A2(W11300), .ZN(W43081));
  NOR2X1 G15152 (.A1(W16837), .A2(I245), .ZN(W22727));
  NOR2X1 G15153 (.A1(W5365), .A2(W6298), .ZN(O12841));
  NOR2X1 G15154 (.A1(W2654), .A2(W7358), .ZN(W7802));
  NOR2X1 G15155 (.A1(W12552), .A2(W6520), .ZN(O12843));
  NOR2X1 G15156 (.A1(W44), .A2(W6371), .ZN(W7800));
  NOR2X1 G15157 (.A1(W2049), .A2(W2501), .ZN(O4316));
  NOR2X1 G15158 (.A1(W1089), .A2(W5635), .ZN(W7751));
  NOR2X1 G15159 (.A1(W15323), .A2(W28433), .ZN(O12874));
  NOR2X1 G15160 (.A1(W27934), .A2(W27631), .ZN(O12875));
  NOR2X1 G15161 (.A1(W24161), .A2(W43025), .ZN(W43135));
  NOR2X1 G15162 (.A1(I1004), .A2(W6673), .ZN(W7756));
  NOR2X1 G15163 (.A1(W20761), .A2(W26810), .ZN(W43137));
  NOR2X1 G15164 (.A1(W42358), .A2(W34921), .ZN(O12877));
  NOR2X1 G15165 (.A1(W6027), .A2(W6929), .ZN(W7753));
  NOR2X1 G15166 (.A1(W40484), .A2(W2869), .ZN(O12879));
  NOR2X1 G15167 (.A1(W12403), .A2(W17420), .ZN(W28003));
  NOR2X1 G15168 (.A1(W19792), .A2(W4112), .ZN(W22744));
  NOR2X1 G15169 (.A1(W7540), .A2(W956), .ZN(W7749));
  NOR2X1 G15170 (.A1(W18422), .A2(W5205), .ZN(W22745));
  NOR2X1 G15171 (.A1(W27842), .A2(W25463), .ZN(O12882));
  NOR2X1 G15172 (.A1(W3476), .A2(W6719), .ZN(W7745));
  NOR2X1 G15173 (.A1(W382), .A2(W20168), .ZN(O12883));
  NOR2X1 G15174 (.A1(I195), .A2(W78), .ZN(W7743));
  NOR2X1 G15175 (.A1(W2414), .A2(W5935), .ZN(W7818));
  NOR2X1 G15176 (.A1(W34417), .A2(W24814), .ZN(W43129));
  NOR2X1 G15177 (.A1(W22032), .A2(W26603), .ZN(O12870));
  NOR2X1 G15178 (.A1(W3908), .A2(W30540), .ZN(O12868));
  NOR2X1 G15179 (.A1(W6314), .A2(W5401), .ZN(W7767));
  NOR2X1 G15180 (.A1(I797), .A2(W3713), .ZN(W7769));
  NOR2X1 G15181 (.A1(I31), .A2(W4041), .ZN(W7770));
  NOR2X1 G15182 (.A1(W16448), .A2(W15073), .ZN(W22738));
  NOR2X1 G15183 (.A1(W12213), .A2(W15447), .ZN(O12864));
  NOR2X1 G15184 (.A1(W7337), .A2(W7682), .ZN(W7773));
  NOR2X1 G15185 (.A1(I622), .A2(W6533), .ZN(W7774));
  NOR2X1 G15186 (.A1(W3922), .A2(W6383), .ZN(W7775));
  NOR2X1 G15187 (.A1(W22042), .A2(W17157), .ZN(W28011));
  NOR2X1 G15188 (.A1(I382), .A2(W3175), .ZN(W7777));
  NOR2X1 G15189 (.A1(W40486), .A2(W37610), .ZN(O12861));
  NOR2X1 G15190 (.A1(W1074), .A2(W715), .ZN(W7779));
  NOR2X1 G15191 (.A1(W973), .A2(W1418), .ZN(W7863));
  NOR2X1 G15192 (.A1(W25556), .A2(W7213), .ZN(W28044));
  NOR2X1 G15193 (.A1(W31247), .A2(W17325), .ZN(O12784));
  NOR2X1 G15194 (.A1(W19990), .A2(W21021), .ZN(W28041));
  NOR2X1 G15195 (.A1(W5403), .A2(W4046), .ZN(W7868));
  NOR2X1 G15196 (.A1(W14961), .A2(W26358), .ZN(W28038));
  NOR2X1 G15197 (.A1(W16743), .A2(W6542), .ZN(W22704));
  NOR2X1 G15198 (.A1(I415), .A2(W307), .ZN(W7865));
  NOR2X1 G15199 (.A1(W39061), .A2(W31773), .ZN(O12787));
  NOR2X1 G15200 (.A1(W23136), .A2(W27607), .ZN(O12782));
  NOR2X1 G15201 (.A1(W9025), .A2(W6851), .ZN(W22705));
  NOR2X1 G15202 (.A1(W5266), .A2(I1366), .ZN(W7861));
  NOR2X1 G15203 (.A1(W972), .A2(W6915), .ZN(W7860));
  NOR2X1 G15204 (.A1(W19010), .A2(W22399), .ZN(W28037));
  NOR2X1 G15205 (.A1(W3196), .A2(W7122), .ZN(O12789));
  NOR2X1 G15206 (.A1(W2208), .A2(W2241), .ZN(W7857));
  NOR2X1 G15207 (.A1(W16500), .A2(W27150), .ZN(O12790));
  NOR2X1 G15208 (.A1(W26836), .A2(W2482), .ZN(O12776));
  NOR2X1 G15209 (.A1(W37803), .A2(W14674), .ZN(W43002));
  NOR2X1 G15210 (.A1(W4890), .A2(W14202), .ZN(W43003));
  NOR2X1 G15211 (.A1(I296), .A2(W4237), .ZN(W7886));
  NOR2X1 G15212 (.A1(W6201), .A2(W3313), .ZN(W7885));
  NOR2X1 G15213 (.A1(W29315), .A2(W34791), .ZN(O12774));
  NOR2X1 G15214 (.A1(W2603), .A2(W5832), .ZN(W7883));
  NOR2X1 G15215 (.A1(I1768), .A2(W4694), .ZN(O205));
  NOR2X1 G15216 (.A1(W12346), .A2(W7901), .ZN(O4325));
  NOR2X1 G15217 (.A1(W6249), .A2(W4971), .ZN(W7855));
  NOR2X1 G15218 (.A1(W32843), .A2(W22703), .ZN(O12777));
  NOR2X1 G15219 (.A1(W11391), .A2(W4789), .ZN(O2586));
  NOR2X1 G15220 (.A1(W6082), .A2(W4286), .ZN(W7877));
  NOR2X1 G15221 (.A1(W27285), .A2(W13062), .ZN(O4324));
  NOR2X1 G15222 (.A1(W2356), .A2(W5581), .ZN(W7875));
  NOR2X1 G15223 (.A1(W5795), .A2(W1443), .ZN(W22700));
  NOR2X1 G15224 (.A1(W37041), .A2(W25882), .ZN(O12781));
  NOR2X1 G15225 (.A1(W30911), .A2(W21369), .ZN(O12819));
  NOR2X1 G15226 (.A1(I1428), .A2(W3512), .ZN(W7837));
  NOR2X1 G15227 (.A1(W4128), .A2(W16598), .ZN(O4320));
  NOR2X1 G15228 (.A1(W39276), .A2(W3382), .ZN(O12813));
  NOR2X1 G15229 (.A1(W12999), .A2(W3429), .ZN(O12814));
  NOR2X1 G15230 (.A1(I578), .A2(W10232), .ZN(W22715));
  NOR2X1 G15231 (.A1(W39344), .A2(W5025), .ZN(W43055));
  NOR2X1 G15232 (.A1(W10825), .A2(W22013), .ZN(O2591));
  NOR2X1 G15233 (.A1(W16460), .A2(W13510), .ZN(W22717));
  NOR2X1 G15234 (.A1(W527), .A2(W16636), .ZN(O12810));
  NOR2X1 G15235 (.A1(W13965), .A2(W11781), .ZN(W22718));
  NOR2X1 G15236 (.A1(W13172), .A2(W35375), .ZN(O12821));
  NOR2X1 G15237 (.A1(W301), .A2(I68), .ZN(W7823));
  NOR2X1 G15238 (.A1(W2257), .A2(I1129), .ZN(W7822));
  NOR2X1 G15239 (.A1(W5467), .A2(W805), .ZN(W7821));
  NOR2X1 G15240 (.A1(W5320), .A2(I175), .ZN(W22721));
  NOR2X1 G15241 (.A1(W7212), .A2(W7813), .ZN(W7819));
  NOR2X1 G15242 (.A1(W7693), .A2(W5752), .ZN(W8036));
  NOR2X1 G15243 (.A1(W13639), .A2(W9764), .ZN(W28033));
  NOR2X1 G15244 (.A1(W12544), .A2(W12967), .ZN(O12807));
  NOR2X1 G15245 (.A1(W8608), .A2(W18147), .ZN(O12806));
  NOR2X1 G15246 (.A1(W24124), .A2(W23261), .ZN(O12805));
  NOR2X1 G15247 (.A1(W8108), .A2(W7371), .ZN(W22711));
  NOR2X1 G15248 (.A1(W35298), .A2(I61), .ZN(O12798));
  NOR2X1 G15249 (.A1(W24690), .A2(I1706), .ZN(W43035));
  NOR2X1 G15250 (.A1(W823), .A2(I354), .ZN(O2588));
  NOR2X1 G15251 (.A1(W20572), .A2(W12593), .ZN(W22708));
  NOR2X1 G15252 (.A1(I1966), .A2(W5008), .ZN(W7849));
  NOR2X1 G15253 (.A1(W24766), .A2(W15012), .ZN(W43030));
  NOR2X1 G15254 (.A1(W31351), .A2(W33741), .ZN(O12794));
  NOR2X1 G15255 (.A1(W3356), .A2(W6758), .ZN(W7852));
  NOR2X1 G15256 (.A1(W38207), .A2(W29822), .ZN(O12792));
  NOR2X1 G15257 (.A1(W4320), .A2(W4961), .ZN(W28036));
  NOR2X1 G15258 (.A1(W12927), .A2(I215), .ZN(W28175));
  NOR2X1 G15259 (.A1(W36317), .A2(W28671), .ZN(O12506));
  NOR2X1 G15260 (.A1(W3979), .A2(I1323), .ZN(W8245));
  NOR2X1 G15261 (.A1(W4011), .A2(W31010), .ZN(O12508));
  NOR2X1 G15262 (.A1(W1729), .A2(W15832), .ZN(O12510));
  NOR2X1 G15263 (.A1(W4547), .A2(I563), .ZN(W42655));
  NOR2X1 G15264 (.A1(W5264), .A2(W1044), .ZN(W8240));
  NOR2X1 G15265 (.A1(W4466), .A2(W6933), .ZN(W8238));
  NOR2X1 G15266 (.A1(W35566), .A2(W38226), .ZN(O12512));
  NOR2X1 G15267 (.A1(I1182), .A2(W13027), .ZN(O4386));
  NOR2X1 G15268 (.A1(W33827), .A2(W35156), .ZN(O12516));
  NOR2X1 G15269 (.A1(W20004), .A2(W9522), .ZN(W22568));
  NOR2X1 G15270 (.A1(W4254), .A2(W6869), .ZN(W8233));
  NOR2X1 G15271 (.A1(I1746), .A2(W2461), .ZN(W8232));
  NOR2X1 G15272 (.A1(W30045), .A2(W23697), .ZN(O12519));
  NOR2X1 G15273 (.A1(W2849), .A2(W3349), .ZN(W8230));
  NOR2X1 G15274 (.A1(W813), .A2(W24911), .ZN(O12521));
  NOR2X1 G15275 (.A1(W7217), .A2(W11390), .ZN(W28183));
  NOR2X1 G15276 (.A1(W4265), .A2(W5226), .ZN(W22557));
  NOR2X1 G15277 (.A1(W5090), .A2(W7434), .ZN(O219));
  NOR2X1 G15278 (.A1(W23636), .A2(W6625), .ZN(O12496));
  NOR2X1 G15279 (.A1(W2546), .A2(W9653), .ZN(O12498));
  NOR2X1 G15280 (.A1(W726), .A2(W5862), .ZN(W8259));
  NOR2X1 G15281 (.A1(W7852), .A2(W14732), .ZN(O4388));
  NOR2X1 G15282 (.A1(W87), .A2(W1680), .ZN(W8257));
  NOR2X1 G15283 (.A1(W21852), .A2(W24786), .ZN(O12499));
  NOR2X1 G15284 (.A1(W6622), .A2(I885), .ZN(W8228));
  NOR2X1 G15285 (.A1(W4016), .A2(W10659), .ZN(O4387));
  NOR2X1 G15286 (.A1(I834), .A2(W378), .ZN(W8253));
  NOR2X1 G15287 (.A1(W851), .A2(W18398), .ZN(W22561));
  NOR2X1 G15288 (.A1(I668), .A2(W26129), .ZN(W28180));
  NOR2X1 G15289 (.A1(W6860), .A2(W5289), .ZN(W8250));
  NOR2X1 G15290 (.A1(W6622), .A2(W1757), .ZN(O217));
  NOR2X1 G15291 (.A1(W12545), .A2(W5415), .ZN(W22563));
  NOR2X1 G15292 (.A1(W355), .A2(W3473), .ZN(W8199));
  NOR2X1 G15293 (.A1(W24764), .A2(W24309), .ZN(O4384));
  NOR2X1 G15294 (.A1(W5948), .A2(W2797), .ZN(W28172));
  NOR2X1 G15295 (.A1(W2211), .A2(W6649), .ZN(W8207));
  NOR2X1 G15296 (.A1(W2193), .A2(W8076), .ZN(W8206));
  NOR2X1 G15297 (.A1(W1646), .A2(W100), .ZN(W8204));
  NOR2X1 G15298 (.A1(W2880), .A2(W33485), .ZN(O12538));
  NOR2X1 G15299 (.A1(W5130), .A2(W10264), .ZN(W28168));
  NOR2X1 G15300 (.A1(W24102), .A2(W10559), .ZN(O4381));
  NOR2X1 G15301 (.A1(W19484), .A2(W806), .ZN(W22574));
  NOR2X1 G15302 (.A1(W24721), .A2(W37367), .ZN(O12542));
  NOR2X1 G15303 (.A1(W29572), .A2(W6939), .ZN(O12543));
  NOR2X1 G15304 (.A1(W460), .A2(W326), .ZN(W8196));
  NOR2X1 G15305 (.A1(W16913), .A2(W16343), .ZN(W28166));
  NOR2X1 G15306 (.A1(W6426), .A2(W34688), .ZN(O12545));
  NOR2X1 G15307 (.A1(W10821), .A2(W19249), .ZN(O12546));
  NOR2X1 G15308 (.A1(W4848), .A2(W2648), .ZN(W8191));
  NOR2X1 G15309 (.A1(I1493), .A2(W6382), .ZN(W8218));
  NOR2X1 G15310 (.A1(W3407), .A2(W10941), .ZN(W22569));
  NOR2X1 G15311 (.A1(W3622), .A2(W30726), .ZN(W42670));
  NOR2X1 G15312 (.A1(W916), .A2(W5384), .ZN(W8225));
  NOR2X1 G15313 (.A1(W10059), .A2(W7611), .ZN(W22570));
  NOR2X1 G15314 (.A1(W26198), .A2(W25986), .ZN(W42673));
  NOR2X1 G15315 (.A1(W1312), .A2(W1830), .ZN(W8222));
  NOR2X1 G15316 (.A1(W16161), .A2(W35994), .ZN(W42674));
  NOR2X1 G15317 (.A1(W19856), .A2(W6476), .ZN(W22571));
  NOR2X1 G15318 (.A1(W6708), .A2(I338), .ZN(W8264));
  NOR2X1 G15319 (.A1(W832), .A2(W4937), .ZN(W8217));
  NOR2X1 G15320 (.A1(W16736), .A2(W5439), .ZN(W22573));
  NOR2X1 G15321 (.A1(W3679), .A2(W2993), .ZN(W8215));
  NOR2X1 G15322 (.A1(W7377), .A2(W40674), .ZN(O12530));
  NOR2X1 G15323 (.A1(W5433), .A2(W3281), .ZN(W8213));
  NOR2X1 G15324 (.A1(W5939), .A2(W3853), .ZN(W8212));
  NOR2X1 G15325 (.A1(W4546), .A2(W6462), .ZN(W8211));
  NOR2X1 G15326 (.A1(W673), .A2(W6018), .ZN(W8312));
  NOR2X1 G15327 (.A1(W22097), .A2(W19934), .ZN(O4400));
  NOR2X1 G15328 (.A1(W6325), .A2(W20025), .ZN(W22540));
  NOR2X1 G15329 (.A1(W11887), .A2(W35310), .ZN(W42575));
  NOR2X1 G15330 (.A1(W10650), .A2(I1255), .ZN(O12451));
  NOR2X1 G15331 (.A1(W2243), .A2(W3875), .ZN(W8316));
  NOR2X1 G15332 (.A1(W1896), .A2(W2305), .ZN(W8315));
  NOR2X1 G15333 (.A1(W9559), .A2(W27363), .ZN(O12452));
  NOR2X1 G15334 (.A1(I351), .A2(W7737), .ZN(W8313));
  NOR2X1 G15335 (.A1(W6137), .A2(W5305), .ZN(W8321));
  NOR2X1 G15336 (.A1(W16148), .A2(I1666), .ZN(W22541));
  NOR2X1 G15337 (.A1(W18261), .A2(W17631), .ZN(O12454));
  NOR2X1 G15338 (.A1(W5278), .A2(W3933), .ZN(W8309));
  NOR2X1 G15339 (.A1(W22979), .A2(W17373), .ZN(O12455));
  NOR2X1 G15340 (.A1(W30272), .A2(W18098), .ZN(O12456));
  NOR2X1 G15341 (.A1(W36555), .A2(W494), .ZN(O12457));
  NOR2X1 G15342 (.A1(W27905), .A2(W40071), .ZN(W42585));
  NOR2X1 G15343 (.A1(I60), .A2(W3680), .ZN(W8329));
  NOR2X1 G15344 (.A1(W3884), .A2(W12443), .ZN(O2543));
  NOR2X1 G15345 (.A1(W3214), .A2(W1204), .ZN(W8337));
  NOR2X1 G15346 (.A1(W5918), .A2(W7117), .ZN(O223));
  NOR2X1 G15347 (.A1(W19038), .A2(I1759), .ZN(O4402));
  NOR2X1 G15348 (.A1(I1819), .A2(W1558), .ZN(W8334));
  NOR2X1 G15349 (.A1(I1633), .A2(W4806), .ZN(W8333));
  NOR2X1 G15350 (.A1(W19753), .A2(W26627), .ZN(W28211));
  NOR2X1 G15351 (.A1(W4720), .A2(W254), .ZN(O4401));
  NOR2X1 G15352 (.A1(W2064), .A2(W3333), .ZN(W8302));
  NOR2X1 G15353 (.A1(W34158), .A2(W12777), .ZN(O12446));
  NOR2X1 G15354 (.A1(W15579), .A2(W16849), .ZN(W28209));
  NOR2X1 G15355 (.A1(W4479), .A2(W586), .ZN(W8326));
  NOR2X1 G15356 (.A1(I432), .A2(W1492), .ZN(W8325));
  NOR2X1 G15357 (.A1(W2329), .A2(W7556), .ZN(W8324));
  NOR2X1 G15358 (.A1(I268), .A2(W2352), .ZN(W8323));
  NOR2X1 G15359 (.A1(W504), .A2(W41681), .ZN(O12448));
  NOR2X1 G15360 (.A1(W4091), .A2(W36424), .ZN(W42631));
  NOR2X1 G15361 (.A1(W14236), .A2(W11063), .ZN(W42616));
  NOR2X1 G15362 (.A1(W7170), .A2(W6230), .ZN(W8284));
  NOR2X1 G15363 (.A1(W1515), .A2(W942), .ZN(W8283));
  NOR2X1 G15364 (.A1(W7755), .A2(W17963), .ZN(O12480));
  NOR2X1 G15365 (.A1(W8224), .A2(I1895), .ZN(W8280));
  NOR2X1 G15366 (.A1(W17749), .A2(W6338), .ZN(O12484));
  NOR2X1 G15367 (.A1(I272), .A2(W2567), .ZN(O12486));
  NOR2X1 G15368 (.A1(W9810), .A2(W2733), .ZN(O2547));
  NOR2X1 G15369 (.A1(W30943), .A2(W38746), .ZN(W42614));
  NOR2X1 G15370 (.A1(I1418), .A2(I1092), .ZN(W8273));
  NOR2X1 G15371 (.A1(W2359), .A2(W1229), .ZN(O220));
  NOR2X1 G15372 (.A1(W4849), .A2(I309), .ZN(W8270));
  NOR2X1 G15373 (.A1(W6060), .A2(W1246), .ZN(W8269));
  NOR2X1 G15374 (.A1(I1930), .A2(W4490), .ZN(W8268));
  NOR2X1 G15375 (.A1(W12457), .A2(W5328), .ZN(W42633));
  NOR2X1 G15376 (.A1(W22050), .A2(W21953), .ZN(O12493));
  NOR2X1 G15377 (.A1(W37359), .A2(W33149), .ZN(O12547));
  NOR2X1 G15378 (.A1(W6145), .A2(W2901), .ZN(W8287));
  NOR2X1 G15379 (.A1(W15094), .A2(W7486), .ZN(W28194));
  NOR2X1 G15380 (.A1(W40275), .A2(W150), .ZN(O12476));
  NOR2X1 G15381 (.A1(W14608), .A2(W12979), .ZN(W42609));
  NOR2X1 G15382 (.A1(W6727), .A2(W8243), .ZN(W8291));
  NOR2X1 G15383 (.A1(W8826), .A2(W12472), .ZN(W42605));
  NOR2X1 G15384 (.A1(W2593), .A2(W11254), .ZN(O4395));
  NOR2X1 G15385 (.A1(W20026), .A2(W23947), .ZN(W28199));
  NOR2X1 G15386 (.A1(W14836), .A2(W27632), .ZN(W28200));
  NOR2X1 G15387 (.A1(W24846), .A2(W16731), .ZN(W42599));
  NOR2X1 G15388 (.A1(W2825), .A2(W6063), .ZN(W8297));
  NOR2X1 G15389 (.A1(W17281), .A2(W2231), .ZN(W22546));
  NOR2X1 G15390 (.A1(W100), .A2(W638), .ZN(O4397));
  NOR2X1 G15391 (.A1(W20595), .A2(W11834), .ZN(W28203));
  NOR2X1 G15392 (.A1(W24830), .A2(W17186), .ZN(O12461));
  NOR2X1 G15393 (.A1(W4174), .A2(W5086), .ZN(O4356));
  NOR2X1 G15394 (.A1(I496), .A2(W7840), .ZN(W8093));
  NOR2X1 G15395 (.A1(W10788), .A2(W13873), .ZN(O12615));
  NOR2X1 G15396 (.A1(W3607), .A2(W2191), .ZN(W8090));
  NOR2X1 G15397 (.A1(W9977), .A2(W1690), .ZN(O12617));
  NOR2X1 G15398 (.A1(I1391), .A2(I151), .ZN(W8088));
  NOR2X1 G15399 (.A1(W1456), .A2(W1384), .ZN(W8087));
  NOR2X1 G15400 (.A1(W573), .A2(W29688), .ZN(W42796));
  NOR2X1 G15401 (.A1(I132), .A2(W7257), .ZN(W8085));
  NOR2X1 G15402 (.A1(W1824), .A2(W1337), .ZN(W8094));
  NOR2X1 G15403 (.A1(I1914), .A2(I619), .ZN(W8083));
  NOR2X1 G15404 (.A1(W8128), .A2(W16501), .ZN(O2559));
  NOR2X1 G15405 (.A1(W3832), .A2(W4783), .ZN(W8080));
  NOR2X1 G15406 (.A1(W14774), .A2(W17898), .ZN(O12622));
  NOR2X1 G15407 (.A1(W25645), .A2(W41780), .ZN(O12624));
  NOR2X1 G15408 (.A1(I1960), .A2(W2189), .ZN(W8077));
  NOR2X1 G15409 (.A1(W34078), .A2(W4355), .ZN(O12625));
  NOR2X1 G15410 (.A1(W7216), .A2(W3971), .ZN(W8103));
  NOR2X1 G15411 (.A1(W5029), .A2(W8022), .ZN(W8111));
  NOR2X1 G15412 (.A1(W3306), .A2(W6163), .ZN(W8110));
  NOR2X1 G15413 (.A1(W6059), .A2(W16023), .ZN(O12610));
  NOR2X1 G15414 (.A1(W7251), .A2(W30503), .ZN(W42782));
  NOR2X1 G15415 (.A1(W6223), .A2(W1094), .ZN(W8107));
  NOR2X1 G15416 (.A1(W19380), .A2(W27608), .ZN(W28125));
  NOR2X1 G15417 (.A1(W9021), .A2(W27367), .ZN(W28124));
  NOR2X1 G15418 (.A1(W915), .A2(W5942), .ZN(W8104));
  NOR2X1 G15419 (.A1(W18326), .A2(W3171), .ZN(O4354));
  NOR2X1 G15420 (.A1(W6441), .A2(W7561), .ZN(W8102));
  NOR2X1 G15421 (.A1(I1333), .A2(W1289), .ZN(W8101));
  NOR2X1 G15422 (.A1(W3596), .A2(W4708), .ZN(W8100));
  NOR2X1 G15423 (.A1(W20290), .A2(W6443), .ZN(W22617));
  NOR2X1 G15424 (.A1(I56), .A2(I1575), .ZN(W8097));
  NOR2X1 G15425 (.A1(I793), .A2(W17303), .ZN(O4359));
  NOR2X1 G15426 (.A1(W66), .A2(I75), .ZN(W8095));
  NOR2X1 G15427 (.A1(W8337), .A2(W15154), .ZN(W28096));
  NOR2X1 G15428 (.A1(W13037), .A2(W15566), .ZN(W28106));
  NOR2X1 G15429 (.A1(W7468), .A2(W12709), .ZN(O12645));
  NOR2X1 G15430 (.A1(W14296), .A2(W12086), .ZN(W28104));
  NOR2X1 G15431 (.A1(I1620), .A2(W4793), .ZN(W8051));
  NOR2X1 G15432 (.A1(W299), .A2(W3959), .ZN(W8050));
  NOR2X1 G15433 (.A1(W14596), .A2(W23348), .ZN(W28100));
  NOR2X1 G15434 (.A1(W25124), .A2(W18539), .ZN(O12653));
  NOR2X1 G15435 (.A1(W35565), .A2(W35432), .ZN(O12654));
  NOR2X1 G15436 (.A1(W4602), .A2(W18985), .ZN(W22631));
  NOR2X1 G15437 (.A1(W4980), .A2(W682), .ZN(W8043));
  NOR2X1 G15438 (.A1(W12055), .A2(W25446), .ZN(O4345));
  NOR2X1 G15439 (.A1(W28336), .A2(W16078), .ZN(W42846));
  NOR2X1 G15440 (.A1(W6544), .A2(W7634), .ZN(W8040));
  NOR2X1 G15441 (.A1(W40082), .A2(W33030), .ZN(O12659));
  NOR2X1 G15442 (.A1(W27232), .A2(W17458), .ZN(W28092));
  NOR2X1 G15443 (.A1(I646), .A2(W24857), .ZN(W28091));
  NOR2X1 G15444 (.A1(I552), .A2(I1640), .ZN(O2557));
  NOR2X1 G15445 (.A1(W36178), .A2(W1748), .ZN(W42824));
  NOR2X1 G15446 (.A1(W1344), .A2(W3639), .ZN(W28107));
  NOR2X1 G15447 (.A1(W2471), .A2(W12157), .ZN(W22629));
  NOR2X1 G15448 (.A1(W4080), .A2(I1959), .ZN(W8062));
  NOR2X1 G15449 (.A1(W28270), .A2(W7789), .ZN(O12640));
  NOR2X1 G15450 (.A1(W15331), .A2(W18202), .ZN(O4350));
  NOR2X1 G15451 (.A1(W21629), .A2(W32338), .ZN(O12638));
  NOR2X1 G15452 (.A1(W10234), .A2(W32319), .ZN(W42816));
  NOR2X1 G15453 (.A1(W5112), .A2(W5553), .ZN(W8067));
  NOR2X1 G15454 (.A1(W298), .A2(W5513), .ZN(W22627));
  NOR2X1 G15455 (.A1(W203), .A2(W5141), .ZN(W22626));
  NOR2X1 G15456 (.A1(W8946), .A2(W14691), .ZN(O12631));
  NOR2X1 G15457 (.A1(I354), .A2(W18979), .ZN(O4351));
  NOR2X1 G15458 (.A1(W32604), .A2(W30870), .ZN(O12628));
  NOR2X1 G15459 (.A1(W3583), .A2(W2921), .ZN(O12627));
  NOR2X1 G15460 (.A1(I1118), .A2(W1262), .ZN(W8162));
  NOR2X1 G15461 (.A1(W32166), .A2(W30468), .ZN(O12567));
  NOR2X1 G15462 (.A1(W2753), .A2(W36664), .ZN(O12568));
  NOR2X1 G15463 (.A1(W23435), .A2(W41234), .ZN(O12569));
  NOR2X1 G15464 (.A1(W17485), .A2(W16376), .ZN(O4378));
  NOR2X1 G15465 (.A1(I672), .A2(I1901), .ZN(W8167));
  NOR2X1 G15466 (.A1(W10834), .A2(W19285), .ZN(W22591));
  NOR2X1 G15467 (.A1(I565), .A2(W785), .ZN(W8164));
  NOR2X1 G15468 (.A1(W21113), .A2(W9289), .ZN(O2552));
  NOR2X1 G15469 (.A1(W2664), .A2(W6089), .ZN(W8172));
  NOR2X1 G15470 (.A1(W2804), .A2(W3475), .ZN(W8161));
  NOR2X1 G15471 (.A1(W7328), .A2(W2350), .ZN(W8159));
  NOR2X1 G15472 (.A1(W27176), .A2(W15488), .ZN(W42733));
  NOR2X1 G15473 (.A1(W27993), .A2(W14610), .ZN(W28156));
  NOR2X1 G15474 (.A1(I696), .A2(I1775), .ZN(W8156));
  NOR2X1 G15475 (.A1(W997), .A2(W3254), .ZN(W8155));
  NOR2X1 G15476 (.A1(W21066), .A2(W24574), .ZN(W28153));
  NOR2X1 G15477 (.A1(W32049), .A2(W24200), .ZN(O12561));
  NOR2X1 G15478 (.A1(W1470), .A2(W6991), .ZN(W22583));
  NOR2X1 G15479 (.A1(W7266), .A2(W38608), .ZN(O12551));
  NOR2X1 G15480 (.A1(W17929), .A2(W24198), .ZN(W28164));
  NOR2X1 G15481 (.A1(W20903), .A2(W414), .ZN(W22585));
  NOR2X1 G15482 (.A1(W15805), .A2(W30061), .ZN(W42708));
  NOR2X1 G15483 (.A1(W40976), .A2(W4648), .ZN(O12556));
  NOR2X1 G15484 (.A1(W7485), .A2(W6395), .ZN(W8182));
  NOR2X1 G15485 (.A1(W22407), .A2(I1956), .ZN(O12557));
  NOR2X1 G15486 (.A1(I875), .A2(W6628), .ZN(W22596));
  NOR2X1 G15487 (.A1(W4946), .A2(W15759), .ZN(W22587));
  NOR2X1 G15488 (.A1(W22550), .A2(W6331), .ZN(O2551));
  NOR2X1 G15489 (.A1(W12113), .A2(W20261), .ZN(O12564));
  NOR2X1 G15490 (.A1(W10406), .A2(W5616), .ZN(W42723));
  NOR2X1 G15491 (.A1(I428), .A2(I501), .ZN(W8175));
  NOR2X1 G15492 (.A1(W6858), .A2(W8145), .ZN(W8174));
  NOR2X1 G15493 (.A1(W703), .A2(W3818), .ZN(W8173));
  NOR2X1 G15494 (.A1(W13088), .A2(W38506), .ZN(W42769));
  NOR2X1 G15495 (.A1(W31740), .A2(W6611), .ZN(W42752));
  NOR2X1 G15496 (.A1(W20763), .A2(W11038), .ZN(W28145));
  NOR2X1 G15497 (.A1(W23850), .A2(W13150), .ZN(W28142));
  NOR2X1 G15498 (.A1(W6625), .A2(W1340), .ZN(W8132));
  NOR2X1 G15499 (.A1(W4257), .A2(W641), .ZN(W8129));
  NOR2X1 G15500 (.A1(I1372), .A2(W6490), .ZN(W8128));
  NOR2X1 G15501 (.A1(W19200), .A2(W13870), .ZN(O4368));
  NOR2X1 G15502 (.A1(W28082), .A2(W24178), .ZN(O4366));
  NOR2X1 G15503 (.A1(W5829), .A2(W581), .ZN(W8136));
  NOR2X1 G15504 (.A1(I1744), .A2(W2856), .ZN(W8121));
  NOR2X1 G15505 (.A1(I267), .A2(W28686), .ZN(W42770));
  NOR2X1 G15506 (.A1(W8382), .A2(W29370), .ZN(W42773));
  NOR2X1 G15507 (.A1(W37199), .A2(I1461), .ZN(O12604));
  NOR2X1 G15508 (.A1(W2930), .A2(W3570), .ZN(W8117));
  NOR2X1 G15509 (.A1(W25679), .A2(W10745), .ZN(O12605));
  NOR2X1 G15510 (.A1(I1676), .A2(W6098), .ZN(W8115));
  NOR2X1 G15511 (.A1(W16902), .A2(W15108), .ZN(O13467));
  NOR2X1 G15512 (.A1(W13157), .A2(W5367), .ZN(W28148));
  NOR2X1 G15513 (.A1(W2689), .A2(W7639), .ZN(W8138));
  NOR2X1 G15514 (.A1(W8011), .A2(W17282), .ZN(W22600));
  NOR2X1 G15515 (.A1(W3619), .A2(W5319), .ZN(W8140));
  NOR2X1 G15516 (.A1(W16990), .A2(W41152), .ZN(O12585));
  NOR2X1 G15517 (.A1(W18255), .A2(I1883), .ZN(O12583));
  NOR2X1 G15518 (.A1(W957), .A2(W4386), .ZN(W8144));
  NOR2X1 G15519 (.A1(W18311), .A2(W41732), .ZN(O12580));
  NOR2X1 G15520 (.A1(W8119), .A2(W6706), .ZN(W8146));
  NOR2X1 G15521 (.A1(W5665), .A2(W15129), .ZN(O12579));
  NOR2X1 G15522 (.A1(W6511), .A2(W23914), .ZN(W28152));
  NOR2X1 G15523 (.A1(W5237), .A2(W21360), .ZN(W22597));
  NOR2X1 G15524 (.A1(W6944), .A2(W4331), .ZN(W8150));
  NOR2X1 G15525 (.A1(W26394), .A2(W37739), .ZN(W42738));
  NOR2X1 G15526 (.A1(W5690), .A2(I1266), .ZN(W8152));
  NOR2X1 G15527 (.A1(I1546), .A2(W5516), .ZN(W6129));
  NOR2X1 G15528 (.A1(I710), .A2(W5029), .ZN(W6125));
  NOR2X1 G15529 (.A1(W35156), .A2(W39681), .ZN(W45569));
  NOR2X1 G15530 (.A1(W37329), .A2(W34190), .ZN(O14195));
  NOR2X1 G15531 (.A1(W14690), .A2(W40299), .ZN(O14945));
  NOR2X1 G15532 (.A1(W2633), .A2(W3482), .ZN(W6127));
  NOR2X1 G15533 (.A1(W13095), .A2(W13830), .ZN(O14946));
  NOR2X1 G15534 (.A1(W2818), .A2(W20), .ZN(W5733));
  NOR2X1 G15535 (.A1(I1574), .A2(W1209), .ZN(W5484));
  NOR2X1 G15536 (.A1(W11827), .A2(W10778), .ZN(O14389));
  NOR2X1 G15537 (.A1(W1978), .A2(W4120), .ZN(W6128));
  NOR2X1 G15538 (.A1(W6573), .A2(W15458), .ZN(W27227));
  NOR2X1 G15539 (.A1(I1425), .A2(W1877), .ZN(W6130));
  NOR2X1 G15540 (.A1(I1585), .A2(W4792), .ZN(W5732));
  NOR2X1 G15541 (.A1(W11371), .A2(W8166), .ZN(O14510));
  NOR2X1 G15542 (.A1(I1368), .A2(W1264), .ZN(W23425));
  NOR2X1 G15543 (.A1(W5347), .A2(W33642), .ZN(O14947));
  NOR2X1 G15544 (.A1(W3711), .A2(W896), .ZN(W5226));
  NOR2X1 G15545 (.A1(W17370), .A2(W30351), .ZN(O14191));
  NOR2X1 G15546 (.A1(I1606), .A2(W4000), .ZN(W44794));
  NOR2X1 G15547 (.A1(W38132), .A2(W36846), .ZN(O14515));
  NOR2X1 G15548 (.A1(I1091), .A2(W5121), .ZN(W5422));
  NOR2X1 G15549 (.A1(W45337), .A2(W37601), .ZN(W45443));
  NOR2X1 G15550 (.A1(W1374), .A2(W45206), .ZN(O14726));
  NOR2X1 G15551 (.A1(W3680), .A2(W2404), .ZN(W5365));
  NOR2X1 G15552 (.A1(I1667), .A2(W39547), .ZN(O14205));
  NOR2X1 G15553 (.A1(W9561), .A2(W34012), .ZN(W45445));
  NOR2X1 G15554 (.A1(W291), .A2(W410), .ZN(W6117));
  NOR2X1 G15555 (.A1(W14578), .A2(I52), .ZN(O14204));
  NOR2X1 G15556 (.A1(W4323), .A2(W2599), .ZN(W5891));
  NOR2X1 G15557 (.A1(W627), .A2(I1597), .ZN(W6119));
  NOR2X1 G15558 (.A1(W27060), .A2(W9291), .ZN(W27438));
  NOR2X1 G15559 (.A1(W28569), .A2(W17157), .ZN(O14202));
  NOR2X1 G15560 (.A1(W9785), .A2(W6122), .ZN(W23427));
  NOR2X1 G15561 (.A1(W16570), .A2(W7217), .ZN(W23291));
  NOR2X1 G15562 (.A1(W14527), .A2(W4291), .ZN(O14506));
  NOR2X1 G15563 (.A1(W3336), .A2(W17525), .ZN(W23511));
  NOR2X1 G15564 (.A1(W35526), .A2(I1495), .ZN(O14198));
  NOR2X1 G15565 (.A1(W36795), .A2(W38982), .ZN(O14196));
  NOR2X1 G15566 (.A1(W4289), .A2(W4445), .ZN(W5231));
  NOR2X1 G15567 (.A1(I683), .A2(W404), .ZN(W5734));
  NOR2X1 G15568 (.A1(W11982), .A2(W8281), .ZN(O14722));
  NOR2X1 G15569 (.A1(W1179), .A2(W19482), .ZN(W27129));
  NOR2X1 G15570 (.A1(W5276), .A2(W20469), .ZN(O3993));
  NOR2X1 G15571 (.A1(W27156), .A2(W25728), .ZN(O14774));
  NOR2X1 G15572 (.A1(W19684), .A2(W860), .ZN(W23431));
  NOR2X1 G15573 (.A1(W19341), .A2(W9285), .ZN(W45566));
  NOR2X1 G15574 (.A1(W24008), .A2(W13532), .ZN(W27230));
  NOR2X1 G15575 (.A1(W29971), .A2(W28689), .ZN(O14823));
  NOR2X1 G15576 (.A1(W16335), .A2(W41718), .ZN(O14524));
  NOR2X1 G15577 (.A1(W17922), .A2(W23569), .ZN(W44789));
  NOR2X1 G15578 (.A1(I1294), .A2(I184), .ZN(W5370));
  NOR2X1 G15579 (.A1(W27325), .A2(W33402), .ZN(O14526));
  NOR2X1 G15580 (.A1(W23471), .A2(W7308), .ZN(O14718));
  NOR2X1 G15581 (.A1(I748), .A2(W865), .ZN(W6140));
  NOR2X1 G15582 (.A1(W5433), .A2(W8244), .ZN(W23603));
  NOR2X1 G15583 (.A1(W19618), .A2(W22097), .ZN(O14392));
  NOR2X1 G15584 (.A1(W10338), .A2(W29744), .ZN(O14185));
  NOR2X1 G15585 (.A1(W1665), .A2(W4899), .ZN(W5217));
  NOR2X1 G15586 (.A1(W15525), .A2(W9540), .ZN(O14393));
  NOR2X1 G15587 (.A1(I1572), .A2(W18060), .ZN(W27232));
  NOR2X1 G15588 (.A1(W1705), .A2(W5468), .ZN(W6143));
  NOR2X1 G15589 (.A1(I1825), .A2(W3259), .ZN(W23288));
  NOR2X1 G15590 (.A1(I726), .A2(W5045), .ZN(W6145));
  NOR2X1 G15591 (.A1(W15722), .A2(W38825), .ZN(O14520));
  NOR2X1 G15592 (.A1(W19209), .A2(W23483), .ZN(O14189));
  NOR2X1 G15593 (.A1(W27286), .A2(W29077), .ZN(O14948));
  NOR2X1 G15594 (.A1(W3244), .A2(W5491), .ZN(W6135));
  NOR2X1 G15595 (.A1(W8691), .A2(W3567), .ZN(W27312));
  NOR2X1 G15596 (.A1(W11386), .A2(W3721), .ZN(W23289));
  NOR2X1 G15597 (.A1(W6796), .A2(W248), .ZN(O2771));
  NOR2X1 G15598 (.A1(W43587), .A2(W21859), .ZN(O14390));
  NOR2X1 G15599 (.A1(W2336), .A2(W3728), .ZN(W5724));
  NOR2X1 G15600 (.A1(W23579), .A2(W10634), .ZN(W44790));
  NOR2X1 G15601 (.A1(W17777), .A2(W19361), .ZN(W27179));
  NOR2X1 G15602 (.A1(W228), .A2(W5173), .ZN(W6115));
  NOR2X1 G15603 (.A1(W667), .A2(W11078), .ZN(W23373));
  NOR2X1 G15604 (.A1(W3202), .A2(W18310), .ZN(W23599));
  NOR2X1 G15605 (.A1(W5366), .A2(W981), .ZN(W5722));
  NOR2X1 G15606 (.A1(W26708), .A2(W19481), .ZN(W27125));
  NOR2X1 G15607 (.A1(W21029), .A2(W5911), .ZN(W27310));
  NOR2X1 G15608 (.A1(W15233), .A2(W33739), .ZN(W45720));
  NOR2X1 G15609 (.A1(I884), .A2(I1656), .ZN(W6138));
  NOR2X1 G15610 (.A1(I1140), .A2(W426), .ZN(W6139));
  NOR2X1 G15611 (.A1(W30262), .A2(W30001), .ZN(O14522));
  NOR2X1 G15612 (.A1(I1856), .A2(W5929), .ZN(W6090));
  NOR2X1 G15613 (.A1(W19013), .A2(W36388), .ZN(W44844));
  NOR2X1 G15614 (.A1(W16605), .A2(W13527), .ZN(O2737));
  NOR2X1 G15615 (.A1(W1796), .A2(W3097), .ZN(W5469));
  NOR2X1 G15616 (.A1(W39768), .A2(W40392), .ZN(O14732));
  NOR2X1 G15617 (.A1(W6727), .A2(W1962), .ZN(O14923));
  NOR2X1 G15618 (.A1(W25278), .A2(W931), .ZN(W44842));
  NOR2X1 G15619 (.A1(W21894), .A2(W2254), .ZN(O14229));
  NOR2X1 G15620 (.A1(W1630), .A2(W13621), .ZN(O14228));
  NOR2X1 G15621 (.A1(W39292), .A2(W36593), .ZN(O14384));
  NOR2X1 G15622 (.A1(W5574), .A2(W5649), .ZN(W6089));
  NOR2X1 G15623 (.A1(W7929), .A2(W16473), .ZN(W23515));
  NOR2X1 G15624 (.A1(W983), .A2(I530), .ZN(W5805));
  NOR2X1 G15625 (.A1(W2914), .A2(W3079), .ZN(W6091));
  NOR2X1 G15626 (.A1(W6581), .A2(W2709), .ZN(O4020));
  NOR2X1 G15627 (.A1(W29490), .A2(W2896), .ZN(O14227));
  NOR2X1 G15628 (.A1(W3466), .A2(W1781), .ZN(W5741));
  NOR2X1 G15629 (.A1(I912), .A2(W17944), .ZN(O14461));
  NOR2X1 G15630 (.A1(I1337), .A2(I1407), .ZN(W6094));
  NOR2X1 G15631 (.A1(W27967), .A2(W40934), .ZN(O14827));
  NOR2X1 G15632 (.A1(I20), .A2(W1759), .ZN(W5247));
  NOR2X1 G15633 (.A1(W12633), .A2(W34059), .ZN(O14380));
  NOR2X1 G15634 (.A1(W2496), .A2(W1397), .ZN(W6073));
  NOR2X1 G15635 (.A1(W17865), .A2(W15657), .ZN(O14239));
  NOR2X1 G15636 (.A1(W36644), .A2(W37611), .ZN(W44852));
  NOR2X1 G15637 (.A1(W14301), .A2(W38530), .ZN(O14735));
  NOR2X1 G15638 (.A1(W2622), .A2(I1726), .ZN(W5900));
  NOR2X1 G15639 (.A1(W4309), .A2(I1054), .ZN(W5744));
  NOR2X1 G15640 (.A1(W18950), .A2(W26775), .ZN(O14921));
  NOR2X1 G15641 (.A1(W2678), .A2(W5717), .ZN(W6077));
  NOR2X1 G15642 (.A1(W4439), .A2(W7659), .ZN(O4101));
  NOR2X1 G15643 (.A1(W10172), .A2(W28910), .ZN(O14378));
  NOR2X1 G15644 (.A1(W1612), .A2(W5202), .ZN(O86));
  NOR2X1 G15645 (.A1(W33052), .A2(W3258), .ZN(O14235));
  NOR2X1 G15646 (.A1(I1921), .A2(W3310), .ZN(W6080));
  NOR2X1 G15647 (.A1(W1042), .A2(W3192), .ZN(W5249));
  NOR2X1 G15648 (.A1(W10329), .A2(W25071), .ZN(W27222));
  NOR2X1 G15649 (.A1(W1410), .A2(W5670), .ZN(O106));
  NOR2X1 G15650 (.A1(W26905), .A2(W21600), .ZN(O14233));
  NOR2X1 G15651 (.A1(I1639), .A2(W7581), .ZN(W45033));
  NOR2X1 G15652 (.A1(W2540), .A2(W3451), .ZN(W6082));
  NOR2X1 G15653 (.A1(W5162), .A2(W5899), .ZN(W27431));
  NOR2X1 G15654 (.A1(W20436), .A2(W41165), .ZN(W44820));
  NOR2X1 G15655 (.A1(W43843), .A2(W18665), .ZN(O14932));
  NOR2X1 G15656 (.A1(W17716), .A2(W38219), .ZN(O14934));
  NOR2X1 G15657 (.A1(W26657), .A2(W41056), .ZN(W45699));
  NOR2X1 G15658 (.A1(W2065), .A2(W3706), .ZN(W5893));
  NOR2X1 G15659 (.A1(W13197), .A2(W20608), .ZN(W23296));
  NOR2X1 G15660 (.A1(W17957), .A2(W4048), .ZN(O14212));
  NOR2X1 G15661 (.A1(W6634), .A2(W44135), .ZN(W45570));
  NOR2X1 G15662 (.A1(W5326), .A2(W1167), .ZN(W5473));
  NOR2X1 G15663 (.A1(W1125), .A2(W1088), .ZN(W27372));
  NOR2X1 G15664 (.A1(W8479), .A2(W1721), .ZN(W23295));
  NOR2X1 G15665 (.A1(W2620), .A2(W4430), .ZN(W6105));
  NOR2X1 G15666 (.A1(W15365), .A2(W16011), .ZN(O4103));
  NOR2X1 G15667 (.A1(W56), .A2(W27635), .ZN(O14208));
  NOR2X1 G15668 (.A1(W3552), .A2(W923), .ZN(W6112));
  NOR2X1 G15669 (.A1(W9432), .A2(W34963), .ZN(O14729));
  NOR2X1 G15670 (.A1(W16976), .A2(W2847), .ZN(W23595));
  NOR2X1 G15671 (.A1(W8676), .A2(W39600), .ZN(W45449));
  NOR2X1 G15672 (.A1(I1701), .A2(W16758), .ZN(W45704));
  NOR2X1 G15673 (.A1(W3254), .A2(W37220), .ZN(O14505));
  NOR2X1 G15674 (.A1(W10805), .A2(W43095), .ZN(O14206));
  NOR2X1 G15675 (.A1(W5433), .A2(I1766), .ZN(W5737));
  NOR2X1 G15676 (.A1(I1962), .A2(W945), .ZN(W5246));
  NOR2X1 G15677 (.A1(W25655), .A2(I1599), .ZN(O14502));
  NOR2X1 G15678 (.A1(W13518), .A2(W22430), .ZN(W27433));
  NOR2X1 G15679 (.A1(W38281), .A2(W35303), .ZN(O14224));
  NOR2X1 G15680 (.A1(W31208), .A2(W13940), .ZN(O14924));
  NOR2X1 G15681 (.A1(W2665), .A2(W1727), .ZN(W6097));
  NOR2X1 G15682 (.A1(W8729), .A2(W10722), .ZN(W23300));
  NOR2X1 G15683 (.A1(W5402), .A2(W2850), .ZN(W5739));
  NOR2X1 G15684 (.A1(W10849), .A2(W17938), .ZN(O14221));
  NOR2X1 G15685 (.A1(W33992), .A2(W23103), .ZN(O14460));
  NOR2X1 G15686 (.A1(I1267), .A2(W4079), .ZN(W5489));
  NOR2X1 G15687 (.A1(W27302), .A2(W12556), .ZN(W27435));
  NOR2X1 G15688 (.A1(W1502), .A2(W22906), .ZN(W27178));
  NOR2X1 G15689 (.A1(W42895), .A2(W21247), .ZN(O14386));
  NOR2X1 G15690 (.A1(W4360), .A2(W4496), .ZN(W6102));
  NOR2X1 G15691 (.A1(W7973), .A2(W38796), .ZN(O14929));
  NOR2X1 G15692 (.A1(I956), .A2(W15692), .ZN(W23297));
  NOR2X1 G15693 (.A1(W8239), .A2(W17489), .ZN(O2822));
  NOR2X1 G15694 (.A1(W23741), .A2(W27332), .ZN(O14216));
  NOR2X1 G15695 (.A1(W4890), .A2(W2995), .ZN(W5240));
  NOR2X1 G15696 (.A1(W42508), .A2(W23291), .ZN(O14149));
  NOR2X1 G15697 (.A1(W20863), .A2(W24430), .ZN(W27305));
  NOR2X1 G15698 (.A1(W27380), .A2(W32743), .ZN(O14699));
  NOR2X1 G15699 (.A1(W4900), .A2(W38908), .ZN(O14997));
  NOR2X1 G15700 (.A1(W14322), .A2(W33498), .ZN(W45121));
  NOR2X1 G15701 (.A1(W3315), .A2(W13704), .ZN(O14153));
  NOR2X1 G15702 (.A1(W1683), .A2(W21334), .ZN(W23274));
  NOR2X1 G15703 (.A1(W831), .A2(W46), .ZN(W5182));
  NOR2X1 G15704 (.A1(W28393), .A2(W104), .ZN(O14998));
  NOR2X1 G15705 (.A1(W3773), .A2(W7696), .ZN(W27457));
  NOR2X1 G15706 (.A1(I501), .A2(W22002), .ZN(W27458));
  NOR2X1 G15707 (.A1(W4670), .A2(W2229), .ZN(W5184));
  NOR2X1 G15708 (.A1(W33032), .A2(W643), .ZN(O14775));
  NOR2X1 G15709 (.A1(W18135), .A2(W6885), .ZN(O2829));
  NOR2X1 G15710 (.A1(W38168), .A2(W21923), .ZN(O14815));
  NOR2X1 G15711 (.A1(W22393), .A2(W19612), .ZN(W27303));
  NOR2X1 G15712 (.A1(W3002), .A2(W4767), .ZN(W5876));
  NOR2X1 G15713 (.A1(W19787), .A2(I1690), .ZN(O3986));
  NOR2X1 G15714 (.A1(W40759), .A2(W10140), .ZN(O14814));
  NOR2X1 G15715 (.A1(W2707), .A2(W4072), .ZN(W6196));
  NOR2X1 G15716 (.A1(W11066), .A2(W17130), .ZN(O14812));
  NOR2X1 G15717 (.A1(W24286), .A2(W17012), .ZN(O14158));
  NOR2X1 G15718 (.A1(W19155), .A2(W14229), .ZN(W27452));
  NOR2X1 G15719 (.A1(W3677), .A2(I1900), .ZN(W44753));
  NOR2X1 G15720 (.A1(I895), .A2(W6113), .ZN(W6183));
  NOR2X1 G15721 (.A1(W22885), .A2(W14350), .ZN(W27115));
  NOR2X1 G15722 (.A1(W24117), .A2(W28682), .ZN(W44751));
  NOR2X1 G15723 (.A1(I18), .A2(W2404), .ZN(W6185));
  NOR2X1 G15724 (.A1(W6259), .A2(W1526), .ZN(O14991));
  NOR2X1 G15725 (.A1(W5089), .A2(W1153), .ZN(W6186));
  NOR2X1 G15726 (.A1(W1549), .A2(I1528), .ZN(W5705));
  NOR2X1 G15727 (.A1(W14455), .A2(W15296), .ZN(O2754));
  NOR2X1 G15728 (.A1(W4837), .A2(W5580), .ZN(W5875));
  NOR2X1 G15729 (.A1(W30785), .A2(W25577), .ZN(O14536));
  NOR2X1 G15730 (.A1(W44247), .A2(I1634), .ZN(O14402));
  NOR2X1 G15731 (.A1(W402), .A2(W2590), .ZN(W5187));
  NOR2X1 G15732 (.A1(W34448), .A2(W24880), .ZN(O14154));
  NOR2X1 G15733 (.A1(W28993), .A2(W43593), .ZN(O14700));
  NOR2X1 G15734 (.A1(I1494), .A2(I912), .ZN(W5703));
  NOR2X1 G15735 (.A1(W17798), .A2(W3675), .ZN(O2828));
  NOR2X1 G15736 (.A1(W21508), .A2(W6711), .ZN(O14537));
  NOR2X1 G15737 (.A1(W2020), .A2(W2461), .ZN(W6190));
  NOR2X1 G15738 (.A1(I1528), .A2(W5801), .ZN(W6211));
  NOR2X1 G15739 (.A1(W28485), .A2(W7228), .ZN(O14129));
  NOR2X1 G15740 (.A1(W4473), .A2(W2065), .ZN(W5873));
  NOR2X1 G15741 (.A1(W9100), .A2(W30780), .ZN(O14548));
  NOR2X1 G15742 (.A1(W44241), .A2(W13974), .ZN(O14128));
  NOR2X1 G15743 (.A1(W1197), .A2(I362), .ZN(W6207));
  NOR2X1 G15744 (.A1(W2422), .A2(W1488), .ZN(W5692));
  NOR2X1 G15745 (.A1(I191), .A2(W12387), .ZN(W23621));
  NOR2X1 G15746 (.A1(W17960), .A2(W32343), .ZN(W44714));
  NOR2X1 G15747 (.A1(W8516), .A2(W3057), .ZN(W45412));
  NOR2X1 G15748 (.A1(W5382), .A2(W8967), .ZN(O14126));
  NOR2X1 G15749 (.A1(I1334), .A2(I1870), .ZN(W27107));
  NOR2X1 G15750 (.A1(W6890), .A2(W20188), .ZN(W23441));
  NOR2X1 G15751 (.A1(I1579), .A2(W1681), .ZN(W6212));
  NOR2X1 G15752 (.A1(W1696), .A2(W5157), .ZN(W5690));
  NOR2X1 G15753 (.A1(W43750), .A2(W19177), .ZN(O15011));
  NOR2X1 G15754 (.A1(W1710), .A2(W851), .ZN(W5168));
  NOR2X1 G15755 (.A1(W21047), .A2(W19414), .ZN(W27469));
  NOR2X1 G15756 (.A1(W3315), .A2(W2787), .ZN(W6214));
  NOR2X1 G15757 (.A1(W40570), .A2(W33029), .ZN(O14123));
  NOR2X1 G15758 (.A1(W5700), .A2(W2344), .ZN(W23624));
  NOR2X1 G15759 (.A1(W20746), .A2(W32672), .ZN(O14137));
  NOR2X1 G15760 (.A1(W9576), .A2(I299), .ZN(W27466));
  NOR2X1 G15761 (.A1(W5457), .A2(I1184), .ZN(W5698));
  NOR2X1 G15762 (.A1(W25542), .A2(W6804), .ZN(O15005));
  NOR2X1 G15763 (.A1(W5883), .A2(W20793), .ZN(O14543));
  NOR2X1 G15764 (.A1(W4255), .A2(W20445), .ZN(W23270));
  NOR2X1 G15765 (.A1(W30506), .A2(W43244), .ZN(O15007));
  NOR2X1 G15766 (.A1(W5624), .A2(W10411), .ZN(W23400));
  NOR2X1 G15767 (.A1(W23454), .A2(I196), .ZN(O14138));
  NOR2X1 G15768 (.A1(W4325), .A2(W703), .ZN(W5696));
  NOR2X1 G15769 (.A1(W15099), .A2(W385), .ZN(O2755));
  NOR2X1 G15770 (.A1(W7501), .A2(W793), .ZN(O3990));
  NOR2X1 G15771 (.A1(W29702), .A2(W19489), .ZN(O14135));
  NOR2X1 G15772 (.A1(W40911), .A2(W21716), .ZN(O14134));
  NOR2X1 G15773 (.A1(W20397), .A2(W33041), .ZN(O14130));
  NOR2X1 G15774 (.A1(W17924), .A2(W44225), .ZN(W44718));
  NOR2X1 G15775 (.A1(I519), .A2(I1253), .ZN(W5381));
  NOR2X1 G15776 (.A1(W3258), .A2(W2032), .ZN(W45119));
  NOR2X1 G15777 (.A1(W35711), .A2(W29283), .ZN(O14544));
  NOR2X1 G15778 (.A1(W32928), .A2(W36443), .ZN(O14545));
  NOR2X1 G15779 (.A1(I430), .A2(W2880), .ZN(W5501));
  NOR2X1 G15780 (.A1(W42346), .A2(W2644), .ZN(O14978));
  NOR2X1 G15781 (.A1(W1116), .A2(W17489), .ZN(W27122));
  NOR2X1 G15782 (.A1(W33856), .A2(W11403), .ZN(O14972));
  NOR2X1 G15783 (.A1(W4406), .A2(W506), .ZN(W5811));
  NOR2X1 G15784 (.A1(I82), .A2(W38043), .ZN(O14182));
  NOR2X1 G15785 (.A1(W4164), .A2(W11124), .ZN(W23606));
  NOR2X1 G15786 (.A1(W19764), .A2(W31235), .ZN(O14819));
  NOR2X1 G15787 (.A1(W19502), .A2(W22524), .ZN(W23433));
  NOR2X1 G15788 (.A1(W30180), .A2(W38226), .ZN(O14181));
  NOR2X1 G15789 (.A1(W25281), .A2(W31155), .ZN(O14180));
  NOR2X1 G15790 (.A1(W20453), .A2(W4291), .ZN(O14974));
  NOR2X1 G15791 (.A1(W5090), .A2(W2573), .ZN(W6150));
  NOR2X1 G15792 (.A1(W20175), .A2(W31624), .ZN(O14531));
  NOR2X1 G15793 (.A1(W5895), .A2(W3555), .ZN(W6155));
  NOR2X1 G15794 (.A1(I1388), .A2(W17042), .ZN(W23286));
  NOR2X1 G15795 (.A1(W31614), .A2(W18653), .ZN(O14980));
  NOR2X1 G15796 (.A1(W8358), .A2(W7585), .ZN(O14818));
  NOR2X1 G15797 (.A1(W1846), .A2(I1802), .ZN(W5200));
  NOR2X1 G15798 (.A1(I1790), .A2(W1004), .ZN(W6157));
  NOR2X1 G15799 (.A1(I1685), .A2(W4441), .ZN(W6158));
  NOR2X1 G15800 (.A1(W1154), .A2(W4488), .ZN(W5882));
  NOR2X1 G15801 (.A1(W16380), .A2(W11887), .ZN(O14964));
  NOR2X1 G15802 (.A1(W3327), .A2(W25852), .ZN(O14956));
  NOR2X1 G15803 (.A1(I1677), .A2(W3360), .ZN(W5371));
  NOR2X1 G15804 (.A1(W45078), .A2(I1554), .ZN(O14959));
  NOR2X1 G15805 (.A1(W39034), .A2(W14719), .ZN(O14961));
  NOR2X1 G15806 (.A1(W4706), .A2(W2289), .ZN(W5213));
  NOR2X1 G15807 (.A1(I756), .A2(W2954), .ZN(W5212));
  NOR2X1 G15808 (.A1(W3526), .A2(W191), .ZN(O14394));
  NOR2X1 G15809 (.A1(W3687), .A2(W1099), .ZN(W6146));
  NOR2X1 G15810 (.A1(W26648), .A2(W10492), .ZN(O14962));
  NOR2X1 G15811 (.A1(W4115), .A2(W6029), .ZN(W6147));
  NOR2X1 G15812 (.A1(W12349), .A2(W6743), .ZN(O2735));
  NOR2X1 G15813 (.A1(W15095), .A2(W43365), .ZN(O14965));
  NOR2X1 G15814 (.A1(W16570), .A2(W43437), .ZN(O14969));
  NOR2X1 G15815 (.A1(W41154), .A2(W3809), .ZN(W45124));
  NOR2X1 G15816 (.A1(W4974), .A2(W16088), .ZN(W27368));
  NOR2X1 G15817 (.A1(W3848), .A2(W1899), .ZN(W5715));
  NOR2X1 G15818 (.A1(W39906), .A2(W38794), .ZN(O14458));
  NOR2X1 G15819 (.A1(W5365), .A2(W5493), .ZN(W6148));
  NOR2X1 G15820 (.A1(W3664), .A2(W12559), .ZN(O14183));
  NOR2X1 G15821 (.A1(W20766), .A2(W23483), .ZN(W23604));
  NOR2X1 G15822 (.A1(W15880), .A2(W19119), .ZN(W23280));
  NOR2X1 G15823 (.A1(W1493), .A2(W4476), .ZN(W5377));
  NOR2X1 G15824 (.A1(W2878), .A2(W24993), .ZN(O14171));
  NOR2X1 G15825 (.A1(W1327), .A2(W5427), .ZN(W5495));
  NOR2X1 G15826 (.A1(I1456), .A2(W18527), .ZN(W23282));
  NOR2X1 G15827 (.A1(W18396), .A2(W1927), .ZN(O14168));
  NOR2X1 G15828 (.A1(W15863), .A2(W11008), .ZN(W23281));
  NOR2X1 G15829 (.A1(W27914), .A2(W35817), .ZN(W44765));
  NOR2X1 G15830 (.A1(W144), .A2(W12488), .ZN(W27119));
  NOR2X1 G15831 (.A1(W10419), .A2(W36061), .ZN(W45761));
  NOR2X1 G15832 (.A1(W3515), .A2(W3492), .ZN(W5193));
  NOR2X1 G15833 (.A1(W19137), .A2(W44181), .ZN(O14707));
  NOR2X1 G15834 (.A1(W37585), .A2(W42578), .ZN(O14165));
  NOR2X1 G15835 (.A1(W19332), .A2(W32114), .ZN(O14400));
  NOR2X1 G15836 (.A1(I212), .A2(W2957), .ZN(W5707));
  NOR2X1 G15837 (.A1(W4236), .A2(W4428), .ZN(W5706));
  NOR2X1 G15838 (.A1(W7823), .A2(W24755), .ZN(W27446));
  NOR2X1 G15839 (.A1(W3549), .A2(W2377), .ZN(W6178));
  NOR2X1 G15840 (.A1(W2927), .A2(W20643), .ZN(W27447));
  NOR2X1 G15841 (.A1(W16912), .A2(W19779), .ZN(O4108));
  NOR2X1 G15842 (.A1(W11373), .A2(W12824), .ZN(W23610));
  NOR2X1 G15843 (.A1(W15679), .A2(W9942), .ZN(W27367));
  NOR2X1 G15844 (.A1(W14878), .A2(W8020), .ZN(O14816));
  NOR2X1 G15845 (.A1(W43592), .A2(W8594), .ZN(O14176));
  NOR2X1 G15846 (.A1(W24576), .A2(W11898), .ZN(O14712));
  NOR2X1 G15847 (.A1(W481), .A2(W4467), .ZN(W6161));
  NOR2X1 G15848 (.A1(W23964), .A2(W2602), .ZN(O14981));
  NOR2X1 G15849 (.A1(W2424), .A2(W4452), .ZN(W5881));
  NOR2X1 G15850 (.A1(W43679), .A2(W25367), .ZN(O14982));
  NOR2X1 G15851 (.A1(W1276), .A2(W3678), .ZN(W6162));
  NOR2X1 G15852 (.A1(W5406), .A2(W209), .ZN(W6163));
  NOR2X1 G15853 (.A1(W20078), .A2(W37156), .ZN(O14174));
  NOR2X1 G15854 (.A1(W25520), .A2(W14768), .ZN(O4021));
  NOR2X1 G15855 (.A1(W1762), .A2(I1216), .ZN(W6165));
  NOR2X1 G15856 (.A1(W2573), .A2(I1904), .ZN(W6166));
  NOR2X1 G15857 (.A1(W12220), .A2(W26461), .ZN(W44775));
  NOR2X1 G15858 (.A1(W19921), .A2(I157), .ZN(W23435));
  NOR2X1 G15859 (.A1(W3692), .A2(I1484), .ZN(W5197));
  NOR2X1 G15860 (.A1(W4859), .A2(I30), .ZN(W5376));
  NOR2X1 G15861 (.A1(W4150), .A2(I486), .ZN(W5710));
  NOR2X1 G15862 (.A1(W42674), .A2(W5950), .ZN(O14709));
  NOR2X1 G15863 (.A1(W17123), .A2(W9508), .ZN(W23607));
  NOR2X1 G15864 (.A1(W1389), .A2(I889), .ZN(W5442));
  NOR2X1 G15865 (.A1(W2916), .A2(W5262), .ZN(W5970));
  NOR2X1 G15866 (.A1(W320), .A2(W17647), .ZN(W23344));
  NOR2X1 G15867 (.A1(W12390), .A2(W3391), .ZN(W27395));
  NOR2X1 G15868 (.A1(W12840), .A2(W4535), .ZN(W27396));
  NOR2X1 G15869 (.A1(W21716), .A2(W1070), .ZN(W27397));
  NOR2X1 G15870 (.A1(W15015), .A2(W5720), .ZN(W27382));
  NOR2X1 G15871 (.A1(W2983), .A2(W3505), .ZN(W5975));
  NOR2X1 G15872 (.A1(W2281), .A2(W528), .ZN(W5976));
  NOR2X1 G15873 (.A1(I1592), .A2(W17621), .ZN(W27399));
  NOR2X1 G15874 (.A1(W285), .A2(I1606), .ZN(W5351));
  NOR2X1 G15875 (.A1(W10995), .A2(W21774), .ZN(W27394));
  NOR2X1 G15876 (.A1(W9117), .A2(W38970), .ZN(O14362));
  NOR2X1 G15877 (.A1(W9648), .A2(W20858), .ZN(W23339));
  NOR2X1 G15878 (.A1(W5207), .A2(I1073), .ZN(W5979));
  NOR2X1 G15879 (.A1(W12673), .A2(W23997), .ZN(O14864));
  NOR2X1 G15880 (.A1(W16917), .A2(W1940), .ZN(W27211));
  NOR2X1 G15881 (.A1(I1486), .A2(W5451), .ZN(W5785));
  NOR2X1 G15882 (.A1(I181), .A2(W24597), .ZN(W27340));
  NOR2X1 G15883 (.A1(W700), .A2(W28392), .ZN(O14865));
  NOR2X1 G15884 (.A1(W6405), .A2(W2037), .ZN(W23338));
  NOR2X1 G15885 (.A1(W9978), .A2(W31599), .ZN(O14755));
  NOR2X1 G15886 (.A1(I1100), .A2(W3326), .ZN(W5319));
  NOR2X1 G15887 (.A1(W16852), .A2(W37128), .ZN(O14473));
  NOR2X1 G15888 (.A1(W2947), .A2(W1699), .ZN(W5324));
  NOR2X1 G15889 (.A1(W1109), .A2(W2107), .ZN(O100));
  NOR2X1 G15890 (.A1(W3423), .A2(W2385), .ZN(W5802));
  NOR2X1 G15891 (.A1(W33519), .A2(W37781), .ZN(O14359));
  NOR2X1 G15892 (.A1(W3864), .A2(W449), .ZN(W5323));
  NOR2X1 G15893 (.A1(W75), .A2(W3721), .ZN(W5321));
  NOR2X1 G15894 (.A1(W3699), .A2(I376), .ZN(W5320));
  NOR2X1 G15895 (.A1(W9332), .A2(W14069), .ZN(O2747));
  NOR2X1 G15896 (.A1(W4751), .A2(I794), .ZN(O101));
  NOR2X1 G15897 (.A1(W86), .A2(W3048), .ZN(W5782));
  NOR2X1 G15898 (.A1(W22727), .A2(W6058), .ZN(W23363));
  NOR2X1 G15899 (.A1(W7430), .A2(W22561), .ZN(O14859));
  NOR2X1 G15900 (.A1(W689), .A2(W4711), .ZN(W5317));
  NOR2X1 G15901 (.A1(W12038), .A2(W3691), .ZN(O2818));
  NOR2X1 G15902 (.A1(W4810), .A2(W4845), .ZN(W5919));
  NOR2X1 G15903 (.A1(W4074), .A2(I481), .ZN(W5966));
  NOR2X1 G15904 (.A1(W38634), .A2(W10266), .ZN(W45008));
  NOR2X1 G15905 (.A1(I905), .A2(I633), .ZN(O111));
  NOR2X1 G15906 (.A1(W1375), .A2(W19601), .ZN(O14316));
  NOR2X1 G15907 (.A1(W21029), .A2(W4952), .ZN(O14877));
  NOR2X1 G15908 (.A1(W5017), .A2(W2323), .ZN(W5777));
  NOR2X1 G15909 (.A1(W19426), .A2(W44516), .ZN(O14754));
  NOR2X1 G15910 (.A1(W5859), .A2(W1595), .ZN(W5993));
  NOR2X1 G15911 (.A1(W10421), .A2(W23621), .ZN(W27332));
  NOR2X1 G15912 (.A1(W25163), .A2(W1319), .ZN(O14872));
  NOR2X1 G15913 (.A1(W19770), .A2(W4236), .ZN(W23555));
  NOR2X1 G15914 (.A1(I308), .A2(W215), .ZN(W5353));
  NOR2X1 G15915 (.A1(W5031), .A2(W32166), .ZN(O14304));
  NOR2X1 G15916 (.A1(W15458), .A2(W40404), .ZN(O14366));
  NOR2X1 G15917 (.A1(W39216), .A2(W26872), .ZN(O14835));
  NOR2X1 G15918 (.A1(W5546), .A2(W5749), .ZN(W5992));
  NOR2X1 G15919 (.A1(W1714), .A2(W5143), .ZN(W5303));
  NOR2X1 G15920 (.A1(W10958), .A2(W28496), .ZN(O14301));
  NOR2X1 G15921 (.A1(I522), .A2(W454), .ZN(O115));
  NOR2X1 G15922 (.A1(W19414), .A2(W4342), .ZN(O14300));
  NOR2X1 G15923 (.A1(W3180), .A2(W10255), .ZN(O14878));
  NOR2X1 G15924 (.A1(W271), .A2(W423), .ZN(W6000));
  NOR2X1 G15925 (.A1(I1435), .A2(I1497), .ZN(W5301));
  NOR2X1 G15926 (.A1(W4394), .A2(W2627), .ZN(W5428));
  NOR2X1 G15927 (.A1(I629), .A2(W862), .ZN(W5449));
  NOR2X1 G15928 (.A1(W1152), .A2(I494), .ZN(W5308));
  NOR2X1 G15929 (.A1(W22882), .A2(W24673), .ZN(O14868));
  NOR2X1 G15930 (.A1(W1630), .A2(W1557), .ZN(W5981));
  NOR2X1 G15931 (.A1(W5023), .A2(W2149), .ZN(W5915));
  NOR2X1 G15932 (.A1(W2093), .A2(W11986), .ZN(O14476));
  NOR2X1 G15933 (.A1(W1180), .A2(I294), .ZN(W5982));
  NOR2X1 G15934 (.A1(W27086), .A2(W15305), .ZN(O4085));
  NOR2X1 G15935 (.A1(I392), .A2(W4304), .ZN(W5984));
  NOR2X1 G15936 (.A1(W797), .A2(W3541), .ZN(W5985));
  NOR2X1 G15937 (.A1(W964), .A2(W5773), .ZN(W23336));
  NOR2X1 G15938 (.A1(W15479), .A2(W2387), .ZN(W23570));
  NOR2X1 G15939 (.A1(W23282), .A2(W6949), .ZN(W27393));
  NOR2X1 G15940 (.A1(W1254), .A2(W28786), .ZN(O14477));
  NOR2X1 G15941 (.A1(W2688), .A2(I712), .ZN(W5988));
  NOR2X1 G15942 (.A1(I152), .A2(W2581), .ZN(W5989));
  NOR2X1 G15943 (.A1(W2367), .A2(W1589), .ZN(W5990));
  NOR2X1 G15944 (.A1(W3319), .A2(W5413), .ZN(W5445));
  NOR2X1 G15945 (.A1(W3788), .A2(W5891), .ZN(W5991));
  NOR2X1 G15946 (.A1(W24925), .A2(W7878), .ZN(O14478));
  NOR2X1 G15947 (.A1(I235), .A2(W277), .ZN(W5307));
  NOR2X1 G15948 (.A1(W3778), .A2(W1424), .ZN(W5446));
  NOR2X1 G15949 (.A1(W20649), .A2(W22668), .ZN(W45594));
  NOR2X1 G15950 (.A1(W2963), .A2(W17152), .ZN(W23354));
  NOR2X1 G15951 (.A1(W21040), .A2(W839), .ZN(W23559));
  NOR2X1 G15952 (.A1(W3958), .A2(W4670), .ZN(W5343));
  NOR2X1 G15953 (.A1(W26035), .A2(W10568), .ZN(O14348));
  NOR2X1 G15954 (.A1(W19611), .A2(W10471), .ZN(W23353));
  NOR2X1 G15955 (.A1(I688), .A2(W5246), .ZN(W5342));
  NOR2X1 G15956 (.A1(I1448), .A2(W1539), .ZN(W5943));
  NOR2X1 G15957 (.A1(I1104), .A2(W1978), .ZN(W5341));
  NOR2X1 G15958 (.A1(W34639), .A2(W29989), .ZN(W44998));
  NOR2X1 G15959 (.A1(W7394), .A2(W16540), .ZN(W23405));
  NOR2X1 G15960 (.A1(W35353), .A2(W41128), .ZN(O14767));
  NOR2X1 G15961 (.A1(I798), .A2(W1883), .ZN(W5339));
  NOR2X1 G15962 (.A1(W3395), .A2(W40158), .ZN(O14344));
  NOR2X1 G15963 (.A1(W10205), .A2(W14547), .ZN(O14343));
  NOR2X1 G15964 (.A1(W14594), .A2(W15126), .ZN(O14341));
  NOR2X1 G15965 (.A1(W3539), .A2(W1424), .ZN(W5947));
  NOR2X1 G15966 (.A1(W227), .A2(W5132), .ZN(W5434));
  NOR2X1 G15967 (.A1(W3863), .A2(W496), .ZN(W5435));
  NOR2X1 G15968 (.A1(I725), .A2(I255), .ZN(W5796));
  NOR2X1 G15969 (.A1(W7684), .A2(W41036), .ZN(O14768));
  NOR2X1 G15970 (.A1(W10003), .A2(W14420), .ZN(W27346));
  NOR2X1 G15971 (.A1(W885), .A2(W1729), .ZN(W5927));
  NOR2X1 G15972 (.A1(W1578), .A2(I13), .ZN(W5801));
  NOR2X1 G15973 (.A1(W14874), .A2(W31133), .ZN(O14766));
  NOR2X1 G15974 (.A1(W22969), .A2(W3896), .ZN(O4088));
  NOR2X1 G15975 (.A1(W389), .A2(W2290), .ZN(W5929));
  NOR2X1 G15976 (.A1(W5832), .A2(W44187), .ZN(W44996));
  NOR2X1 G15977 (.A1(W308), .A2(W3023), .ZN(W5349));
  NOR2X1 G15978 (.A1(W16569), .A2(W10553), .ZN(W23358));
  NOR2X1 G15979 (.A1(W4626), .A2(W1720), .ZN(W5933));
  NOR2X1 G15980 (.A1(W40536), .A2(W29546), .ZN(W44993));
  NOR2X1 G15981 (.A1(W12792), .A2(W35145), .ZN(O14340));
  NOR2X1 G15982 (.A1(W33989), .A2(W26118), .ZN(O14838));
  NOR2X1 G15983 (.A1(W9229), .A2(W6476), .ZN(W23357));
  NOR2X1 G15984 (.A1(I559), .A2(W4152), .ZN(W5346));
  NOR2X1 G15985 (.A1(W43813), .A2(W4469), .ZN(O14349));
  NOR2X1 G15986 (.A1(W2439), .A2(W4197), .ZN(W5432));
  NOR2X1 G15987 (.A1(W6081), .A2(W2846), .ZN(W23356));
  NOR2X1 G15988 (.A1(I725), .A2(I950), .ZN(W5798));
  NOR2X1 G15989 (.A1(W11716), .A2(W18933), .ZN(W27389));
  NOR2X1 G15990 (.A1(W5622), .A2(W1671), .ZN(W5939));
  NOR2X1 G15991 (.A1(W843), .A2(I1575), .ZN(W5441));
  NOR2X1 G15992 (.A1(I870), .A2(I499), .ZN(W5958));
  NOR2X1 G15993 (.A1(W5447), .A2(W4248), .ZN(W5923));
  NOR2X1 G15994 (.A1(W39590), .A2(W8124), .ZN(O14469));
  NOR2X1 G15995 (.A1(W2433), .A2(W4498), .ZN(W5330));
  NOR2X1 G15996 (.A1(W1446), .A2(W2312), .ZN(O4009));
  NOR2X1 G15997 (.A1(I825), .A2(I1651), .ZN(W5791));
  NOR2X1 G15998 (.A1(I1353), .A2(W1602), .ZN(W5328));
  NOR2X1 G15999 (.A1(W25402), .A2(W36485), .ZN(O14327));
  NOR2X1 G16000 (.A1(W35096), .A2(W29003), .ZN(O14759));
  NOR2X1 G16001 (.A1(W13609), .A2(W26063), .ZN(O4024));
  NOR2X1 G16002 (.A1(W12879), .A2(W38495), .ZN(O14330));
  NOR2X1 G16003 (.A1(W19558), .A2(W13706), .ZN(O14857));
  NOR2X1 G16004 (.A1(W1534), .A2(W11447), .ZN(O4069));
  NOR2X1 G16005 (.A1(W32778), .A2(W15231), .ZN(O14324));
  NOR2X1 G16006 (.A1(W10929), .A2(W5011), .ZN(W27383));
  NOR2X1 G16007 (.A1(W302), .A2(W3804), .ZN(W5789));
  NOR2X1 G16008 (.A1(W895), .A2(I7), .ZN(W5788));
  NOR2X1 G16009 (.A1(W27812), .A2(W11450), .ZN(O14322));
  NOR2X1 G16010 (.A1(I1444), .A2(W941), .ZN(W5325));
  NOR2X1 G16011 (.A1(W15757), .A2(I499), .ZN(W23348));
  NOR2X1 G16012 (.A1(W39154), .A2(W20065), .ZN(O14852));
  NOR2X1 G16013 (.A1(I1660), .A2(I636), .ZN(W5949));
  NOR2X1 G16014 (.A1(W7958), .A2(W25751), .ZN(O4072));
  NOR2X1 G16015 (.A1(W41749), .A2(W21684), .ZN(W44976));
  NOR2X1 G16016 (.A1(W15514), .A2(W38116), .ZN(O14845));
  NOR2X1 G16017 (.A1(W23199), .A2(W3285), .ZN(W27391));
  NOR2X1 G16018 (.A1(W2250), .A2(I1388), .ZN(W5952));
  NOR2X1 G16019 (.A1(W22464), .A2(W17371), .ZN(O2816));
  NOR2X1 G16020 (.A1(W1214), .A2(W2599), .ZN(W5334));
  NOR2X1 G16021 (.A1(W1934), .A2(W11412), .ZN(W23407));
  NOR2X1 G16022 (.A1(W10450), .A2(W19104), .ZN(O14335));
  NOR2X1 G16023 (.A1(W3672), .A2(W377), .ZN(W6001));
  NOR2X1 G16024 (.A1(W14703), .A2(W32476), .ZN(O14334));
  NOR2X1 G16025 (.A1(W41302), .A2(W27222), .ZN(O14354));
  NOR2X1 G16026 (.A1(W1757), .A2(W3821), .ZN(O82));
  NOR2X1 G16027 (.A1(W17580), .A2(W9274), .ZN(O14853));
  NOR2X1 G16028 (.A1(W25331), .A2(W6123), .ZN(W27206));
  NOR2X1 G16029 (.A1(W19782), .A2(W22837), .ZN(W23351));
  NOR2X1 G16030 (.A1(W12231), .A2(W24140), .ZN(W27208));
  NOR2X1 G16031 (.A1(W12860), .A2(W17494), .ZN(W23361));
  NOR2X1 G16032 (.A1(W3304), .A2(W970), .ZN(W23350));
  NOR2X1 G16033 (.A1(W632), .A2(W5416), .ZN(W5905));
  NOR2X1 G16034 (.A1(W4102), .A2(W5023), .ZN(W5360));
  NOR2X1 G16035 (.A1(I1518), .A2(W754), .ZN(W6052));
  NOR2X1 G16036 (.A1(W19249), .A2(W4178), .ZN(O14492));
  NOR2X1 G16037 (.A1(W42454), .A2(W30856), .ZN(O14772));
  NOR2X1 G16038 (.A1(W5153), .A2(W21756), .ZN(O14901));
  NOR2X1 G16039 (.A1(I1402), .A2(W9405), .ZN(O14902));
  NOR2X1 G16040 (.A1(I884), .A2(W713), .ZN(W6054));
  NOR2X1 G16041 (.A1(W2845), .A2(W401), .ZN(W5275));
  NOR2X1 G16042 (.A1(I1036), .A2(W2744), .ZN(W5274));
  NOR2X1 G16043 (.A1(W2432), .A2(W2288), .ZN(W6055));
  NOR2X1 G16044 (.A1(W37197), .A2(W32309), .ZN(W45161));
  NOR2X1 G16045 (.A1(W13239), .A2(W16185), .ZN(W23551));
  NOR2X1 G16046 (.A1(W21595), .A2(W26154), .ZN(O14493));
  NOR2X1 G16047 (.A1(I1998), .A2(W42989), .ZN(O14495));
  NOR2X1 G16048 (.A1(W26023), .A2(W15497), .ZN(O3996));
  NOR2X1 G16049 (.A1(W4687), .A2(W19909), .ZN(O14496));
  NOR2X1 G16050 (.A1(W258), .A2(W26247), .ZN(W27219));
  NOR2X1 G16051 (.A1(W21712), .A2(W17221), .ZN(O3995));
  NOR2X1 G16052 (.A1(W2916), .A2(W593), .ZN(W5462));
  NOR2X1 G16053 (.A1(W2447), .A2(W366), .ZN(W5904));
  NOR2X1 G16054 (.A1(W810), .A2(W1251), .ZN(W6047));
  NOR2X1 G16055 (.A1(W11427), .A2(W44312), .ZN(O14898));
  NOR2X1 G16056 (.A1(W16628), .A2(W21448), .ZN(W23519));
  NOR2X1 G16057 (.A1(W41561), .A2(W42322), .ZN(O14269));
  NOR2X1 G16058 (.A1(W1078), .A2(W2098), .ZN(W27417));
  NOR2X1 G16059 (.A1(W26973), .A2(W25369), .ZN(O14266));
  NOR2X1 G16060 (.A1(W4262), .A2(W6203), .ZN(W23418));
  NOR2X1 G16061 (.A1(W22872), .A2(W16913), .ZN(O4001));
  NOR2X1 G16062 (.A1(W31424), .A2(W9029), .ZN(O14491));
  NOR2X1 G16063 (.A1(W24), .A2(I388), .ZN(O79));
  NOR2X1 G16064 (.A1(W5682), .A2(W906), .ZN(W6046));
  NOR2X1 G16065 (.A1(W22100), .A2(W16479), .ZN(O14253));
  NOR2X1 G16066 (.A1(W23007), .A2(W7004), .ZN(W23552));
  NOR2X1 G16067 (.A1(W1987), .A2(W2497), .ZN(W5280));
  NOR2X1 G16068 (.A1(W19617), .A2(W21371), .ZN(O14900));
  NOR2X1 G16069 (.A1(W11277), .A2(W21230), .ZN(W23317));
  NOR2X1 G16070 (.A1(W40792), .A2(W26853), .ZN(W45467));
  NOR2X1 G16071 (.A1(W44836), .A2(W11670), .ZN(W44882));
  NOR2X1 G16072 (.A1(I893), .A2(W3410), .ZN(W6050));
  NOR2X1 G16073 (.A1(W13269), .A2(W18991), .ZN(O14260));
  NOR2X1 G16074 (.A1(W995), .A2(I1819), .ZN(W5278));
  NOR2X1 G16075 (.A1(W7246), .A2(W15978), .ZN(O14919));
  NOR2X1 G16076 (.A1(W3973), .A2(I1606), .ZN(O117));
  NOR2X1 G16077 (.A1(W13043), .A2(W5410), .ZN(W27139));
  NOR2X1 G16078 (.A1(W19340), .A2(W14583), .ZN(O14912));
  NOR2X1 G16079 (.A1(W16546), .A2(W6420), .ZN(W23587));
  NOR2X1 G16080 (.A1(W30883), .A2(W18170), .ZN(W45674));
  NOR2X1 G16081 (.A1(W3869), .A2(W3792), .ZN(W5750));
  NOR2X1 G16082 (.A1(W93), .A2(I836), .ZN(W5749));
  NOR2X1 G16083 (.A1(W3046), .A2(W4757), .ZN(W5258));
  NOR2X1 G16084 (.A1(W27613), .A2(W37926), .ZN(O14916));
  NOR2X1 G16085 (.A1(W10457), .A2(W1999), .ZN(W27138));
  NOR2X1 G16086 (.A1(W28719), .A2(W4293), .ZN(O14244));
  NOR2X1 G16087 (.A1(W1716), .A2(W2092), .ZN(W5254));
  NOR2X1 G16088 (.A1(W1589), .A2(W242), .ZN(W5253));
  NOR2X1 G16089 (.A1(W23036), .A2(W19987), .ZN(W23309));
  NOR2X1 G16090 (.A1(I1243), .A2(I1280), .ZN(W5748));
  NOR2X1 G16091 (.A1(W32537), .A2(W13963), .ZN(O14736));
  NOR2X1 G16092 (.A1(W9387), .A2(W18740), .ZN(O14920));
  NOR2X1 G16093 (.A1(I1888), .A2(W2012), .ZN(W5747));
  NOR2X1 G16094 (.A1(W5139), .A2(W3119), .ZN(W5746));
  NOR2X1 G16095 (.A1(W5238), .A2(W362), .ZN(W5901));
  NOR2X1 G16096 (.A1(W5168), .A2(W14799), .ZN(O2820));
  NOR2X1 G16097 (.A1(W4877), .A2(W30431), .ZN(W45025));
  NOR2X1 G16098 (.A1(I416), .A2(I444), .ZN(W5269));
  NOR2X1 G16099 (.A1(W20613), .A2(W35510), .ZN(O14907));
  NOR2X1 G16100 (.A1(W3392), .A2(W7329), .ZN(O2768));
  NOR2X1 G16101 (.A1(W3331), .A2(W5138), .ZN(W5267));
  NOR2X1 G16102 (.A1(W2019), .A2(W85), .ZN(W6059));
  NOR2X1 G16103 (.A1(W9544), .A2(W30436), .ZN(O14251));
  NOR2X1 G16104 (.A1(I468), .A2(W2864), .ZN(W6061));
  NOR2X1 G16105 (.A1(W2007), .A2(W1392), .ZN(W6062));
  NOR2X1 G16106 (.A1(W25930), .A2(W34439), .ZN(O14908));
  NOR2X1 G16107 (.A1(W22765), .A2(W11845), .ZN(O4097));
  NOR2X1 G16108 (.A1(W9718), .A2(W35144), .ZN(O14248));
  NOR2X1 G16109 (.A1(W16160), .A2(W743), .ZN(W27422));
  NOR2X1 G16110 (.A1(I100), .A2(W5182), .ZN(W5264));
  NOR2X1 G16111 (.A1(W10870), .A2(W4001), .ZN(O4100));
  NOR2X1 G16112 (.A1(W13024), .A2(W16074), .ZN(W27140));
  NOR2X1 G16113 (.A1(W4904), .A2(W7954), .ZN(W23371));
  NOR2X1 G16114 (.A1(W38721), .A2(W19243), .ZN(O14738));
  NOR2X1 G16115 (.A1(W22809), .A2(W9025), .ZN(O2740));
  NOR2X1 G16116 (.A1(W23694), .A2(W11061), .ZN(W27221));
  NOR2X1 G16117 (.A1(W13135), .A2(W16767), .ZN(O2743));
  NOR2X1 G16118 (.A1(W31223), .A2(W13489), .ZN(O14884));
  NOR2X1 G16119 (.A1(I584), .A2(I422), .ZN(W5295));
  NOR2X1 G16120 (.A1(I309), .A2(W1287), .ZN(W5770));
  NOR2X1 G16121 (.A1(W1415), .A2(W2373), .ZN(W5452));
  NOR2X1 G16122 (.A1(W21203), .A2(W16362), .ZN(W45641));
  NOR2X1 G16123 (.A1(W4912), .A2(I196), .ZN(W5768));
  NOR2X1 G16124 (.A1(I1892), .A2(I1464), .ZN(W5358));
  NOR2X1 G16125 (.A1(I1541), .A2(W17750), .ZN(W23328));
  NOR2X1 G16126 (.A1(W7341), .A2(W9845), .ZN(W23575));
  NOR2X1 G16127 (.A1(W21947), .A2(W766), .ZN(W23326));
  NOR2X1 G16128 (.A1(W2172), .A2(W12835), .ZN(O2744));
  NOR2X1 G16129 (.A1(W2133), .A2(W41375), .ZN(O14290));
  NOR2X1 G16130 (.A1(W12105), .A2(W13950), .ZN(W23324));
  NOR2X1 G16131 (.A1(I968), .A2(W270), .ZN(O14285));
  NOR2X1 G16132 (.A1(W4834), .A2(W3663), .ZN(W5292));
  NOR2X1 G16133 (.A1(W38622), .A2(W3931), .ZN(O14746));
  NOR2X1 G16134 (.A1(W1801), .A2(I1794), .ZN(W5767));
  NOR2X1 G16135 (.A1(W4357), .A2(I200), .ZN(W6018));
  NOR2X1 G16136 (.A1(W28313), .A2(W27540), .ZN(O14284));
  NOR2X1 G16137 (.A1(W9286), .A2(W13691), .ZN(O14283));
  NOR2X1 G16138 (.A1(W173), .A2(W2565), .ZN(W6005));
  NOR2X1 G16139 (.A1(W26702), .A2(W9822), .ZN(O14881));
  NOR2X1 G16140 (.A1(W13774), .A2(W11724), .ZN(O14369));
  NOR2X1 G16141 (.A1(W6055), .A2(W13380), .ZN(O4004));
  NOR2X1 G16142 (.A1(I889), .A2(W976), .ZN(W5356));
  NOR2X1 G16143 (.A1(W8184), .A2(W22023), .ZN(W23332));
  NOR2X1 G16144 (.A1(W31170), .A2(W41905), .ZN(O14481));
  NOR2X1 G16145 (.A1(W32888), .A2(W1925), .ZN(O14482));
  NOR2X1 G16146 (.A1(W6201), .A2(W12995), .ZN(W23553));
  NOR2X1 G16147 (.A1(W10324), .A2(W2243), .ZN(W23415));
  NOR2X1 G16148 (.A1(W38218), .A2(W27610), .ZN(O14297));
  NOR2X1 G16149 (.A1(W22928), .A2(W42107), .ZN(O14282));
  NOR2X1 G16150 (.A1(I1648), .A2(W13748), .ZN(O4095));
  NOR2X1 G16151 (.A1(W31554), .A2(W28967), .ZN(O14295));
  NOR2X1 G16152 (.A1(W1436), .A2(W2814), .ZN(W5771));
  NOR2X1 G16153 (.A1(W18710), .A2(W12556), .ZN(W23524));
  NOR2X1 G16154 (.A1(W2704), .A2(W4883), .ZN(W6008));
  NOR2X1 G16155 (.A1(W1048), .A2(W12138), .ZN(W27153));
  NOR2X1 G16156 (.A1(W3663), .A2(W2995), .ZN(W23574));
  NOR2X1 G16157 (.A1(W5830), .A2(W725), .ZN(O116));
  NOR2X1 G16158 (.A1(W12840), .A2(W7002), .ZN(O14748));
  NOR2X1 G16159 (.A1(W21979), .A2(W3687), .ZN(W27415));
  NOR2X1 G16160 (.A1(W14992), .A2(W37700), .ZN(W44902));
  NOR2X1 G16161 (.A1(W5986), .A2(W4320), .ZN(W6034));
  NOR2X1 G16162 (.A1(W35889), .A2(W8562), .ZN(O14277));
  NOR2X1 G16163 (.A1(W43541), .A2(W18369), .ZN(O14891));
  NOR2X1 G16164 (.A1(W29715), .A2(W6262), .ZN(O14276));
  NOR2X1 G16165 (.A1(W4203), .A2(W4107), .ZN(O99));
  NOR2X1 G16166 (.A1(W26288), .A2(W16), .ZN(O4074));
  NOR2X1 G16167 (.A1(I243), .A2(W41486), .ZN(W45470));
  NOR2X1 G16168 (.A1(W21264), .A2(W23149), .ZN(W27326));
  NOR2X1 G16169 (.A1(W38754), .A2(W40100), .ZN(O14488));
  NOR2X1 G16170 (.A1(W11323), .A2(W34488), .ZN(W45500));
  NOR2X1 G16171 (.A1(W9538), .A2(W24523), .ZN(O4002));
  NOR2X1 G16172 (.A1(W27727), .A2(W9716), .ZN(O14371));
  NOR2X1 G16173 (.A1(I1132), .A2(W4571), .ZN(W5760));
  NOR2X1 G16174 (.A1(W4867), .A2(W22819), .ZN(W23369));
  NOR2X1 G16175 (.A1(W3468), .A2(W18204), .ZN(W23320));
  NOR2X1 G16176 (.A1(W4017), .A2(W36), .ZN(W44895));
  NOR2X1 G16177 (.A1(W18791), .A2(W32035), .ZN(O14272));
  NOR2X1 G16178 (.A1(W1172), .A2(W22023), .ZN(W27218));
  NOR2X1 G16179 (.A1(W40196), .A2(W2484), .ZN(O14271));
  NOR2X1 G16180 (.A1(W40340), .A2(W29958), .ZN(W44907));
  NOR2X1 G16181 (.A1(W350), .A2(W4034), .ZN(W5766));
  NOR2X1 G16182 (.A1(W11394), .A2(W16842), .ZN(O4027));
  NOR2X1 G16183 (.A1(W5732), .A2(W10050), .ZN(W23323));
  NOR2X1 G16184 (.A1(W15650), .A2(W29727), .ZN(O14888));
  NOR2X1 G16185 (.A1(W6061), .A2(W4182), .ZN(W23368));
  NOR2X1 G16186 (.A1(W1675), .A2(W12288), .ZN(W23322));
  NOR2X1 G16187 (.A1(W688), .A2(W4969), .ZN(W5289));
  NOR2X1 G16188 (.A1(W4017), .A2(W12598), .ZN(W44908));
  NOR2X1 G16189 (.A1(W2466), .A2(I1955), .ZN(W5288));
  NOR2X1 G16190 (.A1(W3251), .A2(I296), .ZN(W6025));
  NOR2X1 G16191 (.A1(I810), .A2(W23354), .ZN(W23623));
  NOR2X1 G16192 (.A1(W3132), .A2(I66), .ZN(W6027));
  NOR2X1 G16193 (.A1(W38537), .A2(W43884), .ZN(O14279));
  NOR2X1 G16194 (.A1(I1546), .A2(W3445), .ZN(W5765));
  NOR2X1 G16195 (.A1(W35799), .A2(W25170), .ZN(O14486));
  NOR2X1 G16196 (.A1(W26599), .A2(W41870), .ZN(O14278));
  NOR2X1 G16197 (.A1(W33703), .A2(W8427), .ZN(O14889));
  NOR2X1 G16198 (.A1(W2860), .A2(W2865), .ZN(W6030));
  NOR2X1 G16199 (.A1(W12131), .A2(W40538), .ZN(W44904));
  NOR2X1 G16200 (.A1(W42658), .A2(W44501), .ZN(W44903));
  NOR2X1 G16201 (.A1(W1165), .A2(I1935), .ZN(W6402));
  NOR2X1 G16202 (.A1(W41069), .A2(W16991), .ZN(O13969));
  NOR2X1 G16203 (.A1(W3518), .A2(W4975), .ZN(W5603));
  NOR2X1 G16204 (.A1(W41349), .A2(W1029), .ZN(O15103));
  NOR2X1 G16205 (.A1(W589), .A2(W1052), .ZN(W5052));
  NOR2X1 G16206 (.A1(W3308), .A2(W6269), .ZN(W6400));
  NOR2X1 G16207 (.A1(W7012), .A2(W9232), .ZN(W27253));
  NOR2X1 G16208 (.A1(W613), .A2(I1425), .ZN(W5844));
  NOR2X1 G16209 (.A1(I640), .A2(W1138), .ZN(W5051));
  NOR2X1 G16210 (.A1(W29675), .A2(W39398), .ZN(O14613));
  NOR2X1 G16211 (.A1(W32653), .A2(W36016), .ZN(W44516));
  NOR2X1 G16212 (.A1(W15494), .A2(W3687), .ZN(W27279));
  NOR2X1 G16213 (.A1(W2146), .A2(W497), .ZN(W6403));
  NOR2X1 G16214 (.A1(W4784), .A2(W5826), .ZN(W5843));
  NOR2X1 G16215 (.A1(I1361), .A2(W3244), .ZN(W5050));
  NOR2X1 G16216 (.A1(W42950), .A2(I91), .ZN(O14435));
  NOR2X1 G16217 (.A1(W41548), .A2(W19247), .ZN(O13965));
  NOR2X1 G16218 (.A1(W19780), .A2(W6560), .ZN(W23660));
  NOR2X1 G16219 (.A1(W20448), .A2(W31955), .ZN(O15104));
  NOR2X1 G16220 (.A1(W19315), .A2(W15240), .ZN(W23485));
  NOR2X1 G16221 (.A1(I969), .A2(W1663), .ZN(O13964));
  NOR2X1 G16222 (.A1(W14136), .A2(W14762), .ZN(W27528));
  NOR2X1 G16223 (.A1(W16655), .A2(W4362), .ZN(O14609));
  NOR2X1 G16224 (.A1(W12360), .A2(W37588), .ZN(O14799));
  NOR2X1 G16225 (.A1(W3757), .A2(W1365), .ZN(W5845));
  NOR2X1 G16226 (.A1(W2290), .A2(W2663), .ZN(W5540));
  NOR2X1 G16227 (.A1(W2994), .A2(W3072), .ZN(W5541));
  NOR2X1 G16228 (.A1(I42), .A2(W3126), .ZN(W5825));
  NOR2X1 G16229 (.A1(W1602), .A2(I638), .ZN(O73));
  NOR2X1 G16230 (.A1(W32755), .A2(W6124), .ZN(O15100));
  NOR2X1 G16231 (.A1(W4249), .A2(W3206), .ZN(W6391));
  NOR2X1 G16232 (.A1(W4001), .A2(I693), .ZN(W6392));
  NOR2X1 G16233 (.A1(I441), .A2(W2517), .ZN(W5047));
  NOR2X1 G16234 (.A1(W4946), .A2(W1137), .ZN(W5413));
  NOR2X1 G16235 (.A1(W4254), .A2(W1862), .ZN(W6394));
  NOR2X1 G16236 (.A1(I548), .A2(W2303), .ZN(W6395));
  NOR2X1 G16237 (.A1(W5011), .A2(I1523), .ZN(W6396));
  NOR2X1 G16238 (.A1(W6875), .A2(W22340), .ZN(O4014));
  NOR2X1 G16239 (.A1(W32970), .A2(W7346), .ZN(O14610));
  NOR2X1 G16240 (.A1(W916), .A2(W15811), .ZN(W23205));
  NOR2X1 G16241 (.A1(W26962), .A2(W33608), .ZN(O13972));
  NOR2X1 G16242 (.A1(W156), .A2(W5407), .ZN(W5542));
  NOR2X1 G16243 (.A1(W660), .A2(W1710), .ZN(W5547));
  NOR2X1 G16244 (.A1(W1527), .A2(W5119), .ZN(W6423));
  NOR2X1 G16245 (.A1(W29852), .A2(W17914), .ZN(O13947));
  NOR2X1 G16246 (.A1(W4543), .A2(W2347), .ZN(W5546));
  NOR2X1 G16247 (.A1(W3579), .A2(W4906), .ZN(W5043));
  NOR2X1 G16248 (.A1(W4308), .A2(W22489), .ZN(O3973));
  NOR2X1 G16249 (.A1(W772), .A2(W2666), .ZN(W5041));
  NOR2X1 G16250 (.A1(I375), .A2(I929), .ZN(W6425));
  NOR2X1 G16251 (.A1(W7797), .A2(W13076), .ZN(W27062));
  NOR2X1 G16252 (.A1(W41233), .A2(W31628), .ZN(W45314));
  NOR2X1 G16253 (.A1(W35758), .A2(W26031), .ZN(O13946));
  NOR2X1 G16254 (.A1(W29678), .A2(W44305), .ZN(O13948));
  NOR2X1 G16255 (.A1(I1507), .A2(W2395), .ZN(W5841));
  NOR2X1 G16256 (.A1(W1999), .A2(W4588), .ZN(O131));
  NOR2X1 G16257 (.A1(W33408), .A2(W31159), .ZN(O14616));
  NOR2X1 G16258 (.A1(W469), .A2(W3822), .ZN(W5038));
  NOR2X1 G16259 (.A1(W5642), .A2(W932), .ZN(W6428));
  NOR2X1 G16260 (.A1(W5754), .A2(I242), .ZN(W5840));
  NOR2X1 G16261 (.A1(W1895), .A2(W15436), .ZN(W27274));
  NOR2X1 G16262 (.A1(W2265), .A2(W3140), .ZN(W5400));
  NOR2X1 G16263 (.A1(I877), .A2(W2673), .ZN(W5037));
  NOR2X1 G16264 (.A1(W23251), .A2(W30761), .ZN(O15107));
  NOR2X1 G16265 (.A1(W36746), .A2(W28807), .ZN(O13962));
  NOR2X1 G16266 (.A1(I1095), .A2(W3900), .ZN(W6408));
  NOR2X1 G16267 (.A1(W2997), .A2(W10015), .ZN(O4140));
  NOR2X1 G16268 (.A1(W3602), .A2(W2357), .ZN(W6410));
  NOR2X1 G16269 (.A1(W26457), .A2(W42782), .ZN(O13959));
  NOR2X1 G16270 (.A1(W6419), .A2(W4986), .ZN(W45532));
  NOR2X1 G16271 (.A1(W12545), .A2(W13516), .ZN(W23202));
  NOR2X1 G16272 (.A1(W30260), .A2(W300), .ZN(O14614));
  NOR2X1 G16273 (.A1(W8221), .A2(W16655), .ZN(W23201));
  NOR2X1 G16274 (.A1(W21621), .A2(W21583), .ZN(O2706));
  NOR2X1 G16275 (.A1(W43128), .A2(W4507), .ZN(O14434));
  NOR2X1 G16276 (.A1(W38487), .A2(W24409), .ZN(O14661));
  NOR2X1 G16277 (.A1(W22781), .A2(W18758), .ZN(O13955));
  NOR2X1 G16278 (.A1(W42989), .A2(W21202), .ZN(O13953));
  NOR2X1 G16279 (.A1(W15917), .A2(W22047), .ZN(W27067));
  NOR2X1 G16280 (.A1(I464), .A2(W20405), .ZN(W27534));
  NOR2X1 G16281 (.A1(W5317), .A2(W1189), .ZN(W6418));
  NOR2X1 G16282 (.A1(W26560), .A2(W31830), .ZN(O13952));
  NOR2X1 G16283 (.A1(W41889), .A2(W2104), .ZN(O13950));
  NOR2X1 G16284 (.A1(I122), .A2(W4456), .ZN(O2705));
  NOR2X1 G16285 (.A1(W33994), .A2(W33908), .ZN(W45299));
  NOR2X1 G16286 (.A1(W2021), .A2(W4585), .ZN(W6366));
  NOR2X1 G16287 (.A1(W5265), .A2(W2056), .ZN(W5620));
  NOR2X1 G16288 (.A1(W1839), .A2(W6522), .ZN(W23213));
  NOR2X1 G16289 (.A1(I1448), .A2(W2085), .ZN(W5072));
  NOR2X1 G16290 (.A1(W37540), .A2(W5627), .ZN(O14600));
  NOR2X1 G16291 (.A1(W2322), .A2(W2184), .ZN(W5071));
  NOR2X1 G16292 (.A1(W16667), .A2(W31699), .ZN(W44548));
  NOR2X1 G16293 (.A1(W26776), .A2(W4472), .ZN(O13993));
  NOR2X1 G16294 (.A1(W5058), .A2(W1008), .ZN(W6370));
  NOR2X1 G16295 (.A1(W17596), .A2(W18007), .ZN(W44542));
  NOR2X1 G16296 (.A1(W20224), .A2(W17606), .ZN(W27283));
  NOR2X1 G16297 (.A1(W1182), .A2(I1854), .ZN(W5617));
  NOR2X1 G16298 (.A1(W2844), .A2(W17221), .ZN(O15091));
  NOR2X1 G16299 (.A1(W2240), .A2(W4730), .ZN(O2711));
  NOR2X1 G16300 (.A1(I858), .A2(W3803), .ZN(W5068));
  NOR2X1 G16301 (.A1(W36788), .A2(W14193), .ZN(W44540));
  NOR2X1 G16302 (.A1(W25675), .A2(W12843), .ZN(O4051));
  NOR2X1 G16303 (.A1(W14886), .A2(W6159), .ZN(W27524));
  NOR2X1 G16304 (.A1(W16156), .A2(W3702), .ZN(W23492));
  NOR2X1 G16305 (.A1(W16229), .A2(W15902), .ZN(W23491));
  NOR2X1 G16306 (.A1(W19724), .A2(W17325), .ZN(O2758));
  NOR2X1 G16307 (.A1(W442), .A2(W23714), .ZN(O15089));
  NOR2X1 G16308 (.A1(W1381), .A2(W22490), .ZN(O14673));
  NOR2X1 G16309 (.A1(W3285), .A2(W980), .ZN(W5074));
  NOR2X1 G16310 (.A1(W7646), .A2(W22666), .ZN(W23217));
  NOR2X1 G16311 (.A1(W17839), .A2(W6577), .ZN(W45890));
  NOR2X1 G16312 (.A1(W2359), .A2(I895), .ZN(W6357));
  NOR2X1 G16313 (.A1(I1730), .A2(W893), .ZN(W5823));
  NOR2X1 G16314 (.A1(W20772), .A2(W7610), .ZN(O2782));
  NOR2X1 G16315 (.A1(W16768), .A2(W6690), .ZN(W45086));
  NOR2X1 G16316 (.A1(W836), .A2(W2189), .ZN(W5530));
  NOR2X1 G16317 (.A1(I1825), .A2(W520), .ZN(W6375));
  NOR2X1 G16318 (.A1(W4295), .A2(W4211), .ZN(W5393));
  NOR2X1 G16319 (.A1(W16238), .A2(W36690), .ZN(O14001));
  NOR2X1 G16320 (.A1(W2231), .A2(W2217), .ZN(W6360));
  NOR2X1 G16321 (.A1(W4142), .A2(W2918), .ZN(W6361));
  NOR2X1 G16322 (.A1(W8828), .A2(W7409), .ZN(W27285));
  NOR2X1 G16323 (.A1(W4615), .A2(W4965), .ZN(W6362));
  NOR2X1 G16324 (.A1(W1348), .A2(W4242), .ZN(W6363));
  NOR2X1 G16325 (.A1(W2885), .A2(I1110), .ZN(W5824));
  NOR2X1 G16326 (.A1(W19660), .A2(W16829), .ZN(W23215));
  NOR2X1 G16327 (.A1(I963), .A2(W4103), .ZN(W6387));
  NOR2X1 G16328 (.A1(W3397), .A2(I1484), .ZN(W5063));
  NOR2X1 G16329 (.A1(I1182), .A2(I1052), .ZN(W5062));
  NOR2X1 G16330 (.A1(W3617), .A2(W3036), .ZN(W5847));
  NOR2X1 G16331 (.A1(W3136), .A2(W1171), .ZN(W5061));
  NOR2X1 G16332 (.A1(W350), .A2(W4314), .ZN(W5060));
  NOR2X1 G16333 (.A1(W4612), .A2(W1051), .ZN(W6385));
  NOR2X1 G16334 (.A1(W12326), .A2(W3177), .ZN(W27281));
  NOR2X1 G16335 (.A1(W1489), .A2(W4380), .ZN(W6386));
  NOR2X1 G16336 (.A1(W15712), .A2(W23752), .ZN(W27185));
  NOR2X1 G16337 (.A1(W2790), .A2(W18905), .ZN(W23463));
  NOR2X1 G16338 (.A1(W14670), .A2(W3155), .ZN(W23490));
  NOR2X1 G16339 (.A1(W18966), .A2(W28757), .ZN(O14802));
  NOR2X1 G16340 (.A1(W951), .A2(W2364), .ZN(W5609));
  NOR2X1 G16341 (.A1(W3430), .A2(W13579), .ZN(W27252));
  NOR2X1 G16342 (.A1(W36592), .A2(W40686), .ZN(O14607));
  NOR2X1 G16343 (.A1(W24546), .A2(W9809), .ZN(W27525));
  NOR2X1 G16344 (.A1(W24587), .A2(W9941), .ZN(W27527));
  NOR2X1 G16345 (.A1(W17335), .A2(W27956), .ZN(O14608));
  NOR2X1 G16346 (.A1(W25689), .A2(W44540), .ZN(O14663));
  NOR2X1 G16347 (.A1(W21269), .A2(W5009), .ZN(O2709));
  NOR2X1 G16348 (.A1(W9403), .A2(W2860), .ZN(O13982));
  NOR2X1 G16349 (.A1(W1033), .A2(W7663), .ZN(W23210));
  NOR2X1 G16350 (.A1(W11588), .A2(W30046), .ZN(O14670));
  NOR2X1 G16351 (.A1(W10893), .A2(W21734), .ZN(O2841));
  NOR2X1 G16352 (.A1(W36873), .A2(W27048), .ZN(O13987));
  NOR2X1 G16353 (.A1(W3814), .A2(W4943), .ZN(W5534));
  NOR2X1 G16354 (.A1(W3135), .A2(W5301), .ZN(W6378));
  NOR2X1 G16355 (.A1(I1812), .A2(W4776), .ZN(W5615));
  NOR2X1 G16356 (.A1(W43173), .A2(W26219), .ZN(O14784));
  NOR2X1 G16357 (.A1(W8370), .A2(I52), .ZN(O13984));
  NOR2X1 G16358 (.A1(W1095), .A2(W1922), .ZN(W6380));
  NOR2X1 G16359 (.A1(W17076), .A2(W38614), .ZN(O15113));
  NOR2X1 G16360 (.A1(W27487), .A2(W8672), .ZN(O13981));
  NOR2X1 G16361 (.A1(W490), .A2(I1225), .ZN(W23544));
  NOR2X1 G16362 (.A1(W4391), .A2(W3792), .ZN(W5414));
  NOR2X1 G16363 (.A1(W30210), .A2(W44023), .ZN(O14603));
  NOR2X1 G16364 (.A1(W2412), .A2(W5227), .ZN(W5613));
  NOR2X1 G16365 (.A1(W6007), .A2(W8726), .ZN(W27359));
  NOR2X1 G16366 (.A1(W20105), .A2(W43654), .ZN(O15096));
  NOR2X1 G16367 (.A1(W935), .A2(W547), .ZN(W6383));
  NOR2X1 G16368 (.A1(W30997), .A2(W23153), .ZN(W44529));
  NOR2X1 G16369 (.A1(I1332), .A2(W4923), .ZN(W6487));
  NOR2X1 G16370 (.A1(W34876), .A2(W8867), .ZN(O13906));
  NOR2X1 G16371 (.A1(W3330), .A2(W250), .ZN(O72));
  NOR2X1 G16372 (.A1(W4731), .A2(W1914), .ZN(W5831));
  NOR2X1 G16373 (.A1(W5753), .A2(W3021), .ZN(W6483));
  NOR2X1 G16374 (.A1(W26964), .A2(I447), .ZN(O4045));
  NOR2X1 G16375 (.A1(W12901), .A2(W5130), .ZN(W27049));
  NOR2X1 G16376 (.A1(W14978), .A2(W18237), .ZN(W27258));
  NOR2X1 G16377 (.A1(W8260), .A2(W25646), .ZN(O4144));
  NOR2X1 G16378 (.A1(W4058), .A2(W24900), .ZN(W27551));
  NOR2X1 G16379 (.A1(W25841), .A2(W3730), .ZN(O13901));
  NOR2X1 G16380 (.A1(W2322), .A2(W20089), .ZN(O13907));
  NOR2X1 G16381 (.A1(W23367), .A2(W12839), .ZN(O13900));
  NOR2X1 G16382 (.A1(W38195), .A2(W10711), .ZN(O15138));
  NOR2X1 G16383 (.A1(W44131), .A2(W14462), .ZN(O13897));
  NOR2X1 G16384 (.A1(W21640), .A2(W44167), .ZN(O14791));
  NOR2X1 G16385 (.A1(W289), .A2(W31014), .ZN(O13895));
  NOR2X1 G16386 (.A1(W4131), .A2(I676), .ZN(W6492));
  NOR2X1 G16387 (.A1(W4308), .A2(I1743), .ZN(W27266));
  NOR2X1 G16388 (.A1(W1623), .A2(W31890), .ZN(O15140));
  NOR2X1 G16389 (.A1(W2839), .A2(W14903), .ZN(W23174));
  NOR2X1 G16390 (.A1(W21589), .A2(W25683), .ZN(O4046));
  NOR2X1 G16391 (.A1(W4742), .A2(W4033), .ZN(W6470));
  NOR2X1 G16392 (.A1(W4554), .A2(I1669), .ZN(W6471));
  NOR2X1 G16393 (.A1(W2218), .A2(W3999), .ZN(W5584));
  NOR2X1 G16394 (.A1(W36319), .A2(W23255), .ZN(W45328));
  NOR2X1 G16395 (.A1(I565), .A2(W797), .ZN(O133));
  NOR2X1 G16396 (.A1(W1691), .A2(I1648), .ZN(W6473));
  NOR2X1 G16397 (.A1(W5487), .A2(W19117), .ZN(O2698));
  NOR2X1 G16398 (.A1(W1297), .A2(W323), .ZN(W5582));
  NOR2X1 G16399 (.A1(W2611), .A2(W4500), .ZN(W5016));
  NOR2X1 G16400 (.A1(W5768), .A2(W839), .ZN(W6475));
  NOR2X1 G16401 (.A1(W26411), .A2(W27171), .ZN(O14631));
  NOR2X1 G16402 (.A1(W2930), .A2(W874), .ZN(W6477));
  NOR2X1 G16403 (.A1(W14155), .A2(W12853), .ZN(W27189));
  NOR2X1 G16404 (.A1(W36914), .A2(I580), .ZN(O13911));
  NOR2X1 G16405 (.A1(W26396), .A2(W13769), .ZN(O13910));
  NOR2X1 G16406 (.A1(W4046), .A2(W2528), .ZN(W5580));
  NOR2X1 G16407 (.A1(W4047), .A2(W12924), .ZN(O14647));
  NOR2X1 G16408 (.A1(W7587), .A2(W14498), .ZN(O13909));
  NOR2X1 G16409 (.A1(W22243), .A2(W14316), .ZN(W45948));
  NOR2X1 G16410 (.A1(W38882), .A2(W21608), .ZN(O14443));
  NOR2X1 G16411 (.A1(W6139), .A2(W18843), .ZN(O2761));
  NOR2X1 G16412 (.A1(W29440), .A2(W5052), .ZN(W44406));
  NOR2X1 G16413 (.A1(W1460), .A2(W5118), .ZN(O134));
  NOR2X1 G16414 (.A1(W5517), .A2(W3080), .ZN(W5571));
  NOR2X1 G16415 (.A1(W29752), .A2(I806), .ZN(O15141));
  NOR2X1 G16416 (.A1(W25137), .A2(W15407), .ZN(O14637));
  NOR2X1 G16417 (.A1(I1258), .A2(W2242), .ZN(W5827));
  NOR2X1 G16418 (.A1(W3493), .A2(W3866), .ZN(W5007));
  NOR2X1 G16419 (.A1(W4778), .A2(W462), .ZN(W5006));
  NOR2X1 G16420 (.A1(W7835), .A2(W39101), .ZN(O15144));
  NOR2X1 G16421 (.A1(W4601), .A2(W5081), .ZN(W5569));
  NOR2X1 G16422 (.A1(W20050), .A2(W31703), .ZN(O13875));
  NOR2X1 G16423 (.A1(W9273), .A2(W1769), .ZN(O4043));
  NOR2X1 G16424 (.A1(W37583), .A2(W8297), .ZN(O15145));
  NOR2X1 G16425 (.A1(W14970), .A2(W5885), .ZN(O4146));
  NOR2X1 G16426 (.A1(W9279), .A2(W26548), .ZN(W44403));
  NOR2X1 G16427 (.A1(W2979), .A2(W2119), .ZN(O14639));
  NOR2X1 G16428 (.A1(W4867), .A2(I660), .ZN(W6513));
  NOR2X1 G16429 (.A1(W17568), .A2(W8942), .ZN(W27354));
  NOR2X1 G16430 (.A1(W29722), .A2(W6126), .ZN(O13872));
  NOR2X1 G16431 (.A1(W3004), .A2(W5309), .ZN(W5566));
  NOR2X1 G16432 (.A1(I943), .A2(W3517), .ZN(W6502));
  NOR2X1 G16433 (.A1(I175), .A2(W3771), .ZN(W6495));
  NOR2X1 G16434 (.A1(W43538), .A2(W18349), .ZN(O13891));
  NOR2X1 G16435 (.A1(W28330), .A2(I1020), .ZN(O13890));
  NOR2X1 G16436 (.A1(W40714), .A2(W29507), .ZN(W45336));
  NOR2X1 G16437 (.A1(W3851), .A2(W4326), .ZN(O13885));
  NOR2X1 G16438 (.A1(W13941), .A2(W20480), .ZN(O13884));
  NOR2X1 G16439 (.A1(W5078), .A2(I660), .ZN(O14634));
  NOR2X1 G16440 (.A1(W9856), .A2(W18255), .ZN(W44415));
  NOR2X1 G16441 (.A1(W10046), .A2(W2927), .ZN(O4041));
  NOR2X1 G16442 (.A1(W34342), .A2(W37418), .ZN(W44414));
  NOR2X1 G16443 (.A1(W3138), .A2(I350), .ZN(W6469));
  NOR2X1 G16444 (.A1(I1972), .A2(W1541), .ZN(W5409));
  NOR2X1 G16445 (.A1(W4121), .A2(W1032), .ZN(W5574));
  NOR2X1 G16446 (.A1(W481), .A2(W3139), .ZN(W6503));
  NOR2X1 G16447 (.A1(W5809), .A2(W3171), .ZN(W6504));
  NOR2X1 G16448 (.A1(W6308), .A2(W14576), .ZN(O4044));
  NOR2X1 G16449 (.A1(W198), .A2(I1175), .ZN(W5010));
  NOR2X1 G16450 (.A1(W4025), .A2(W6471), .ZN(W6505));
  NOR2X1 G16451 (.A1(W2206), .A2(W4893), .ZN(W6506));
  NOR2X1 G16452 (.A1(W15416), .A2(W13237), .ZN(W27558));
  NOR2X1 G16453 (.A1(W4350), .A2(W3386), .ZN(W5553));
  NOR2X1 G16454 (.A1(W12358), .A2(W6647), .ZN(W44478));
  NOR2X1 G16455 (.A1(W44603), .A2(W23826), .ZN(O14659));
  NOR2X1 G16456 (.A1(W26640), .A2(W12440), .ZN(O13936));
  NOR2X1 G16457 (.A1(W4332), .A2(W19830), .ZN(W23193));
  NOR2X1 G16458 (.A1(W22328), .A2(I330), .ZN(W45322));
  NOR2X1 G16459 (.A1(W11575), .A2(I1005), .ZN(O13934));
  NOR2X1 G16460 (.A1(W5824), .A2(W2955), .ZN(W5839));
  NOR2X1 G16461 (.A1(I1179), .A2(W1747), .ZN(W5590));
  NOR2X1 G16462 (.A1(W38556), .A2(W33211), .ZN(W44473));
  NOR2X1 G16463 (.A1(W13114), .A2(W26613), .ZN(O3971));
  NOR2X1 G16464 (.A1(W1029), .A2(W1206), .ZN(W5550));
  NOR2X1 G16465 (.A1(I1784), .A2(W13095), .ZN(W27538));
  NOR2X1 G16466 (.A1(I355), .A2(W5778), .ZN(W6447));
  NOR2X1 G16467 (.A1(W14135), .A2(W26045), .ZN(O13932));
  NOR2X1 G16468 (.A1(W13830), .A2(W24983), .ZN(W27539));
  NOR2X1 G16469 (.A1(W1504), .A2(W4525), .ZN(W6450));
  NOR2X1 G16470 (.A1(W1671), .A2(W3761), .ZN(W5031));
  NOR2X1 G16471 (.A1(W18221), .A2(W21748), .ZN(W27256));
  NOR2X1 G16472 (.A1(W19834), .A2(W21320), .ZN(O2792));
  NOR2X1 G16473 (.A1(W7982), .A2(W8950), .ZN(W23189));
  NOR2X1 G16474 (.A1(W1491), .A2(W2937), .ZN(W6434));
  NOR2X1 G16475 (.A1(W27314), .A2(W16568), .ZN(O14619));
  NOR2X1 G16476 (.A1(W9907), .A2(W8647), .ZN(W23196));
  NOR2X1 G16477 (.A1(W3958), .A2(W5435), .ZN(W5596));
  NOR2X1 G16478 (.A1(W2045), .A2(W4098), .ZN(W5401));
  NOR2X1 G16479 (.A1(W33146), .A2(W23520), .ZN(O14620));
  NOR2X1 G16480 (.A1(W15885), .A2(W33095), .ZN(W45919));
  NOR2X1 G16481 (.A1(W19458), .A2(W13824), .ZN(W44487));
  NOR2X1 G16482 (.A1(I794), .A2(W1941), .ZN(W6432));
  NOR2X1 G16483 (.A1(W2743), .A2(W12220), .ZN(O2703));
  NOR2X1 G16484 (.A1(W6062), .A2(W667), .ZN(W23541));
  NOR2X1 G16485 (.A1(W2886), .A2(W6307), .ZN(W44467));
  NOR2X1 G16486 (.A1(I901), .A2(I995), .ZN(W6435));
  NOR2X1 G16487 (.A1(I286), .A2(I5), .ZN(W6436));
  NOR2X1 G16488 (.A1(W1227), .A2(W41833), .ZN(W45367));
  NOR2X1 G16489 (.A1(W5175), .A2(W11467), .ZN(O13942));
  NOR2X1 G16490 (.A1(W3089), .A2(W1484), .ZN(W6438));
  NOR2X1 G16491 (.A1(W290), .A2(W2974), .ZN(W5549));
  NOR2X1 G16492 (.A1(W28820), .A2(W28263), .ZN(O13938));
  NOR2X1 G16493 (.A1(W5146), .A2(W657), .ZN(W5593));
  NOR2X1 G16494 (.A1(I1519), .A2(I1314), .ZN(W5592));
  NOR2X1 G16495 (.A1(W13570), .A2(W15859), .ZN(W23183));
  NOR2X1 G16496 (.A1(W2702), .A2(W43801), .ZN(O14789));
  NOR2X1 G16497 (.A1(W3591), .A2(W1101), .ZN(W6464));
  NOR2X1 G16498 (.A1(W35749), .A2(W19515), .ZN(O15124));
  NOR2X1 G16499 (.A1(W5270), .A2(W3318), .ZN(W5558));
  NOR2X1 G16500 (.A1(I1576), .A2(W18297), .ZN(O2790));
  NOR2X1 G16501 (.A1(W4654), .A2(W18931), .ZN(W23479));
  NOR2X1 G16502 (.A1(W3295), .A2(W36717), .ZN(O14447));
  NOR2X1 G16503 (.A1(W19962), .A2(W32094), .ZN(O15126));
  NOR2X1 G16504 (.A1(W1293), .A2(W25753), .ZN(O15127));
  NOR2X1 G16505 (.A1(I228), .A2(W21639), .ZN(O2789));
  NOR2X1 G16506 (.A1(W27641), .A2(W11848), .ZN(O14625));
  NOR2X1 G16507 (.A1(I1253), .A2(W3375), .ZN(W5586));
  NOR2X1 G16508 (.A1(W37301), .A2(W39235), .ZN(W44456));
  NOR2X1 G16509 (.A1(W6007), .A2(W6205), .ZN(O2847));
  NOR2X1 G16510 (.A1(W14340), .A2(W23464), .ZN(W27051));
  NOR2X1 G16511 (.A1(I1222), .A2(W1865), .ZN(W5834));
  NOR2X1 G16512 (.A1(W14567), .A2(W33224), .ZN(O14793));
  NOR2X1 G16513 (.A1(W2015), .A2(W3313), .ZN(W5585));
  NOR2X1 G16514 (.A1(W8228), .A2(W9256), .ZN(W23181));
  NOR2X1 G16515 (.A1(W4700), .A2(W4295), .ZN(W5833));
  NOR2X1 G16516 (.A1(W5019), .A2(W4083), .ZN(W5836));
  NOR2X1 G16517 (.A1(I1149), .A2(W2289), .ZN(W5030));
  NOR2X1 G16518 (.A1(W25194), .A2(W25984), .ZN(W45929));
  NOR2X1 G16519 (.A1(W24387), .A2(W20613), .ZN(W27541));
  NOR2X1 G16520 (.A1(W3709), .A2(I780), .ZN(W5403));
  NOR2X1 G16521 (.A1(I1909), .A2(W540), .ZN(W6455));
  NOR2X1 G16522 (.A1(W2362), .A2(I726), .ZN(W6456));
  NOR2X1 G16523 (.A1(W19071), .A2(W10028), .ZN(O14437));
  NOR2X1 G16524 (.A1(W17716), .A2(W17395), .ZN(W27542));
  NOR2X1 G16525 (.A1(I1146), .A2(W17933), .ZN(O13926));
  NOR2X1 G16526 (.A1(W3391), .A2(W13487), .ZN(W23399));
  NOR2X1 G16527 (.A1(W10731), .A2(W13525), .ZN(O13923));
  NOR2X1 G16528 (.A1(W12745), .A2(W37586), .ZN(O15118));
  NOR2X1 G16529 (.A1(W17963), .A2(W3800), .ZN(O15119));
  NOR2X1 G16530 (.A1(W22974), .A2(W14531), .ZN(O14622));
  NOR2X1 G16531 (.A1(W32093), .A2(W4908), .ZN(O14651));
  NOR2X1 G16532 (.A1(W2832), .A2(W3392), .ZN(W27056));
  NOR2X1 G16533 (.A1(W11924), .A2(W2182), .ZN(O4143));
  NOR2X1 G16534 (.A1(W5361), .A2(I1281), .ZN(W6463));
  NOR2X1 G16535 (.A1(W1093), .A2(W2644), .ZN(W5405));
  NOR2X1 G16536 (.A1(W6305), .A2(I404), .ZN(W27297));
  NOR2X1 G16537 (.A1(W29947), .A2(W14514), .ZN(W44656));
  NOR2X1 G16538 (.A1(W16), .A2(W3078), .ZN(W5386));
  NOR2X1 G16539 (.A1(W11162), .A2(W26749), .ZN(O14690));
  NOR2X1 G16540 (.A1(W29587), .A2(W5953), .ZN(O14086));
  NOR2X1 G16541 (.A1(I1385), .A2(W7406), .ZN(W23637));
  NOR2X1 G16542 (.A1(W4884), .A2(W2103), .ZN(W5664));
  NOR2X1 G16543 (.A1(W36675), .A2(W37779), .ZN(O14084));
  NOR2X1 G16544 (.A1(W738), .A2(I1768), .ZN(W6262));
  NOR2X1 G16545 (.A1(I713), .A2(W5738), .ZN(W6263));
  NOR2X1 G16546 (.A1(W11697), .A2(W16773), .ZN(O14450));
  NOR2X1 G16547 (.A1(W43402), .A2(W8619), .ZN(W44660));
  NOR2X1 G16548 (.A1(W11225), .A2(W11999), .ZN(W23247));
  NOR2X1 G16549 (.A1(W7568), .A2(W21454), .ZN(W27496));
  NOR2X1 G16550 (.A1(W19407), .A2(W26490), .ZN(O4124));
  NOR2X1 G16551 (.A1(W32179), .A2(W26402), .ZN(W45232));
  NOR2X1 G16552 (.A1(W38136), .A2(W8127), .ZN(O14569));
  NOR2X1 G16553 (.A1(I494), .A2(W3537), .ZN(W6267));
  NOR2X1 G16554 (.A1(W2290), .A2(W8673), .ZN(O4125));
  NOR2X1 G16555 (.A1(W15059), .A2(W22571), .ZN(W27296));
  NOR2X1 G16556 (.A1(W6928), .A2(W6624), .ZN(O14078));
  NOR2X1 G16557 (.A1(W36487), .A2(W39530), .ZN(W44667));
  NOR2X1 G16558 (.A1(W23862), .A2(W6165), .ZN(O14691));
  NOR2X1 G16559 (.A1(I747), .A2(W4427), .ZN(W6218));
  NOR2X1 G16560 (.A1(W13112), .A2(W1148), .ZN(O14565));
  NOR2X1 G16561 (.A1(W25818), .A2(W26993), .ZN(O14096));
  NOR2X1 G16562 (.A1(W17813), .A2(W14111), .ZN(O2723));
  NOR2X1 G16563 (.A1(W14508), .A2(W41670), .ZN(W45249));
  NOR2X1 G16564 (.A1(W12662), .A2(W530), .ZN(W27096));
  NOR2X1 G16565 (.A1(W30534), .A2(W2577), .ZN(O14566));
  NOR2X1 G16566 (.A1(W22707), .A2(W9408), .ZN(O14093));
  NOR2X1 G16567 (.A1(W4386), .A2(W2222), .ZN(W5868));
  NOR2X1 G16568 (.A1(W43926), .A2(W27183), .ZN(O14567));
  NOR2X1 G16569 (.A1(W10108), .A2(W24320), .ZN(O14568));
  NOR2X1 G16570 (.A1(I681), .A2(I1599), .ZN(W5666));
  NOR2X1 G16571 (.A1(W6129), .A2(W1225), .ZN(O4121));
  NOR2X1 G16572 (.A1(W8876), .A2(W34690), .ZN(O14452));
  NOR2X1 G16573 (.A1(W1581), .A2(I1277), .ZN(W5816));
  NOR2X1 G16574 (.A1(I448), .A2(W2570), .ZN(W5134));
  NOR2X1 G16575 (.A1(W21296), .A2(W13087), .ZN(W23380));
  NOR2X1 G16576 (.A1(W1002), .A2(W3090), .ZN(W5665));
  NOR2X1 G16577 (.A1(W31600), .A2(W38174), .ZN(O15047));
  NOR2X1 G16578 (.A1(W12780), .A2(W14305), .ZN(W23241));
  NOR2X1 G16579 (.A1(W16929), .A2(W37738), .ZN(O14068));
  NOR2X1 G16580 (.A1(W41828), .A2(W4574), .ZN(O14067));
  NOR2X1 G16581 (.A1(W29194), .A2(W26746), .ZN(O14065));
  NOR2X1 G16582 (.A1(W23941), .A2(W37735), .ZN(O14064));
  NOR2X1 G16583 (.A1(W27661), .A2(W31062), .ZN(O14063));
  NOR2X1 G16584 (.A1(W3418), .A2(I778), .ZN(W6280));
  NOR2X1 G16585 (.A1(W77), .A2(W44375), .ZN(O14061));
  NOR2X1 G16586 (.A1(I1531), .A2(W3948), .ZN(W5867));
  NOR2X1 G16587 (.A1(W616), .A2(W2972), .ZN(W6282));
  NOR2X1 G16588 (.A1(W8468), .A2(W5774), .ZN(O15046));
  NOR2X1 G16589 (.A1(W25591), .A2(W13152), .ZN(O3980));
  NOR2X1 G16590 (.A1(W20002), .A2(W4783), .ZN(W23240));
  NOR2X1 G16591 (.A1(W2737), .A2(I1196), .ZN(O14687));
  NOR2X1 G16592 (.A1(W11406), .A2(W27758), .ZN(O14059));
  NOR2X1 G16593 (.A1(W13673), .A2(W11285), .ZN(O14122));
  NOR2X1 G16594 (.A1(W3127), .A2(W2764), .ZN(W5866));
  NOR2X1 G16595 (.A1(W35765), .A2(W24958), .ZN(W45837));
  NOR2X1 G16596 (.A1(W42351), .A2(W34895), .ZN(O15050));
  NOR2X1 G16597 (.A1(W15742), .A2(I740), .ZN(O14058));
  NOR2X1 G16598 (.A1(W12593), .A2(W31382), .ZN(O14572));
  NOR2X1 G16599 (.A1(W15991), .A2(W16121), .ZN(O2720));
  NOR2X1 G16600 (.A1(W5041), .A2(W1770), .ZN(W5660));
  NOR2X1 G16601 (.A1(W31599), .A2(W18927), .ZN(O14076));
  NOR2X1 G16602 (.A1(W3411), .A2(W67), .ZN(W5131));
  NOR2X1 G16603 (.A1(W35822), .A2(W21521), .ZN(O15041));
  NOR2X1 G16604 (.A1(W31587), .A2(W9841), .ZN(O14571));
  NOR2X1 G16605 (.A1(W8876), .A2(W21578), .ZN(W27242));
  NOR2X1 G16606 (.A1(W3801), .A2(W9513), .ZN(W23639));
  NOR2X1 G16607 (.A1(W30396), .A2(W34941), .ZN(W45832));
  NOR2X1 G16608 (.A1(W4897), .A2(W5911), .ZN(W6219));
  NOR2X1 G16609 (.A1(W1674), .A2(W3025), .ZN(W5872));
  NOR2X1 G16610 (.A1(I247), .A2(I1404), .ZN(W5657));
  NOR2X1 G16611 (.A1(I230), .A2(W4457), .ZN(W5127));
  NOR2X1 G16612 (.A1(W6995), .A2(W19321), .ZN(W23242));
  NOR2X1 G16613 (.A1(W17691), .A2(W5716), .ZN(O14776));
  NOR2X1 G16614 (.A1(W12925), .A2(W20033), .ZN(O2778));
  NOR2X1 G16615 (.A1(W2300), .A2(W39914), .ZN(O14074));
  NOR2X1 G16616 (.A1(W6911), .A2(W11583), .ZN(O14688));
  NOR2X1 G16617 (.A1(I1770), .A2(W441), .ZN(W5126));
  NOR2X1 G16618 (.A1(W6721), .A2(W15079), .ZN(W23627));
  NOR2X1 G16619 (.A1(W37341), .A2(W24006), .ZN(O14113));
  NOR2X1 G16620 (.A1(W42470), .A2(W2489), .ZN(O14780));
  NOR2X1 G16621 (.A1(W21118), .A2(W16098), .ZN(O15027));
  NOR2X1 G16622 (.A1(I1803), .A2(I936), .ZN(W6230));
  NOR2X1 G16623 (.A1(W22399), .A2(W4168), .ZN(O4033));
  NOR2X1 G16624 (.A1(W20990), .A2(W39507), .ZN(O15020));
  NOR2X1 G16625 (.A1(W16889), .A2(W14310), .ZN(O4058));
  NOR2X1 G16626 (.A1(W3221), .A2(W5363), .ZN(W6231));
  NOR2X1 G16627 (.A1(W29003), .A2(W45075), .ZN(O14695));
  NOR2X1 G16628 (.A1(I1664), .A2(W2236), .ZN(W5680));
  NOR2X1 G16629 (.A1(W1895), .A2(W4506), .ZN(W27476));
  NOR2X1 G16630 (.A1(W14469), .A2(W25536), .ZN(O14112));
  NOR2X1 G16631 (.A1(W6474), .A2(W33869), .ZN(O14693));
  NOR2X1 G16632 (.A1(W4723), .A2(W2920), .ZN(O75));
  NOR2X1 G16633 (.A1(W35107), .A2(W24164), .ZN(W45813));
  NOR2X1 G16634 (.A1(W3921), .A2(W4500), .ZN(O97));
  NOR2X1 G16635 (.A1(W2342), .A2(W3922), .ZN(W5150));
  NOR2X1 G16636 (.A1(W4443), .A2(W3643), .ZN(W5149));
  NOR2X1 G16637 (.A1(W31051), .A2(W4878), .ZN(W45234));
  NOR2X1 G16638 (.A1(W5277), .A2(W2201), .ZN(W23261));
  NOR2X1 G16639 (.A1(W1922), .A2(I1373), .ZN(W6224));
  NOR2X1 G16640 (.A1(W26305), .A2(W22135), .ZN(O14407));
  NOR2X1 G16641 (.A1(W4011), .A2(W4333), .ZN(W5161));
  NOR2X1 G16642 (.A1(W1161), .A2(W1748), .ZN(W5382));
  NOR2X1 G16643 (.A1(W4419), .A2(W23130), .ZN(O15021));
  NOR2X1 G16644 (.A1(W5531), .A2(W4634), .ZN(W27302));
  NOR2X1 G16645 (.A1(W2055), .A2(W2626), .ZN(W5159));
  NOR2X1 G16646 (.A1(W39849), .A2(W28440), .ZN(W44702));
  NOR2X1 G16647 (.A1(W14039), .A2(W21594), .ZN(W45236));
  NOR2X1 G16648 (.A1(W8044), .A2(W9709), .ZN(O2833));
  NOR2X1 G16649 (.A1(W26255), .A2(W21223), .ZN(O14110));
  NOR2X1 G16650 (.A1(W16522), .A2(W1509), .ZN(O15026));
  NOR2X1 G16651 (.A1(W31116), .A2(W21802), .ZN(O14116));
  NOR2X1 G16652 (.A1(W3371), .A2(W80), .ZN(W5156));
  NOR2X1 G16653 (.A1(W26470), .A2(W30356), .ZN(O14556));
  NOR2X1 G16654 (.A1(W40552), .A2(W18630), .ZN(O14697));
  NOR2X1 G16655 (.A1(I802), .A2(W20022), .ZN(W27474));
  NOR2X1 G16656 (.A1(W16716), .A2(W13396), .ZN(W45411));
  NOR2X1 G16657 (.A1(W26663), .A2(W18763), .ZN(W27475));
  NOR2X1 G16658 (.A1(W1711), .A2(I1069), .ZN(W5155));
  NOR2X1 G16659 (.A1(W24196), .A2(W7169), .ZN(W27101));
  NOR2X1 G16660 (.A1(I1912), .A2(W2280), .ZN(W5676));
  NOR2X1 G16661 (.A1(W4202), .A2(W3617), .ZN(W5144));
  NOR2X1 G16662 (.A1(W21719), .A2(W18541), .ZN(O14106));
  NOR2X1 G16663 (.A1(W818), .A2(W2105), .ZN(W27299));
  NOR2X1 G16664 (.A1(W29487), .A2(I1674), .ZN(W45245));
  NOR2X1 G16665 (.A1(W9653), .A2(W3049), .ZN(W23258));
  NOR2X1 G16666 (.A1(W440), .A2(W2232), .ZN(W27481));
  NOR2X1 G16667 (.A1(I435), .A2(W3956), .ZN(W5142));
  NOR2X1 G16668 (.A1(W2164), .A2(I1531), .ZN(W6245));
  NOR2X1 G16669 (.A1(W4394), .A2(I925), .ZN(W5509));
  NOR2X1 G16670 (.A1(W26042), .A2(W18305), .ZN(W27471));
  NOR2X1 G16671 (.A1(I1121), .A2(W163), .ZN(W5140));
  NOR2X1 G16672 (.A1(W23609), .A2(W20627), .ZN(O2834));
  NOR2X1 G16673 (.A1(W1231), .A2(W1085), .ZN(W5385));
  NOR2X1 G16674 (.A1(W19028), .A2(I721), .ZN(W23256));
  NOR2X1 G16675 (.A1(W4539), .A2(I181), .ZN(W5672));
  NOR2X1 G16676 (.A1(I244), .A2(I1214), .ZN(W23633));
  NOR2X1 G16677 (.A1(W12463), .A2(W21952), .ZN(W27483));
  NOR2X1 G16678 (.A1(W22391), .A2(W5201), .ZN(W23634));
  NOR2X1 G16679 (.A1(W27847), .A2(W38906), .ZN(O14692));
  NOR2X1 G16680 (.A1(W21802), .A2(W12974), .ZN(W23628));
  NOR2X1 G16681 (.A1(I490), .A2(W13696), .ZN(W23629));
  NOR2X1 G16682 (.A1(W13481), .A2(W2672), .ZN(O14118));
  NOR2X1 G16683 (.A1(I896), .A2(W5720), .ZN(W6235));
  NOR2X1 G16684 (.A1(W3345), .A2(W4321), .ZN(W5146));
  NOR2X1 G16685 (.A1(W28257), .A2(W25400), .ZN(O14560));
  NOR2X1 G16686 (.A1(W33907), .A2(W27338), .ZN(O14109));
  NOR2X1 G16687 (.A1(W21486), .A2(W22945), .ZN(O14561));
  NOR2X1 G16688 (.A1(W9490), .A2(W22562), .ZN(W27478));
  NOR2X1 G16689 (.A1(W12508), .A2(W19733), .ZN(W23381));
  NOR2X1 G16690 (.A1(W1488), .A2(W2362), .ZN(W5145));
  NOR2X1 G16691 (.A1(W37350), .A2(W42430), .ZN(W44687));
  NOR2X1 G16692 (.A1(W40281), .A2(W41823), .ZN(W44686));
  NOR2X1 G16693 (.A1(W9970), .A2(W32106), .ZN(O14811));
  NOR2X1 G16694 (.A1(I203), .A2(W771), .ZN(W5384));
  NOR2X1 G16695 (.A1(W10128), .A2(W1023), .ZN(W27480));
  NOR2X1 G16696 (.A1(W23571), .A2(W11077), .ZN(O15016));
  NOR2X1 G16697 (.A1(W1171), .A2(W2759), .ZN(W6241));
  NOR2X1 G16698 (.A1(W5420), .A2(W12201), .ZN(O4019));
  NOR2X1 G16699 (.A1(W1803), .A2(W1624), .ZN(W5392));
  NOR2X1 G16700 (.A1(I784), .A2(W3329), .ZN(W6329));
  NOR2X1 G16701 (.A1(W15607), .A2(W43808), .ZN(O14025));
  NOR2X1 G16702 (.A1(W2351), .A2(I1008), .ZN(O14024));
  NOR2X1 G16703 (.A1(W6509), .A2(W16197), .ZN(O2780));
  NOR2X1 G16704 (.A1(W19966), .A2(W44561), .ZN(O14023));
  NOR2X1 G16705 (.A1(W4811), .A2(W1029), .ZN(W27084));
  NOR2X1 G16706 (.A1(W4471), .A2(I1749), .ZN(W5091));
  NOR2X1 G16707 (.A1(W756), .A2(W1257), .ZN(W5090));
  NOR2X1 G16708 (.A1(W1987), .A2(W3245), .ZN(W5522));
  NOR2X1 G16709 (.A1(W2825), .A2(W5262), .ZN(W23225));
  NOR2X1 G16710 (.A1(W8615), .A2(W3610), .ZN(W23226));
  NOR2X1 G16711 (.A1(W21171), .A2(W8616), .ZN(W23650));
  NOR2X1 G16712 (.A1(W2514), .A2(W2725), .ZN(O76));
  NOR2X1 G16713 (.A1(W44487), .A2(W16160), .ZN(O14020));
  NOR2X1 G16714 (.A1(W14435), .A2(I840), .ZN(O2796));
  NOR2X1 G16715 (.A1(W43437), .A2(W19192), .ZN(W45083));
  NOR2X1 G16716 (.A1(W1857), .A2(W6017), .ZN(W6337));
  NOR2X1 G16717 (.A1(W2959), .A2(W42439), .ZN(O14017));
  NOR2X1 G16718 (.A1(W26183), .A2(W26147), .ZN(O14016));
  NOR2X1 G16719 (.A1(W32616), .A2(W36577), .ZN(O15015));
  NOR2X1 G16720 (.A1(W4858), .A2(W812), .ZN(W5689));
  NOR2X1 G16721 (.A1(I457), .A2(W26461), .ZN(W27516));
  NOR2X1 G16722 (.A1(W3636), .A2(W2544), .ZN(W5096));
  NOR2X1 G16723 (.A1(W4911), .A2(W1509), .ZN(W5639));
  NOR2X1 G16724 (.A1(W3026), .A2(W2978), .ZN(W5095));
  NOR2X1 G16725 (.A1(W14065), .A2(W12178), .ZN(O4053));
  NOR2X1 G16726 (.A1(W24144), .A2(W4834), .ZN(W44588));
  NOR2X1 G16727 (.A1(W36995), .A2(W29730), .ZN(W45544));
  NOR2X1 G16728 (.A1(W18306), .A2(W772), .ZN(O14426));
  NOR2X1 G16729 (.A1(W5192), .A2(W2942), .ZN(W6324));
  NOR2X1 G16730 (.A1(W17316), .A2(W3674), .ZN(W27353));
  NOR2X1 G16731 (.A1(W977), .A2(W1401), .ZN(W5854));
  NOR2X1 G16732 (.A1(W4196), .A2(I1843), .ZN(W5637));
  NOR2X1 G16733 (.A1(W2789), .A2(W4820), .ZN(W6325));
  NOR2X1 G16734 (.A1(W300), .A2(W941), .ZN(W5636));
  NOR2X1 G16735 (.A1(W9652), .A2(W12534), .ZN(W27288));
  NOR2X1 G16736 (.A1(W155), .A2(W24920), .ZN(W44587));
  NOR2X1 G16737 (.A1(W40226), .A2(W588), .ZN(O14587));
  NOR2X1 G16738 (.A1(W15184), .A2(W160), .ZN(W27085));
  NOR2X1 G16739 (.A1(I1042), .A2(W5129), .ZN(W6327));
  NOR2X1 G16740 (.A1(W5251), .A2(W22715), .ZN(W27364));
  NOR2X1 G16741 (.A1(W56), .A2(W1821), .ZN(O90));
  NOR2X1 G16742 (.A1(W834), .A2(I1407), .ZN(W5081));
  NOR2X1 G16743 (.A1(W38926), .A2(W36047), .ZN(O14009));
  NOR2X1 G16744 (.A1(W14372), .A2(W17818), .ZN(O2712));
  NOR2X1 G16745 (.A1(W585), .A2(I1982), .ZN(W6350));
  NOR2X1 G16746 (.A1(W18832), .A2(W5762), .ZN(W45879));
  NOR2X1 G16747 (.A1(W36469), .A2(W35069), .ZN(O15082));
  NOR2X1 G16748 (.A1(W19662), .A2(I558), .ZN(W23219));
  NOR2X1 G16749 (.A1(I1778), .A2(W1721), .ZN(O4034));
  NOR2X1 G16750 (.A1(W38471), .A2(W42841), .ZN(O15083));
  NOR2X1 G16751 (.A1(W1926), .A2(W3516), .ZN(W5626));
  NOR2X1 G16752 (.A1(W1521), .A2(W33967), .ZN(O14592));
  NOR2X1 G16753 (.A1(I235), .A2(I1168), .ZN(W5077));
  NOR2X1 G16754 (.A1(W23852), .A2(W20258), .ZN(W45288));
  NOR2X1 G16755 (.A1(W41992), .A2(W17115), .ZN(W44560));
  NOR2X1 G16756 (.A1(W25550), .A2(W13962), .ZN(O14429));
  NOR2X1 G16757 (.A1(W20222), .A2(W23898), .ZN(W27521));
  NOR2X1 G16758 (.A1(W44486), .A2(W43684), .ZN(O14594));
  NOR2X1 G16759 (.A1(I1089), .A2(W4253), .ZN(W6354));
  NOR2X1 G16760 (.A1(W1523), .A2(W5712), .ZN(W6355));
  NOR2X1 G16761 (.A1(W20936), .A2(W1071), .ZN(O15086));
  NOR2X1 G16762 (.A1(W37762), .A2(W15146), .ZN(W44570));
  NOR2X1 G16763 (.A1(W40684), .A2(W14667), .ZN(O14015));
  NOR2X1 G16764 (.A1(W4972), .A2(W23692), .ZN(O14589));
  NOR2X1 G16765 (.A1(W2869), .A2(I868), .ZN(W5087));
  NOR2X1 G16766 (.A1(W9478), .A2(W36897), .ZN(O15077));
  NOR2X1 G16767 (.A1(W11361), .A2(W995), .ZN(O14014));
  NOR2X1 G16768 (.A1(W4850), .A2(W5218), .ZN(W6342));
  NOR2X1 G16769 (.A1(W15717), .A2(W36941), .ZN(O14591));
  NOR2X1 G16770 (.A1(W37215), .A2(W2848), .ZN(O14013));
  NOR2X1 G16771 (.A1(W30806), .A2(W28), .ZN(O14675));
  NOR2X1 G16772 (.A1(I1341), .A2(W2654), .ZN(W5097));
  NOR2X1 G16773 (.A1(I697), .A2(W2026), .ZN(W5085));
  NOR2X1 G16774 (.A1(W2737), .A2(I289), .ZN(W6345));
  NOR2X1 G16775 (.A1(W3885), .A2(W9484), .ZN(O15079));
  NOR2X1 G16776 (.A1(W3376), .A2(I215), .ZN(W5525));
  NOR2X1 G16777 (.A1(W24243), .A2(W12043), .ZN(W45286));
  NOR2X1 G16778 (.A1(W12716), .A2(W17660), .ZN(O15080));
  NOR2X1 G16779 (.A1(W2780), .A2(W94), .ZN(W5628));
  NOR2X1 G16780 (.A1(W15046), .A2(W10546), .ZN(O15081));
  NOR2X1 G16781 (.A1(W201), .A2(I1826), .ZN(O2713));
  NOR2X1 G16782 (.A1(W36999), .A2(W44570), .ZN(O14044));
  NOR2X1 G16783 (.A1(I507), .A2(W4478), .ZN(W5113));
  NOR2X1 G16784 (.A1(W15685), .A2(W6613), .ZN(W23237));
  NOR2X1 G16785 (.A1(W4396), .A2(W422), .ZN(W5112));
  NOR2X1 G16786 (.A1(I1377), .A2(W1227), .ZN(W6299));
  NOR2X1 G16787 (.A1(W28774), .A2(W11504), .ZN(O14577));
  NOR2X1 G16788 (.A1(W11760), .A2(W8315), .ZN(O4079));
  NOR2X1 G16789 (.A1(W18713), .A2(I454), .ZN(W23499));
  NOR2X1 G16790 (.A1(W2031), .A2(W4683), .ZN(W5651));
  NOR2X1 G16791 (.A1(W15689), .A2(W16944), .ZN(O14046));
  NOR2X1 G16792 (.A1(W24697), .A2(W14874), .ZN(O4128));
  NOR2X1 G16793 (.A1(W486), .A2(W26924), .ZN(O14417));
  NOR2X1 G16794 (.A1(W1455), .A2(W4740), .ZN(W6303));
  NOR2X1 G16795 (.A1(W19676), .A2(W33014), .ZN(O14043));
  NOR2X1 G16796 (.A1(W2315), .A2(W1400), .ZN(W5111));
  NOR2X1 G16797 (.A1(W16467), .A2(W15506), .ZN(O14578));
  NOR2X1 G16798 (.A1(W19928), .A2(W2731), .ZN(O15059));
  NOR2X1 G16799 (.A1(W18234), .A2(W37112), .ZN(O14579));
  NOR2X1 G16800 (.A1(W2230), .A2(I339), .ZN(W5108));
  NOR2X1 G16801 (.A1(I344), .A2(W10728), .ZN(O14419));
  NOR2X1 G16802 (.A1(W2692), .A2(W3880), .ZN(W6286));
  NOR2X1 G16803 (.A1(W41492), .A2(W33295), .ZN(O14054));
  NOR2X1 G16804 (.A1(W15124), .A2(I283), .ZN(O14056));
  NOR2X1 G16805 (.A1(W8912), .A2(W9400), .ZN(O4018));
  NOR2X1 G16806 (.A1(W4041), .A2(W12926), .ZN(O2837));
  NOR2X1 G16807 (.A1(W19657), .A2(W13562), .ZN(O14807));
  NOR2X1 G16808 (.A1(W31496), .A2(W37219), .ZN(O15057));
  NOR2X1 G16809 (.A1(W4819), .A2(W2767), .ZN(W5864));
  NOR2X1 G16810 (.A1(W42080), .A2(W250), .ZN(W45265));
  NOR2X1 G16811 (.A1(W18094), .A2(W7201), .ZN(O14055));
  NOR2X1 G16812 (.A1(W2875), .A2(W4247), .ZN(W5116));
  NOR2X1 G16813 (.A1(W42573), .A2(W15543), .ZN(O14042));
  NOR2X1 G16814 (.A1(W24570), .A2(W16072), .ZN(O14053));
  NOR2X1 G16815 (.A1(W3726), .A2(W3612), .ZN(W5115));
  NOR2X1 G16816 (.A1(W5189), .A2(W4840), .ZN(W6292));
  NOR2X1 G16817 (.A1(W43305), .A2(W34993), .ZN(O15058));
  NOR2X1 G16818 (.A1(W56), .A2(W1908), .ZN(W6293));
  NOR2X1 G16819 (.A1(W36079), .A2(W25452), .ZN(O14052));
  NOR2X1 G16820 (.A1(W16032), .A2(W4676), .ZN(O4127));
  NOR2X1 G16821 (.A1(W34349), .A2(W42640), .ZN(O14050));
  NOR2X1 G16822 (.A1(W4571), .A2(I362), .ZN(W6297));
  NOR2X1 G16823 (.A1(W16319), .A2(W9302), .ZN(W27184));
  NOR2X1 G16824 (.A1(W142), .A2(W3182), .ZN(W27088));
  NOR2X1 G16825 (.A1(W14905), .A2(W34667), .ZN(O15063));
  NOR2X1 G16826 (.A1(W1092), .A2(I1994), .ZN(W5642));
  NOR2X1 G16827 (.A1(W18318), .A2(W10479), .ZN(O2757));
  NOR2X1 G16828 (.A1(W26870), .A2(W8389), .ZN(O14677));
  NOR2X1 G16829 (.A1(I1674), .A2(W4382), .ZN(W5102));
  NOR2X1 G16830 (.A1(W1918), .A2(W674), .ZN(W5641));
  NOR2X1 G16831 (.A1(W4140), .A2(W6298), .ZN(W6315));
  NOR2X1 G16832 (.A1(W34502), .A2(W38698), .ZN(O14552));
  NOR2X1 G16833 (.A1(W21909), .A2(W5843), .ZN(W45858));
  NOR2X1 G16834 (.A1(W2867), .A2(W4920), .ZN(W5643));
  NOR2X1 G16835 (.A1(W23599), .A2(W42999), .ZN(O14033));
  NOR2X1 G16836 (.A1(W9037), .A2(W13085), .ZN(W27087));
  NOR2X1 G16837 (.A1(W22374), .A2(W20398), .ZN(O4132));
  NOR2X1 G16838 (.A1(W3685), .A2(W3414), .ZN(W5099));
  NOR2X1 G16839 (.A1(W620), .A2(W39909), .ZN(O14585));
  NOR2X1 G16840 (.A1(W2402), .A2(I380), .ZN(W6319));
  NOR2X1 G16841 (.A1(W181), .A2(W979), .ZN(W5688));
  NOR2X1 G16842 (.A1(W42655), .A2(W14061), .ZN(O15065));
  NOR2X1 G16843 (.A1(W35932), .A2(W13460), .ZN(O14031));
  NOR2X1 G16844 (.A1(I12), .A2(W7994), .ZN(W23383));
  NOR2X1 G16845 (.A1(W8324), .A2(W5360), .ZN(W23497));
  NOR2X1 G16846 (.A1(W5346), .A2(W43113), .ZN(O14040));
  NOR2X1 G16847 (.A1(W20447), .A2(W28760), .ZN(W45855));
  NOR2X1 G16848 (.A1(W14228), .A2(W1987), .ZN(O2716));
  NOR2X1 G16849 (.A1(W19573), .A2(W18963), .ZN(O14580));
  NOR2X1 G16850 (.A1(W464), .A2(W286), .ZN(W6309));
  NOR2X1 G16851 (.A1(W13142), .A2(I276), .ZN(O14682));
  NOR2X1 G16852 (.A1(W4507), .A2(W2921), .ZN(W6310));
  NOR2X1 G16853 (.A1(W19071), .A2(W25888), .ZN(W27290));
  NOR2X1 G16854 (.A1(W291), .A2(W1944), .ZN(W5859));
  NOR2X1 G16855 (.A1(W3913), .A2(W197), .ZN(W5646));
  NOR2X1 G16856 (.A1(W17743), .A2(W5988), .ZN(O4054));
  NOR2X1 G16857 (.A1(W447), .A2(I1838), .ZN(W5105));
  NOR2X1 G16858 (.A1(W4788), .A2(W18563), .ZN(W27510));
  NOR2X1 G16859 (.A1(I1939), .A2(W3474), .ZN(W5519));
  NOR2X1 G16860 (.A1(W380), .A2(W6342), .ZN(O15062));
  NOR2X1 G16861 (.A1(W59), .A2(W4850), .ZN(W6314));
  NANDX1 G16862 (.A1(W7164), .A2(W10838), .ZN(O3476));
  NANDX1 G16863 (.A1(W1796), .A2(W17427), .ZN(O5167));
  NANDX1 G16864 (.A1(W6251), .A2(W13947), .ZN(O4392));
  NANDX1 G16865 (.A1(W19955), .A2(W2551), .ZN(O3449));
  NANDX1 G16866 (.A1(W7662), .A2(W4838), .ZN(O5809));
  NANDX1 G16867 (.A1(W745), .A2(W27193), .ZN(W31492));
  NANDX1 G16868 (.A1(W27540), .A2(W17909), .ZN(O5805));
  NANDX1 G16869 (.A1(W1114), .A2(W14331), .ZN(W28693));
  NANDX1 G16870 (.A1(W28149), .A2(W1554), .ZN(W29708));
  NANDX1 G16871 (.A1(W11227), .A2(I1778), .ZN(W28193));
  NANDX1 G16872 (.A1(W25056), .A2(W7864), .ZN(W27200));
  NANDX1 G16873 (.A1(W18230), .A2(W19712), .ZN(O3889));
  NANDX1 G16874 (.A1(W17324), .A2(W31056), .ZN(W31490));
  NANDX1 G16875 (.A1(W11862), .A2(W20357), .ZN(W26840));
  NANDX1 G16876 (.A1(W27582), .A2(W19216), .ZN(O4394));
  NANDX1 G16877 (.A1(W3922), .A2(W12445), .ZN(W25635));
  NANDX1 G16878 (.A1(W9802), .A2(W18563), .ZN(W31499));
  NANDX1 G16879 (.A1(W19309), .A2(I655), .ZN(O4017));
  NANDX1 G16880 (.A1(W9178), .A2(W9360), .ZN(W25633));
  NANDX1 G16881 (.A1(W7428), .A2(W4722), .ZN(W26841));
  NANDX1 G16882 (.A1(W15370), .A2(W4201), .ZN(O4393));
  NANDX1 G16883 (.A1(W20743), .A2(W6735), .ZN(W28696));
  NANDX1 G16884 (.A1(W15840), .A2(W13460), .ZN(O4015));
  NANDX1 G16885 (.A1(W20970), .A2(W18378), .ZN(W28698));
  NANDX1 G16886 (.A1(W10252), .A2(W4976), .ZN(W25637));
  NANDX1 G16887 (.A1(W5078), .A2(W808), .ZN(O5012));
  NANDX1 G16888 (.A1(W5822), .A2(I164), .ZN(O3479));
  NANDX1 G16889 (.A1(W15358), .A2(I222), .ZN(W28751));
  NANDX1 G16890 (.A1(W10626), .A2(W20892), .ZN(W25713));
  NANDX1 G16891 (.A1(W3339), .A2(W15304), .ZN(O4369));
  NANDX1 G16892 (.A1(W3340), .A2(W14507), .ZN(W31417));
  NANDX1 G16893 (.A1(W797), .A2(W28619), .ZN(O5777));
  NANDX1 G16894 (.A1(W18501), .A2(W10510), .ZN(W28136));
  NANDX1 G16895 (.A1(W26134), .A2(W24405), .ZN(W31414));
  NANDX1 G16896 (.A1(W22553), .A2(W15947), .ZN(O5775));
  NANDX1 G16897 (.A1(W1622), .A2(W27994), .ZN(O4367));
  NANDX1 G16898 (.A1(W7890), .A2(W12165), .ZN(W26810));
  NANDX1 G16899 (.A1(W9391), .A2(W10170), .ZN(O4365));
  NANDX1 G16900 (.A1(W22873), .A2(W24014), .ZN(W31408));
  NANDX1 G16901 (.A1(W12434), .A2(W19421), .ZN(W29675));
  NANDX1 G16902 (.A1(W20224), .A2(W22055), .ZN(W27243));
  NANDX1 G16903 (.A1(W4673), .A2(W4961), .ZN(W28141));
  NANDX1 G16904 (.A1(W19203), .A2(I781), .ZN(O5190));
  NANDX1 G16905 (.A1(W27128), .A2(W25717), .ZN(W27244));
  NANDX1 G16906 (.A1(W19805), .A2(W12970), .ZN(W25720));
  NANDX1 G16907 (.A1(I579), .A2(W17662), .ZN(O4364));
  NANDX1 G16908 (.A1(W19979), .A2(W16175), .ZN(O4362));
  NANDX1 G16909 (.A1(W10914), .A2(W21495), .ZN(O3505));
  NANDX1 G16910 (.A1(W8857), .A2(W29578), .ZN(O5191));
  NANDX1 G16911 (.A1(W24633), .A2(W18657), .ZN(W25725));
  NANDX1 G16912 (.A1(W1059), .A2(W14327), .ZN(W28755));
  NANDX1 G16913 (.A1(I1582), .A2(W26141), .ZN(O5770));
  NANDX1 G16914 (.A1(W16934), .A2(W10043), .ZN(W30110));
  NANDX1 G16915 (.A1(W9654), .A2(W10763), .ZN(O4994));
  NANDX1 G16916 (.A1(I24), .A2(W1926), .ZN(W28746));
  NANDX1 G16917 (.A1(W11832), .A2(W25942), .ZN(O5787));
  NANDX1 G16918 (.A1(W12907), .A2(W27629), .ZN(O5786));
  NANDX1 G16919 (.A1(W5153), .A2(W28124), .ZN(O5186));
  NANDX1 G16920 (.A1(W10142), .A2(W12474), .ZN(W30089));
  NANDX1 G16921 (.A1(W22842), .A2(W23152), .ZN(O4032));
  NANDX1 G16922 (.A1(W16424), .A2(W25213), .ZN(W30090));
  NANDX1 G16923 (.A1(W23706), .A2(W24121), .ZN(O4603));
  NANDX1 G16924 (.A1(W11449), .A2(W4340), .ZN(O5187));
  NANDX1 G16925 (.A1(W24413), .A2(W17446), .ZN(W31430));
  NANDX1 G16926 (.A1(W17346), .A2(W6813), .ZN(W26816));
  NANDX1 G16927 (.A1(W1407), .A2(W23529), .ZN(W25709));
  NANDX1 G16928 (.A1(W22405), .A2(W15037), .ZN(W30095));
  NANDX1 G16929 (.A1(W1282), .A2(W13994), .ZN(O4035));
  NANDX1 G16930 (.A1(W13976), .A2(W25986), .ZN(W26815));
  NANDX1 G16931 (.A1(W9046), .A2(W10087), .ZN(W26814));
  NANDX1 G16932 (.A1(W19639), .A2(W11838), .ZN(O4375));
  NANDX1 G16933 (.A1(W5065), .A2(W8321), .ZN(W31425));
  NANDX1 G16934 (.A1(W8540), .A2(W18758), .ZN(W30099));
  NANDX1 G16935 (.A1(I1065), .A2(I683), .ZN(W31423));
  NANDX1 G16936 (.A1(W25341), .A2(W17516), .ZN(W26811));
  NANDX1 G16937 (.A1(I1114), .A2(W3104), .ZN(W25711));
  NANDX1 G16938 (.A1(W11197), .A2(W3993), .ZN(O5188));
  NANDX1 G16939 (.A1(W3519), .A2(W7026), .ZN(O5782));
  NANDX1 G16940 (.A1(W2979), .A2(I417), .ZN(W28748));
  NANDX1 G16941 (.A1(W24873), .A2(W23992), .ZN(O5780));
  NANDX1 G16942 (.A1(W26440), .A2(I587), .ZN(W28103));
  NANDX1 G16943 (.A1(W21235), .A2(W2585), .ZN(O4038));
  NANDX1 G16944 (.A1(W8556), .A2(W5709), .ZN(W30118));
  NANDX1 G16945 (.A1(W23112), .A2(W24963), .ZN(W27257));
  NANDX1 G16946 (.A1(W9228), .A2(W27467), .ZN(O5764));
  NANDX1 G16947 (.A1(W22845), .A2(W28305), .ZN(W28771));
  NANDX1 G16948 (.A1(W20334), .A2(W2799), .ZN(W29659));
  NANDX1 G16949 (.A1(W26916), .A2(W8931), .ZN(O5195));
  NANDX1 G16950 (.A1(I1720), .A2(W1913), .ZN(W25738));
  NANDX1 G16951 (.A1(W19082), .A2(W5943), .ZN(O4349));
  NANDX1 G16952 (.A1(W6226), .A2(W15934), .ZN(W28777));
  NANDX1 G16953 (.A1(W8220), .A2(W9419), .ZN(W25741));
  NANDX1 G16954 (.A1(W20911), .A2(W22238), .ZN(W28778));
  NANDX1 G16955 (.A1(I347), .A2(W10058), .ZN(W29658));
  NANDX1 G16956 (.A1(W17565), .A2(I322), .ZN(W30115));
  NANDX1 G16957 (.A1(W24662), .A2(W24268), .ZN(W25744));
  NANDX1 G16958 (.A1(W8973), .A2(W18154), .ZN(W28101));
  NANDX1 G16959 (.A1(W19180), .A2(W6536), .ZN(W28779));
  NANDX1 G16960 (.A1(W19065), .A2(W15218), .ZN(W29656));
  NANDX1 G16961 (.A1(W11173), .A2(W8539), .ZN(W28099));
  NANDX1 G16962 (.A1(W5580), .A2(W25657), .ZN(W25750));
  NANDX1 G16963 (.A1(W12824), .A2(W8152), .ZN(O3873));
  NANDX1 G16964 (.A1(W25148), .A2(W19851), .ZN(O4042));
  NANDX1 G16965 (.A1(W28743), .A2(W10650), .ZN(W31383));
  NANDX1 G16966 (.A1(W13404), .A2(W4934), .ZN(O4346));
  NANDX1 G16967 (.A1(W17757), .A2(W14258), .ZN(W30127));
  NANDX1 G16968 (.A1(W9125), .A2(W12796), .ZN(W30129));
  NANDX1 G16969 (.A1(W4617), .A2(W9247), .ZN(W28763));
  NANDX1 G16970 (.A1(W11034), .A2(W13815), .ZN(W28758));
  NANDX1 G16971 (.A1(W12067), .A2(W10381), .ZN(O4361));
  NANDX1 G16972 (.A1(W4992), .A2(W5101), .ZN(W29666));
  NANDX1 G16973 (.A1(W1267), .A2(W7444), .ZN(W30112));
  NANDX1 G16974 (.A1(W11466), .A2(W3736), .ZN(O4357));
  NANDX1 G16975 (.A1(I224), .A2(W15693), .ZN(W28760));
  NANDX1 G16976 (.A1(W30859), .A2(W4481), .ZN(O5769));
  NANDX1 G16977 (.A1(W3453), .A2(W21383), .ZN(W28761));
  NANDX1 G16978 (.A1(W26095), .A2(W10079), .ZN(O4036));
  NANDX1 G16979 (.A1(W25723), .A2(W16086), .ZN(W27251));
  NANDX1 G16980 (.A1(W9100), .A2(W31286), .ZN(O5768));
  NANDX1 G16981 (.A1(W9059), .A2(W7714), .ZN(W28762));
  NANDX1 G16982 (.A1(W25519), .A2(W5481), .ZN(W25705));
  NANDX1 G16983 (.A1(W9149), .A2(W11024), .ZN(O5767));
  NANDX1 G16984 (.A1(W2968), .A2(W3963), .ZN(O3878));
  NANDX1 G16985 (.A1(W9768), .A2(W15105), .ZN(W25728));
  NANDX1 G16986 (.A1(W3513), .A2(W23878), .ZN(W25731));
  NANDX1 G16987 (.A1(W27299), .A2(W6931), .ZN(O4355));
  NANDX1 G16988 (.A1(W27220), .A2(W25060), .ZN(O4607));
  NANDX1 G16989 (.A1(W3459), .A2(W17402), .ZN(W25732));
  NANDX1 G16990 (.A1(W13320), .A2(W22890), .ZN(W25733));
  NANDX1 G16991 (.A1(W4269), .A2(W18216), .ZN(O3877));
  NANDX1 G16992 (.A1(W22820), .A2(W10795), .ZN(W28115));
  NANDX1 G16993 (.A1(W22333), .A2(W4810), .ZN(W25736));
  NANDX1 G16994 (.A1(W11948), .A2(W26370), .ZN(W26801));
  NANDX1 G16995 (.A1(W20115), .A2(W6237), .ZN(W26827));
  NANDX1 G16996 (.A1(W12173), .A2(W4497), .ZN(W28177));
  NANDX1 G16997 (.A1(W18742), .A2(W12360), .ZN(W31466));
  NANDX1 G16998 (.A1(I232), .A2(W18355), .ZN(W25657));
  NANDX1 G16999 (.A1(W26704), .A2(W24583), .ZN(W31465));
  NANDX1 G17000 (.A1(W23388), .A2(W5963), .ZN(O3485));
  NANDX1 G17001 (.A1(W423), .A2(W3903), .ZN(W29697));
  NANDX1 G17002 (.A1(W26556), .A2(W13831), .ZN(W26829));
  NANDX1 G17003 (.A1(W5990), .A2(W26770), .ZN(W28176));
  NANDX1 G17004 (.A1(W20496), .A2(W18030), .ZN(W30054));
  NANDX1 G17005 (.A1(W6924), .A2(W21881), .ZN(W25661));
  NANDX1 G17006 (.A1(W14298), .A2(I1563), .ZN(W27216));
  NANDX1 G17007 (.A1(W16317), .A2(W16537), .ZN(W27217));
  NANDX1 G17008 (.A1(I440), .A2(W26759), .ZN(W31462));
  NANDX1 G17009 (.A1(W14399), .A2(W18417), .ZN(O4025));
  NANDX1 G17010 (.A1(W10119), .A2(W9668), .ZN(W25663));
  NANDX1 G17011 (.A1(W5660), .A2(W22112), .ZN(O5006));
  NANDX1 G17012 (.A1(W2209), .A2(W14927), .ZN(W28719));
  NANDX1 G17013 (.A1(W20709), .A2(W1975), .ZN(W25667));
  NANDX1 G17014 (.A1(W10344), .A2(W1194), .ZN(O5797));
  NANDX1 G17015 (.A1(W31452), .A2(W14518), .ZN(O5796));
  NANDX1 G17016 (.A1(W1414), .A2(W6774), .ZN(O3884));
  NANDX1 G17017 (.A1(W2207), .A2(W3408), .ZN(W26823));
  NANDX1 G17018 (.A1(W26136), .A2(W16231), .ZN(O5795));
  NANDX1 G17019 (.A1(W505), .A2(W17030), .ZN(W26822));
  NANDX1 G17020 (.A1(W27355), .A2(W21321), .ZN(W28174));
  NANDX1 G17021 (.A1(W9216), .A2(W26135), .ZN(O5174));
  NANDX1 G17022 (.A1(W23122), .A2(W1527), .ZN(W26832));
  NANDX1 G17023 (.A1(W24151), .A2(I674), .ZN(O5011));
  NANDX1 G17024 (.A1(W24265), .A2(W13986), .ZN(W27202));
  NANDX1 G17025 (.A1(W2857), .A2(W14246), .ZN(W30047));
  NANDX1 G17026 (.A1(W8264), .A2(W9408), .ZN(O4391));
  NANDX1 G17027 (.A1(W19670), .A2(W8866), .ZN(W26836));
  NANDX1 G17028 (.A1(W21269), .A2(W22201), .ZN(W28705));
  NANDX1 G17029 (.A1(W11269), .A2(I1075), .ZN(W31474));
  NANDX1 G17030 (.A1(W23857), .A2(W20597), .ZN(W27203));
  NANDX1 G17031 (.A1(W4248), .A2(W3539), .ZN(W28706));
  NANDX1 G17032 (.A1(W20448), .A2(W16419), .ZN(W28707));
  NANDX1 G17033 (.A1(W21925), .A2(W28220), .ZN(W28708));
  NANDX1 G17034 (.A1(W5588), .A2(W4121), .ZN(W26834));
  NANDX1 G17035 (.A1(W13741), .A2(W3804), .ZN(W28726));
  NANDX1 G17036 (.A1(W582), .A2(W7236), .ZN(W28713));
  NANDX1 G17037 (.A1(W19121), .A2(W15546), .ZN(O4587));
  NANDX1 G17038 (.A1(W11864), .A2(W29409), .ZN(W31473));
  NANDX1 G17039 (.A1(W21898), .A2(W19090), .ZN(W28715));
  NANDX1 G17040 (.A1(W8345), .A2(W18505), .ZN(W25650));
  NANDX1 G17041 (.A1(W15111), .A2(W19656), .ZN(W26831));
  NANDX1 G17042 (.A1(W10670), .A2(W8026), .ZN(O4588));
  NANDX1 G17043 (.A1(W26848), .A2(W16175), .ZN(W31471));
  NANDX1 G17044 (.A1(W5467), .A2(W5306), .ZN(O5168));
  NANDX1 G17045 (.A1(W16339), .A2(W2522), .ZN(W31470));
  NANDX1 G17046 (.A1(W8071), .A2(W18201), .ZN(W25656));
  NANDX1 G17047 (.A1(W14516), .A2(W25053), .ZN(W29700));
  NANDX1 G17048 (.A1(W25152), .A2(W4431), .ZN(O5183));
  NANDX1 G17049 (.A1(W21674), .A2(W9663), .ZN(O4595));
  NANDX1 G17050 (.A1(W17715), .A2(W18200), .ZN(W25693));
  NANDX1 G17051 (.A1(W13000), .A2(W2011), .ZN(W28162));
  NANDX1 G17052 (.A1(W7353), .A2(W25249), .ZN(O5000));
  NANDX1 G17053 (.A1(W17800), .A2(W16553), .ZN(W30069));
  NANDX1 G17054 (.A1(W23436), .A2(W25855), .ZN(W30071));
  NANDX1 G17055 (.A1(W15712), .A2(W17297), .ZN(O5178));
  NANDX1 G17056 (.A1(W362), .A2(W17999), .ZN(W27233));
  NANDX1 G17057 (.A1(W24279), .A2(W6168), .ZN(O5180));
  NANDX1 G17058 (.A1(W14952), .A2(W15508), .ZN(O5181));
  NANDX1 G17059 (.A1(W25530), .A2(W28543), .ZN(W30078));
  NANDX1 G17060 (.A1(W14923), .A2(W29603), .ZN(W31441));
  NANDX1 G17061 (.A1(W6841), .A2(W23980), .ZN(W29684));
  NANDX1 G17062 (.A1(W8721), .A2(W14421), .ZN(W27234));
  NANDX1 G17063 (.A1(W2260), .A2(W17951), .ZN(W25696));
  NANDX1 G17064 (.A1(I802), .A2(W5610), .ZN(O4599));
  NANDX1 G17065 (.A1(W26439), .A2(W6315), .ZN(O5184));
  NANDX1 G17066 (.A1(W11550), .A2(W470), .ZN(W30082));
  NANDX1 G17067 (.A1(W5382), .A2(W19434), .ZN(W28159));
  NANDX1 G17068 (.A1(W22675), .A2(W9973), .ZN(W29680));
  NANDX1 G17069 (.A1(W7378), .A2(W22399), .ZN(W26817));
  NANDX1 G17070 (.A1(W10741), .A2(W1333), .ZN(W28158));
  NANDX1 G17071 (.A1(W12513), .A2(W1667), .ZN(O4031));
  NANDX1 G17072 (.A1(W16038), .A2(W6349), .ZN(W27239));
  NANDX1 G17073 (.A1(I958), .A2(W20238), .ZN(W31434));
  NANDX1 G17074 (.A1(W23356), .A2(W17212), .ZN(O4382));
  NANDX1 G17075 (.A1(W23735), .A2(W7953), .ZN(W30061));
  NANDX1 G17076 (.A1(W7672), .A2(W11810), .ZN(W25669));
  NANDX1 G17077 (.A1(W3782), .A2(W11738), .ZN(O5794));
  NANDX1 G17078 (.A1(W6098), .A2(W4970), .ZN(W26821));
  NANDX1 G17079 (.A1(W17154), .A2(W21985), .ZN(O5004));
  NANDX1 G17080 (.A1(W19343), .A2(I665), .ZN(O3491));
  NANDX1 G17081 (.A1(I843), .A2(W10019), .ZN(W27223));
  NANDX1 G17082 (.A1(W18759), .A2(W22718), .ZN(O4383));
  NANDX1 G17083 (.A1(W13019), .A2(W30556), .ZN(W31454));
  NANDX1 G17084 (.A1(W28365), .A2(W909), .ZN(O5793));
  NANDX1 G17085 (.A1(W6565), .A2(W14570), .ZN(O3492));
  NANDX1 G17086 (.A1(W16189), .A2(W8854), .ZN(O5177));
  NANDX1 G17087 (.A1(W5228), .A2(W19407), .ZN(W28702));
  NANDX1 G17088 (.A1(W27516), .A2(W21957), .ZN(W31451));
  NANDX1 G17089 (.A1(W17712), .A2(W4266), .ZN(O5792));
  NANDX1 G17090 (.A1(W9733), .A2(W20787), .ZN(O5003));
  NANDX1 G17091 (.A1(W22266), .A2(W14880), .ZN(W26820));
  NANDX1 G17092 (.A1(W25774), .A2(W13843), .ZN(O4028));
  NANDX1 G17093 (.A1(W388), .A2(W18530), .ZN(W25681));
  NANDX1 G17094 (.A1(W1526), .A2(I767), .ZN(W27226));
  NANDX1 G17095 (.A1(W12343), .A2(W18565), .ZN(O4380));
  NANDX1 G17096 (.A1(W12311), .A2(W14035), .ZN(W25684));
  NANDX1 G17097 (.A1(W4767), .A2(W24697), .ZN(W27228));
  NANDX1 G17098 (.A1(W9147), .A2(W25407), .ZN(W25687));
  NANDX1 G17099 (.A1(W6045), .A2(I1546), .ZN(W31448));
  NANDX1 G17100 (.A1(W2829), .A2(W20241), .ZN(W27092));
  NANDX1 G17101 (.A1(W28677), .A2(W17976), .ZN(O5917));
  NANDX1 G17102 (.A1(W8669), .A2(W10847), .ZN(W26990));
  NANDX1 G17103 (.A1(W22830), .A2(W12267), .ZN(O3423));
  NANDX1 G17104 (.A1(W11692), .A2(I1398), .ZN(W28322));
  NANDX1 G17105 (.A1(W16340), .A2(W17944), .ZN(O4449));
  NANDX1 G17106 (.A1(W4252), .A2(W13969), .ZN(W26991));
  NANDX1 G17107 (.A1(W917), .A2(W847), .ZN(O5111));
  NANDX1 G17108 (.A1(W10276), .A2(W21364), .ZN(W28329));
  NANDX1 G17109 (.A1(W7327), .A2(W15596), .ZN(O5056));
  NANDX1 G17110 (.A1(W21658), .A2(W8512), .ZN(W28505));
  NANDX1 G17111 (.A1(W17935), .A2(I680), .ZN(W27090));
  NANDX1 G17112 (.A1(I1780), .A2(W8581), .ZN(W25432));
  NANDX1 G17113 (.A1(W13743), .A2(W620), .ZN(W28498));
  NANDX1 G17114 (.A1(W19467), .A2(W3150), .ZN(O3418));
  NANDX1 G17115 (.A1(W26978), .A2(W13047), .ZN(W31739));
  NANDX1 G17116 (.A1(W1272), .A2(I1763), .ZN(W28496));
  NANDX1 G17117 (.A1(W24267), .A2(W18036), .ZN(W25427));
  NANDX1 G17118 (.A1(W23280), .A2(W24137), .ZN(O5921));
  NANDX1 G17119 (.A1(W2653), .A2(W21730), .ZN(W27094));
  NANDX1 G17120 (.A1(W20530), .A2(I640), .ZN(O3427));
  NANDX1 G17121 (.A1(W7287), .A2(W20702), .ZN(W28513));
  NANDX1 G17122 (.A1(W11998), .A2(W11695), .ZN(W29808));
  NANDX1 G17123 (.A1(W10182), .A2(W11184), .ZN(W28318));
  NANDX1 G17124 (.A1(W17736), .A2(W3586), .ZN(W31730));
  NANDX1 G17125 (.A1(W3788), .A2(W7442), .ZN(W26983));
  NANDX1 G17126 (.A1(W16875), .A2(I1253), .ZN(O4523));
  NANDX1 G17127 (.A1(W17990), .A2(W15928), .ZN(W25447));
  NANDX1 G17128 (.A1(W11948), .A2(W15817), .ZN(W28510));
  NANDX1 G17129 (.A1(W22522), .A2(W14091), .ZN(O3417));
  NANDX1 G17130 (.A1(W24298), .A2(W27810), .ZN(O4446));
  NANDX1 G17131 (.A1(W28264), .A2(W4341), .ZN(W28509));
  NANDX1 G17132 (.A1(W24254), .A2(W22384), .ZN(W29921));
  NANDX1 G17133 (.A1(W4920), .A2(W26202), .ZN(W28508));
  NANDX1 G17134 (.A1(I759), .A2(W25146), .ZN(O3424));
  NANDX1 G17135 (.A1(W21171), .A2(W27989), .ZN(W29809));
  NANDX1 G17136 (.A1(W18810), .A2(I1570), .ZN(W28507));
  NANDX1 G17137 (.A1(W24697), .A2(W2270), .ZN(W26987));
  NANDX1 G17138 (.A1(W12303), .A2(W4342), .ZN(W25410));
  NANDX1 G17139 (.A1(W16654), .A2(W7037), .ZN(W25414));
  NANDX1 G17140 (.A1(W27757), .A2(W20540), .ZN(O5928));
  NANDX1 G17141 (.A1(W6401), .A2(W16370), .ZN(W27086));
  NANDX1 G17142 (.A1(W16170), .A2(W18306), .ZN(O5930));
  NANDX1 G17143 (.A1(W437), .A2(W879), .ZN(W28487));
  NANDX1 G17144 (.A1(W14439), .A2(W18339), .ZN(O3412));
  NANDX1 G17145 (.A1(W26959), .A2(W24030), .ZN(W29912));
  NANDX1 G17146 (.A1(W3967), .A2(W14072), .ZN(O4518));
  NANDX1 G17147 (.A1(W19404), .A2(W12339), .ZN(W25411));
  NANDX1 G17148 (.A1(W8216), .A2(W26526), .ZN(W28491));
  NANDX1 G17149 (.A1(I1942), .A2(W21512), .ZN(W28485));
  NANDX1 G17150 (.A1(W16056), .A2(W24091), .ZN(O5103));
  NANDX1 G17151 (.A1(W17161), .A2(W27685), .ZN(W28484));
  NANDX1 G17152 (.A1(W25312), .A2(W31682), .ZN(W31761));
  NANDX1 G17153 (.A1(W26679), .A2(W7694), .ZN(W29823));
  NANDX1 G17154 (.A1(W9195), .A2(W17120), .ZN(O3978));
  NANDX1 G17155 (.A1(W22037), .A2(W16373), .ZN(O5101));
  NANDX1 G17156 (.A1(W17511), .A2(W28387), .ZN(W31763));
  NANDX1 G17157 (.A1(W18334), .A2(W7172), .ZN(O4456));
  NANDX1 G17158 (.A1(W11136), .A2(W210), .ZN(W27089));
  NANDX1 G17159 (.A1(W24821), .A2(W26503), .ZN(O5923));
  NANDX1 G17160 (.A1(W27186), .A2(W14076), .ZN(W29915));
  NANDX1 G17161 (.A1(W21149), .A2(W26084), .ZN(O4453));
  NANDX1 G17162 (.A1(W28417), .A2(W19964), .ZN(O5058));
  NANDX1 G17163 (.A1(I54), .A2(W8493), .ZN(O4454));
  NANDX1 G17164 (.A1(W21314), .A2(W22554), .ZN(O4455));
  NANDX1 G17165 (.A1(W28454), .A2(I1340), .ZN(W31751));
  NANDX1 G17166 (.A1(W23055), .A2(W14492), .ZN(W25423));
  NANDX1 G17167 (.A1(W12713), .A2(W20796), .ZN(O3428));
  NANDX1 G17168 (.A1(W26957), .A2(W1562), .ZN(O4521));
  NANDX1 G17169 (.A1(W11104), .A2(W1064), .ZN(O5926));
  NANDX1 G17170 (.A1(W8781), .A2(W18361), .ZN(O4459));
  NANDX1 G17171 (.A1(W6439), .A2(W2674), .ZN(W25421));
  NANDX1 G17172 (.A1(W19012), .A2(W23159), .ZN(W28348));
  NANDX1 G17173 (.A1(W877), .A2(W17604), .ZN(W31754));
  NANDX1 G17174 (.A1(W6410), .A2(W18076), .ZN(W28351));
  NANDX1 G17175 (.A1(W520), .A2(W18329), .ZN(W25416));
  NANDX1 G17176 (.A1(W15686), .A2(W20276), .ZN(O5903));
  NANDX1 G17177 (.A1(W22889), .A2(W1399), .ZN(O3941));
  NANDX1 G17178 (.A1(W25637), .A2(W23497), .ZN(O3942));
  NANDX1 G17179 (.A1(W17618), .A2(W24779), .ZN(W27108));
  NANDX1 G17180 (.A1(W6214), .A2(W18302), .ZN(W31703));
  NANDX1 G17181 (.A1(W31441), .A2(W25492), .ZN(W31704));
  NANDX1 G17182 (.A1(W10534), .A2(W28647), .ZN(O5052));
  NANDX1 G17183 (.A1(W6859), .A2(W8566), .ZN(W25472));
  NANDX1 G17184 (.A1(W16572), .A2(W14316), .ZN(W25471));
  NANDX1 G17185 (.A1(W8796), .A2(W1151), .ZN(W28293));
  NANDX1 G17186 (.A1(W13557), .A2(W11928), .ZN(O3985));
  NANDX1 G17187 (.A1(W15977), .A2(W18484), .ZN(W26959));
  NANDX1 G17188 (.A1(W25140), .A2(W12704), .ZN(W31708));
  NANDX1 G17189 (.A1(W25635), .A2(W25938), .ZN(O5904));
  NANDX1 G17190 (.A1(W22035), .A2(W10686), .ZN(O3983));
  NANDX1 G17191 (.A1(W1597), .A2(W9285), .ZN(O4530));
  NANDX1 G17192 (.A1(W23046), .A2(W20187), .ZN(W28294));
  NANDX1 G17193 (.A1(W25653), .A2(W28802), .ZN(W31711));
  NANDX1 G17194 (.A1(W5965), .A2(W7942), .ZN(O4435));
  NANDX1 G17195 (.A1(W2991), .A2(W23649), .ZN(O3431));
  NANDX1 G17196 (.A1(W775), .A2(W13585), .ZN(W25487));
  NANDX1 G17197 (.A1(W26856), .A2(W4349), .ZN(W28545));
  NANDX1 G17198 (.A1(W14998), .A2(W12001), .ZN(W29943));
  NANDX1 G17199 (.A1(W18776), .A2(I1868), .ZN(W25484));
  NANDX1 G17200 (.A1(W9439), .A2(W2507), .ZN(O5049));
  NANDX1 G17201 (.A1(W23553), .A2(W12707), .ZN(O3432));
  NANDX1 G17202 (.A1(I72), .A2(W8569), .ZN(W25478));
  NANDX1 G17203 (.A1(W10333), .A2(W1050), .ZN(O5118));
  NANDX1 G17204 (.A1(W23504), .A2(W15556), .ZN(O3989));
  NANDX1 G17205 (.A1(W92), .A2(W8082), .ZN(W26960));
  NANDX1 G17206 (.A1(W5738), .A2(W25186), .ZN(W31700));
  NANDX1 G17207 (.A1(W25601), .A2(W18851), .ZN(W28540));
  NANDX1 G17208 (.A1(W23723), .A2(W16677), .ZN(O4535));
  NANDX1 G17209 (.A1(W947), .A2(W15439), .ZN(O3940));
  NANDX1 G17210 (.A1(W8552), .A2(W22518), .ZN(W26954));
  NANDX1 G17211 (.A1(W8994), .A2(W732), .ZN(O3987));
  NANDX1 G17212 (.A1(W27840), .A2(W20024), .ZN(O4534));
  NANDX1 G17213 (.A1(W27037), .A2(W15379), .ZN(W28536));
  NANDX1 G17214 (.A1(W14759), .A2(W19155), .ZN(O5112));
  NANDX1 G17215 (.A1(I1560), .A2(W6117), .ZN(O5114));
  NANDX1 G17216 (.A1(W21981), .A2(W18852), .ZN(O4440));
  NANDX1 G17217 (.A1(W17906), .A2(W19058), .ZN(W25460));
  NANDX1 G17218 (.A1(W3452), .A2(W11641), .ZN(O3429));
  NANDX1 G17219 (.A1(W12411), .A2(W17234), .ZN(O3948));
  NANDX1 G17220 (.A1(W15403), .A2(I1825), .ZN(W26973));
  NANDX1 G17221 (.A1(W23589), .A2(W21691), .ZN(W28314));
  NANDX1 G17222 (.A1(W17672), .A2(I1940), .ZN(W28518));
  NANDX1 G17223 (.A1(W3837), .A2(W15478), .ZN(W28315));
  NANDX1 G17224 (.A1(I1754), .A2(W751), .ZN(O5912));
  NANDX1 G17225 (.A1(W20210), .A2(W24352), .ZN(W26975));
  NANDX1 G17226 (.A1(W12083), .A2(W8750), .ZN(W29922));
  NANDX1 G17227 (.A1(W9999), .A2(W25411), .ZN(W27102));
  NANDX1 G17228 (.A1(W193), .A2(W14746), .ZN(W26978));
  NANDX1 G17229 (.A1(W16118), .A2(W23374), .ZN(W25457));
  NANDX1 G17230 (.A1(W9800), .A2(W16151), .ZN(O4444));
  NANDX1 G17231 (.A1(W17591), .A2(W12479), .ZN(W27098));
  NANDX1 G17232 (.A1(W3742), .A2(W26364), .ZN(O5914));
  NANDX1 G17233 (.A1(W27643), .A2(W1165), .ZN(O4439));
  NANDX1 G17234 (.A1(W12521), .A2(W8788), .ZN(O4438));
  NANDX1 G17235 (.A1(W214), .A2(W19205), .ZN(W26962));
  NANDX1 G17236 (.A1(W15312), .A2(W5708), .ZN(W29804));
  NANDX1 G17237 (.A1(W15451), .A2(W13016), .ZN(W29934));
  NANDX1 G17238 (.A1(I49), .A2(W24958), .ZN(W28306));
  NANDX1 G17239 (.A1(W13292), .A2(I1411), .ZN(W27103));
  NANDX1 G17240 (.A1(W20606), .A2(W14124), .ZN(O3430));
  NANDX1 G17241 (.A1(W8781), .A2(W20180), .ZN(W28308));
  NANDX1 G17242 (.A1(W23009), .A2(W27648), .ZN(W31764));
  NANDX1 G17243 (.A1(W12528), .A2(W23119), .ZN(W25467));
  NANDX1 G17244 (.A1(W21269), .A2(W12203), .ZN(W28522));
  NANDX1 G17245 (.A1(W6054), .A2(W7920), .ZN(W26967));
  NANDX1 G17246 (.A1(W10311), .A2(W5534), .ZN(W29932));
  NANDX1 G17247 (.A1(I960), .A2(W16956), .ZN(W31719));
  NANDX1 G17248 (.A1(W6171), .A2(W20234), .ZN(O3947));
  NANDX1 G17249 (.A1(W11569), .A2(W16843), .ZN(W25463));
  NANDX1 G17250 (.A1(W14776), .A2(W19509), .ZN(W31721));
  NANDX1 G17251 (.A1(W12018), .A2(W19745), .ZN(W25367));
  NANDX1 G17252 (.A1(W26669), .A2(W2505), .ZN(W28397));
  NANDX1 G17253 (.A1(W7325), .A2(W17408), .ZN(W25369));
  NANDX1 G17254 (.A1(W3549), .A2(W10553), .ZN(O5092));
  NANDX1 G17255 (.A1(W20290), .A2(W21810), .ZN(W27033));
  NANDX1 G17256 (.A1(W17549), .A2(I932), .ZN(W31811));
  NANDX1 G17257 (.A1(W21792), .A2(W26415), .ZN(W29855));
  NANDX1 G17258 (.A1(W19474), .A2(W6855), .ZN(O5081));
  NANDX1 G17259 (.A1(W4126), .A2(I24), .ZN(W27054));
  NANDX1 G17260 (.A1(W23572), .A2(W15906), .ZN(O4483));
  NANDX1 G17261 (.A1(W5692), .A2(I1127), .ZN(O4481));
  NANDX1 G17262 (.A1(W6085), .A2(W26453), .ZN(W28405));
  NANDX1 G17263 (.A1(W27554), .A2(W5399), .ZN(O4502));
  NANDX1 G17264 (.A1(W14840), .A2(W19527), .ZN(W27035));
  NANDX1 G17265 (.A1(W18976), .A2(W22924), .ZN(O3970));
  NANDX1 G17266 (.A1(W26644), .A2(W12379), .ZN(W27052));
  NANDX1 G17267 (.A1(W25185), .A2(W18775), .ZN(W29875));
  NANDX1 G17268 (.A1(W16493), .A2(W27445), .ZN(O5090));
  NANDX1 G17269 (.A1(W5077), .A2(W4065), .ZN(W28440));
  NANDX1 G17270 (.A1(W16840), .A2(I946), .ZN(W27026));
  NANDX1 G17271 (.A1(W23782), .A2(W17385), .ZN(O3394));
  NANDX1 G17272 (.A1(W17370), .A2(W30086), .ZN(W31803));
  NANDX1 G17273 (.A1(W20620), .A2(W26235), .ZN(W29845));
  NANDX1 G17274 (.A1(W26409), .A2(W11427), .ZN(W29883));
  NANDX1 G17275 (.A1(W28915), .A2(W4836), .ZN(W31805));
  NANDX1 G17276 (.A1(W8068), .A2(W24535), .ZN(W28453));
  NANDX1 G17277 (.A1(W18609), .A2(W7350), .ZN(O3393));
  NANDX1 G17278 (.A1(W3209), .A2(W12096), .ZN(W27024));
  NANDX1 G17279 (.A1(W20), .A2(W16945), .ZN(W27060));
  NANDX1 G17280 (.A1(I1751), .A2(W11143), .ZN(O3969));
  NANDX1 G17281 (.A1(W26861), .A2(W22263), .ZN(W27059));
  NANDX1 G17282 (.A1(I1141), .A2(W7193), .ZN(W28451));
  NANDX1 G17283 (.A1(W11678), .A2(W12846), .ZN(W27027));
  NANDX1 G17284 (.A1(W10231), .A2(W3174), .ZN(O4480));
  NANDX1 G17285 (.A1(W3185), .A2(W75), .ZN(W29846));
  NANDX1 G17286 (.A1(W6410), .A2(W8654), .ZN(W25371));
  NANDX1 G17287 (.A1(W189), .A2(W19358), .ZN(O5077));
  NANDX1 G17288 (.A1(W11066), .A2(W5390), .ZN(O5958));
  NANDX1 G17289 (.A1(W25893), .A2(W15149), .ZN(W28426));
  NANDX1 G17290 (.A1(W25470), .A2(W2145), .ZN(O4489));
  NANDX1 G17291 (.A1(W2238), .A2(W5879), .ZN(W28428));
  NANDX1 G17292 (.A1(W9817), .A2(W3871), .ZN(O4490));
  NANDX1 G17293 (.A1(W20779), .A2(W5254), .ZN(W25354));
  NANDX1 G17294 (.A1(W98), .A2(W5461), .ZN(W25353));
  NANDX1 G17295 (.A1(W16136), .A2(W11132), .ZN(W25351));
  NANDX1 G17296 (.A1(W3934), .A2(W12079), .ZN(W31822));
  NANDX1 G17297 (.A1(W20466), .A2(W14940), .ZN(O3968));
  NANDX1 G17298 (.A1(W17400), .A2(W17639), .ZN(W27048));
  NANDX1 G17299 (.A1(W19337), .A2(W19530), .ZN(W27041));
  NANDX1 G17300 (.A1(W17342), .A2(W4791), .ZN(O5085));
  NANDX1 G17301 (.A1(W8994), .A2(W22842), .ZN(O5086));
  NANDX1 G17302 (.A1(W21852), .A2(W13020), .ZN(W25347));
  NANDX1 G17303 (.A1(W13203), .A2(W3164), .ZN(W25346));
  NANDX1 G17304 (.A1(W2670), .A2(W1612), .ZN(O4494));
  NANDX1 G17305 (.A1(W22591), .A2(W19282), .ZN(W28423));
  NANDX1 G17306 (.A1(W6179), .A2(W5213), .ZN(O4493));
  NANDX1 G17307 (.A1(W10827), .A2(W10566), .ZN(O5413));
  NANDX1 G17308 (.A1(W31051), .A2(W24281), .ZN(O5961));
  NANDX1 G17309 (.A1(W14139), .A2(W3090), .ZN(W31815));
  NANDX1 G17310 (.A1(W11972), .A2(W17385), .ZN(O4486));
  NANDX1 G17311 (.A1(W3809), .A2(W24068), .ZN(W28435));
  NANDX1 G17312 (.A1(W3370), .A2(W2397), .ZN(W25362));
  NANDX1 G17313 (.A1(W695), .A2(W12970), .ZN(W27038));
  NANDX1 G17314 (.A1(W16032), .A2(W18727), .ZN(O4498));
  NANDX1 G17315 (.A1(W27984), .A2(W2547), .ZN(W28433));
  NANDX1 G17316 (.A1(W9289), .A2(W27059), .ZN(W29873));
  NANDX1 G17317 (.A1(W16942), .A2(W21087), .ZN(W31801));
  NANDX1 G17318 (.A1(W11590), .A2(W23439), .ZN(O4487));
  NANDX1 G17319 (.A1(W12825), .A2(W18933), .ZN(O4488));
  NANDX1 G17320 (.A1(W916), .A2(W21343), .ZN(W31819));
  NANDX1 G17321 (.A1(W10430), .A2(W11861), .ZN(O4497));
  NANDX1 G17322 (.A1(W28774), .A2(W12311), .ZN(O5083));
  NANDX1 G17323 (.A1(W628), .A2(W25484), .ZN(W28431));
  NANDX1 G17324 (.A1(W2956), .A2(W23921), .ZN(W25358));
  NANDX1 G17325 (.A1(W24986), .A2(W10722), .ZN(O3387));
  NANDX1 G17326 (.A1(W19152), .A2(W18993), .ZN(W29893));
  NANDX1 G17327 (.A1(W14981), .A2(W13302), .ZN(W29899));
  NANDX1 G17328 (.A1(I1724), .A2(W27834), .ZN(O5940));
  NANDX1 G17329 (.A1(W20580), .A2(W5556), .ZN(W28370));
  NANDX1 G17330 (.A1(W2398), .A2(W15942), .ZN(W28371));
  NANDX1 G17331 (.A1(W17010), .A2(W10655), .ZN(O3977));
  NANDX1 G17332 (.A1(W20797), .A2(W18471), .ZN(W25390));
  NANDX1 G17333 (.A1(W1299), .A2(W6166), .ZN(W27007));
  NANDX1 G17334 (.A1(I1851), .A2(W24772), .ZN(O5065));
  NANDX1 G17335 (.A1(W765), .A2(W24076), .ZN(O5942));
  NANDX1 G17336 (.A1(W16767), .A2(W11681), .ZN(W31779));
  NANDX1 G17337 (.A1(W12340), .A2(W24894), .ZN(O5067));
  NANDX1 G17338 (.A1(W6123), .A2(W7409), .ZN(W25387));
  NANDX1 G17339 (.A1(W2522), .A2(W26010), .ZN(W31784));
  NANDX1 G17340 (.A1(W24062), .A2(W19264), .ZN(W27078));
  NANDX1 G17341 (.A1(W19719), .A2(W138), .ZN(W28472));
  NANDX1 G17342 (.A1(W24742), .A2(W2475), .ZN(O5943));
  NANDX1 G17343 (.A1(W27557), .A2(W16195), .ZN(O4469));
  NANDX1 G17344 (.A1(W6715), .A2(W24404), .ZN(W27077));
  NANDX1 G17345 (.A1(W25007), .A2(W10095), .ZN(O3406));
  NANDX1 G17346 (.A1(W11355), .A2(I1296), .ZN(W25404));
  NANDX1 G17347 (.A1(W22192), .A2(W19825), .ZN(W28366));
  NANDX1 G17348 (.A1(W21942), .A2(W23907), .ZN(W25402));
  NANDX1 G17349 (.A1(W1872), .A2(W23049), .ZN(W29904));
  NANDX1 G17350 (.A1(W17102), .A2(W29655), .ZN(W29902));
  NANDX1 G17351 (.A1(W10200), .A2(W12878), .ZN(O4517));
  NANDX1 G17352 (.A1(W21107), .A2(W22807), .ZN(W28367));
  NANDX1 G17353 (.A1(W16782), .A2(W1329), .ZN(W31769));
  NANDX1 G17354 (.A1(W10855), .A2(W9742), .ZN(W25400));
  NANDX1 G17355 (.A1(W5671), .A2(W24679), .ZN(W25386));
  NANDX1 G17356 (.A1(W7580), .A2(W10199), .ZN(O3405));
  NANDX1 G17357 (.A1(W808), .A2(W29451), .ZN(W31773));
  NANDX1 G17358 (.A1(W26124), .A2(W26360), .ZN(O5064));
  NANDX1 G17359 (.A1(W4060), .A2(W27999), .ZN(W31775));
  NANDX1 G17360 (.A1(I696), .A2(W12872), .ZN(O5937));
  NANDX1 G17361 (.A1(W11322), .A2(W27504), .ZN(O5099));
  NANDX1 G17362 (.A1(W6301), .A2(W9966), .ZN(O3404));
  NANDX1 G17363 (.A1(W23145), .A2(W20256), .ZN(W28479));
  NANDX1 G17364 (.A1(W29680), .A2(W15846), .ZN(W31796));
  NANDX1 G17365 (.A1(W3446), .A2(W9219), .ZN(W29836));
  NANDX1 G17366 (.A1(W16524), .A2(W17126), .ZN(O5948));
  NANDX1 G17367 (.A1(W21582), .A2(W8618), .ZN(O5073));
  NANDX1 G17368 (.A1(W23956), .A2(W18367), .ZN(O3974));
  NANDX1 G17369 (.A1(W24912), .A2(I1365), .ZN(O3960));
  NANDX1 G17370 (.A1(W4229), .A2(W15588), .ZN(W27019));
  NANDX1 G17371 (.A1(W1754), .A2(W12757), .ZN(O4475));
  NANDX1 G17372 (.A1(W18817), .A2(W14417), .ZN(W29887));
  NANDX1 G17373 (.A1(I1002), .A2(W26713), .ZN(W27021));
  NANDX1 G17374 (.A1(W16262), .A2(W27057), .ZN(W27070));
  NANDX1 G17375 (.A1(W15474), .A2(W2922), .ZN(W28459));
  NANDX1 G17376 (.A1(W15070), .A2(W6514), .ZN(W27068));
  NANDX1 G17377 (.A1(W19902), .A2(W21795), .ZN(W28389));
  NANDX1 G17378 (.A1(W4068), .A2(W23327), .ZN(O4479));
  NANDX1 G17379 (.A1(W5965), .A2(W16901), .ZN(O5952));
  NANDX1 G17380 (.A1(I475), .A2(W309), .ZN(O3961));
  NANDX1 G17381 (.A1(W2208), .A2(W24491), .ZN(W28454));
  NANDX1 G17382 (.A1(W20093), .A2(W14901), .ZN(O3972));
  NANDX1 G17383 (.A1(W1758), .A2(W13552), .ZN(O4470));
  NANDX1 G17384 (.A1(W22178), .A2(W19150), .ZN(W29832));
  NANDX1 G17385 (.A1(W4034), .A2(W2025), .ZN(W31789));
  NANDX1 G17386 (.A1(W23721), .A2(W5253), .ZN(O3401));
  NANDX1 G17387 (.A1(W11768), .A2(W5747), .ZN(O3397));
  NANDX1 G17388 (.A1(W8828), .A2(W15502), .ZN(O4514));
  NANDX1 G17389 (.A1(W5584), .A2(W26952), .ZN(W28375));
  NANDX1 G17390 (.A1(W1311), .A2(W23493), .ZN(O5946));
  NANDX1 G17391 (.A1(W18390), .A2(W11418), .ZN(W25379));
  NANDX1 G17392 (.A1(W17833), .A2(W25652), .ZN(O3991));
  NANDX1 G17393 (.A1(W1373), .A2(W19481), .ZN(O3396));
  NANDX1 G17394 (.A1(W2820), .A2(W27622), .ZN(W29891));
  NANDX1 G17395 (.A1(W25211), .A2(W27682), .ZN(W31792));
  NANDX1 G17396 (.A1(W17145), .A2(W14836), .ZN(O4473));
  NANDX1 G17397 (.A1(W1113), .A2(W14215), .ZN(O3959));
  NANDX1 G17398 (.A1(W4675), .A2(W24049), .ZN(W27075));
  NANDX1 G17399 (.A1(W7660), .A2(W22318), .ZN(W27072));
  NANDX1 G17400 (.A1(W9552), .A2(W16958), .ZN(W29890));
  NANDX1 G17401 (.A1(W14019), .A2(I616), .ZN(O3458));
  NANDX1 G17402 (.A1(W16708), .A2(W16121), .ZN(W25568));
  NANDX1 G17403 (.A1(W20860), .A2(W11210), .ZN(W26879));
  NANDX1 G17404 (.A1(I1889), .A2(W23965), .ZN(O5837));
  NANDX1 G17405 (.A1(W5665), .A2(W10295), .ZN(W30016));
  NANDX1 G17406 (.A1(W277), .A2(W2673), .ZN(O5154));
  NANDX1 G17407 (.A1(W27182), .A2(W4025), .ZN(O5153));
  NANDX1 G17408 (.A1(W3324), .A2(W5447), .ZN(W30012));
  NANDX1 G17409 (.A1(W7654), .A2(W4579), .ZN(W28227));
  NANDX1 G17410 (.A1(W12857), .A2(W14458), .ZN(W31555));
  NANDX1 G17411 (.A1(W19609), .A2(W2303), .ZN(W27167));
  NANDX1 G17412 (.A1(W18491), .A2(W27326), .ZN(W28646));
  NANDX1 G17413 (.A1(W245), .A2(W7381), .ZN(W27166));
  NANDX1 G17414 (.A1(W16281), .A2(W27074), .ZN(O5022));
  NANDX1 G17415 (.A1(W9501), .A2(W15164), .ZN(W31562));
  NANDX1 G17416 (.A1(W7941), .A2(W5626), .ZN(W31566));
  NANDX1 G17417 (.A1(I422), .A2(W6712), .ZN(W27165));
  NANDX1 G17418 (.A1(W90), .A2(W11772), .ZN(O3904));
  NANDX1 G17419 (.A1(W23730), .A2(W80), .ZN(W25562));
  NANDX1 G17420 (.A1(W18288), .A2(W20841), .ZN(W25572));
  NANDX1 G17421 (.A1(W24970), .A2(W11407), .ZN(W31536));
  NANDX1 G17422 (.A1(W14146), .A2(W31362), .ZN(W31537));
  NANDX1 G17423 (.A1(W758), .A2(W2654), .ZN(O4010));
  NANDX1 G17424 (.A1(W21725), .A2(W766), .ZN(W25574));
  NANDX1 G17425 (.A1(W6827), .A2(W17867), .ZN(O3899));
  NANDX1 G17426 (.A1(W1873), .A2(W18425), .ZN(W31544));
  NANDX1 G17427 (.A1(W23337), .A2(W25797), .ZN(O3900));
  NANDX1 G17428 (.A1(W16357), .A2(W18815), .ZN(O3901));
  NANDX1 G17429 (.A1(W22280), .A2(W16997), .ZN(W27171));
  NANDX1 G17430 (.A1(W12573), .A2(W12446), .ZN(O5024));
  NANDX1 G17431 (.A1(W16914), .A2(W2802), .ZN(O5832));
  NANDX1 G17432 (.A1(W20849), .A2(W15234), .ZN(W25570));
  NANDX1 G17433 (.A1(W22880), .A2(W24694), .ZN(W25569));
  NANDX1 G17434 (.A1(W29424), .A2(W19738), .ZN(O5156));
  NANDX1 G17435 (.A1(I607), .A2(W2672), .ZN(W28225));
  NANDX1 G17436 (.A1(W2255), .A2(W19840), .ZN(W30020));
  NANDX1 G17437 (.A1(W29161), .A2(W26059), .ZN(O5833));
  NANDX1 G17438 (.A1(W17780), .A2(I118), .ZN(O5155));
  NANDX1 G17439 (.A1(W5924), .A2(W27542), .ZN(W28629));
  NANDX1 G17440 (.A1(W15827), .A2(W26647), .ZN(O4411));
  NANDX1 G17441 (.A1(W20918), .A2(W8112), .ZN(W29756));
  NANDX1 G17442 (.A1(W11161), .A2(W13698), .ZN(W25550));
  NANDX1 G17443 (.A1(I1229), .A2(W1872), .ZN(O3910));
  NANDX1 G17444 (.A1(W22297), .A2(W16813), .ZN(O9410));
  NANDX1 G17445 (.A1(W8609), .A2(W26820), .ZN(O5030));
  NANDX1 G17446 (.A1(W7001), .A2(I332), .ZN(W25548));
  NANDX1 G17447 (.A1(W472), .A2(W14147), .ZN(O5146));
  NANDX1 G17448 (.A1(W3588), .A2(W21383), .ZN(O5031));
  NANDX1 G17449 (.A1(W21862), .A2(W12062), .ZN(W27157));
  NANDX1 G17450 (.A1(W24812), .A2(W23253), .ZN(W26898));
  NANDX1 G17451 (.A1(W21254), .A2(W28587), .ZN(W28628));
  NANDX1 G17452 (.A1(W8800), .A2(W28738), .ZN(O5849));
  NANDX1 G17453 (.A1(W12356), .A2(W15040), .ZN(O5850));
  NANDX1 G17454 (.A1(W26797), .A2(I1372), .ZN(W31592));
  NANDX1 G17455 (.A1(W19275), .A2(W16838), .ZN(W25545));
  NANDX1 G17456 (.A1(W16373), .A2(W22233), .ZN(W31594));
  NANDX1 G17457 (.A1(W20938), .A2(W5790), .ZN(W28626));
  NANDX1 G17458 (.A1(W3868), .A2(W12956), .ZN(O4005));
  NANDX1 G17459 (.A1(W808), .A2(W11729), .ZN(W28641));
  NANDX1 G17460 (.A1(W31212), .A2(W28152), .ZN(W31567));
  NANDX1 G17461 (.A1(W14897), .A2(W4270), .ZN(O4410));
  NANDX1 G17462 (.A1(W23644), .A2(W18389), .ZN(O5151));
  NANDX1 G17463 (.A1(W26233), .A2(W1692), .ZN(W27161));
  NANDX1 G17464 (.A1(W11319), .A2(W18031), .ZN(O5025));
  NANDX1 G17465 (.A1(W10448), .A2(W20927), .ZN(O5150));
  NANDX1 G17466 (.A1(W29639), .A2(W24957), .ZN(O5026));
  NANDX1 G17467 (.A1(W7310), .A2(W7657), .ZN(O4406));
  NANDX1 G17468 (.A1(W1193), .A2(W25437), .ZN(W28232));
  NANDX1 G17469 (.A1(W6780), .A2(W3133), .ZN(O3909));
  NANDX1 G17470 (.A1(W13946), .A2(W5013), .ZN(W28633));
  NANDX1 G17471 (.A1(W24571), .A2(W11674), .ZN(W25553));
  NANDX1 G17472 (.A1(W1133), .A2(W21736), .ZN(W30001));
  NANDX1 G17473 (.A1(W19732), .A2(W20315), .ZN(W28632));
  NANDX1 G17474 (.A1(W4989), .A2(I454), .ZN(O5845));
  NANDX1 G17475 (.A1(W25476), .A2(I1939), .ZN(W31578));
  NANDX1 G17476 (.A1(W18507), .A2(I1865), .ZN(W25607));
  NANDX1 G17477 (.A1(W26635), .A2(W9151), .ZN(W27182));
  NANDX1 G17478 (.A1(W17709), .A2(W18294), .ZN(O4013));
  NANDX1 G17479 (.A1(W284), .A2(W19501), .ZN(O3469));
  NANDX1 G17480 (.A1(W20963), .A2(W6035), .ZN(O4579));
  NANDX1 G17481 (.A1(W26143), .A2(W9318), .ZN(W28212));
  NANDX1 G17482 (.A1(W9884), .A2(W382), .ZN(W25611));
  NANDX1 G17483 (.A1(W18200), .A2(W3397), .ZN(O3468));
  NANDX1 G17484 (.A1(W22114), .A2(W8035), .ZN(O5161));
  NANDX1 G17485 (.A1(W20439), .A2(W8505), .ZN(W26863));
  NANDX1 G17486 (.A1(W236), .A2(W14456), .ZN(W31509));
  NANDX1 G17487 (.A1(W19591), .A2(I911), .ZN(O4578));
  NANDX1 G17488 (.A1(W6835), .A2(W9711), .ZN(W25605));
  NANDX1 G17489 (.A1(W15361), .A2(I1709), .ZN(W26864));
  NANDX1 G17490 (.A1(W19449), .A2(W1214), .ZN(O3465));
  NANDX1 G17491 (.A1(W5982), .A2(W11651), .ZN(W26866));
  NANDX1 G17492 (.A1(W17644), .A2(W143), .ZN(W28214));
  NANDX1 G17493 (.A1(W26568), .A2(W20753), .ZN(W28676));
  NANDX1 G17494 (.A1(W12356), .A2(W17416), .ZN(W27180));
  NANDX1 G17495 (.A1(W2339), .A2(W26211), .ZN(W27188));
  NANDX1 G17496 (.A1(W10852), .A2(W16410), .ZN(W25631));
  NANDX1 G17497 (.A1(W24288), .A2(W20211), .ZN(W28205));
  NANDX1 G17498 (.A1(W15759), .A2(W19825), .ZN(O4399));
  NANDX1 G17499 (.A1(W7455), .A2(W5212), .ZN(W25630));
  NANDX1 G17500 (.A1(W22633), .A2(W4984), .ZN(W26849));
  NANDX1 G17501 (.A1(W15937), .A2(W19759), .ZN(W25628));
  NANDX1 G17502 (.A1(W23853), .A2(W29484), .ZN(W29718));
  NANDX1 G17503 (.A1(W13750), .A2(W23671), .ZN(W25627));
  NANDX1 G17504 (.A1(W2156), .A2(W805), .ZN(W31504));
  NANDX1 G17505 (.A1(W21246), .A2(W6673), .ZN(W25599));
  NANDX1 G17506 (.A1(W19474), .A2(W19739), .ZN(W25621));
  NANDX1 G17507 (.A1(W16213), .A2(W10920), .ZN(O5817));
  NANDX1 G17508 (.A1(W3382), .A2(W289), .ZN(O3472));
  NANDX1 G17509 (.A1(W14595), .A2(W1006), .ZN(W28684));
  NANDX1 G17510 (.A1(W6070), .A2(W24010), .ZN(W29721));
  NANDX1 G17511 (.A1(W3605), .A2(W17164), .ZN(W28682));
  NANDX1 G17512 (.A1(W19171), .A2(W22271), .ZN(O4580));
  NANDX1 G17513 (.A1(W8887), .A2(W7266), .ZN(W29722));
  NANDX1 G17514 (.A1(W3383), .A2(W15853), .ZN(W28659));
  NANDX1 G17515 (.A1(W10878), .A2(W13635), .ZN(O4576));
  NANDX1 G17516 (.A1(W11502), .A2(W10904), .ZN(W27176));
  NANDX1 G17517 (.A1(W28166), .A2(W20803), .ZN(W29733));
  NANDX1 G17518 (.A1(W27734), .A2(W22116), .ZN(W28662));
  NANDX1 G17519 (.A1(W1363), .A2(W16640), .ZN(W31526));
  NANDX1 G17520 (.A1(W14960), .A2(I1244), .ZN(O4574));
  NANDX1 G17521 (.A1(W3288), .A2(W25982), .ZN(W31528));
  NANDX1 G17522 (.A1(W14724), .A2(W17984), .ZN(O4573));
  NANDX1 G17523 (.A1(W20219), .A2(W19109), .ZN(O3898));
  NANDX1 G17524 (.A1(W24162), .A2(W5815), .ZN(W31525));
  NANDX1 G17525 (.A1(W2685), .A2(W9886), .ZN(O4572));
  NANDX1 G17526 (.A1(W20052), .A2(W27424), .ZN(W28219));
  NANDX1 G17527 (.A1(W14860), .A2(W24064), .ZN(O4012));
  NANDX1 G17528 (.A1(W11051), .A2(W2867), .ZN(W28656));
  NANDX1 G17529 (.A1(W5126), .A2(I1949), .ZN(O4570));
  NANDX1 G17530 (.A1(W20342), .A2(W16970), .ZN(W28221));
  NANDX1 G17531 (.A1(W19099), .A2(W20951), .ZN(O4011));
  NANDX1 G17532 (.A1(W7961), .A2(W24824), .ZN(W25575));
  NANDX1 G17533 (.A1(W28065), .A2(W21610), .ZN(W28674));
  NANDX1 G17534 (.A1(W21014), .A2(W13178), .ZN(W26868));
  NANDX1 G17535 (.A1(W9809), .A2(W6542), .ZN(W25595));
  NANDX1 G17536 (.A1(W16170), .A2(W15134), .ZN(O5160));
  NANDX1 G17537 (.A1(W1187), .A2(W9314), .ZN(W28675));
  NANDX1 G17538 (.A1(W14838), .A2(W18150), .ZN(W25587));
  NANDX1 G17539 (.A1(W15219), .A2(W16007), .ZN(W25586));
  NANDX1 G17540 (.A1(W3207), .A2(W11427), .ZN(W29730));
  NANDX1 G17541 (.A1(W26158), .A2(W5704), .ZN(W31520));
  NANDX1 G17542 (.A1(W15052), .A2(W16854), .ZN(O3912));
  NANDX1 G17543 (.A1(W2753), .A2(W14401), .ZN(O5823));
  NANDX1 G17544 (.A1(W13051), .A2(W21458), .ZN(W25584));
  NANDX1 G17545 (.A1(W7959), .A2(W25680), .ZN(W28673));
  NANDX1 G17546 (.A1(W17968), .A2(W20984), .ZN(O4404));
  NANDX1 G17547 (.A1(W7159), .A2(I688), .ZN(O3897));
  NANDX1 G17548 (.A1(W20965), .A2(W2192), .ZN(W28672));
  NANDX1 G17549 (.A1(W714), .A2(W26225), .ZN(W28668));
  NANDX1 G17550 (.A1(W19280), .A2(W10717), .ZN(W27177));
  NANDX1 G17551 (.A1(W20456), .A2(W18593), .ZN(O5041));
  NANDX1 G17552 (.A1(W4020), .A2(W17533), .ZN(W31661));
  NANDX1 G17553 (.A1(W27678), .A2(W7089), .ZN(O4421));
  NANDX1 G17554 (.A1(W14049), .A2(W18847), .ZN(W28266));
  NANDX1 G17555 (.A1(W3031), .A2(W29397), .ZN(O5125));
  NANDX1 G17556 (.A1(W14500), .A2(W8219), .ZN(O5884));
  NANDX1 G17557 (.A1(W18254), .A2(W23479), .ZN(O5040));
  NANDX1 G17558 (.A1(W2538), .A2(W12130), .ZN(W27127));
  NANDX1 G17559 (.A1(W21715), .A2(W11635), .ZN(O5885));
  NANDX1 G17560 (.A1(W21379), .A2(W1767), .ZN(W25507));
  NANDX1 G17561 (.A1(W21017), .A2(W18130), .ZN(W31659));
  NANDX1 G17562 (.A1(W7510), .A2(W22462), .ZN(W25505));
  NANDX1 G17563 (.A1(W1303), .A2(W27514), .ZN(O5042));
  NANDX1 G17564 (.A1(W25401), .A2(W20216), .ZN(W31668));
  NANDX1 G17565 (.A1(W10774), .A2(W8557), .ZN(O4547));
  NANDX1 G17566 (.A1(W21507), .A2(W3680), .ZN(W28579));
  NANDX1 G17567 (.A1(W11689), .A2(W25968), .ZN(W28267));
  NANDX1 G17568 (.A1(W22694), .A2(W9366), .ZN(W26931));
  NANDX1 G17569 (.A1(W5343), .A2(W10580), .ZN(O3438));
  NANDX1 G17570 (.A1(W22113), .A2(W15147), .ZN(W28587));
  NANDX1 G17571 (.A1(W2688), .A2(W6818), .ZN(W26921));
  NANDX1 G17572 (.A1(W10027), .A2(I225), .ZN(W28262));
  NANDX1 G17573 (.A1(W10142), .A2(W14692), .ZN(O3994));
  NANDX1 G17574 (.A1(W1897), .A2(W12255), .ZN(W31649));
  NANDX1 G17575 (.A1(W9651), .A2(W18583), .ZN(W27132));
  NANDX1 G17576 (.A1(W14090), .A2(W28517), .ZN(W31652));
  NANDX1 G17577 (.A1(W4269), .A2(W1253), .ZN(O3441));
  NANDX1 G17578 (.A1(W20403), .A2(W11933), .ZN(W28263));
  NANDX1 G17579 (.A1(W12401), .A2(W7818), .ZN(W28588));
  NANDX1 G17580 (.A1(I260), .A2(W14167), .ZN(O5888));
  NANDX1 G17581 (.A1(W24687), .A2(W15556), .ZN(W29783));
  NANDX1 G17582 (.A1(W6219), .A2(W6716), .ZN(W28586));
  NANDX1 G17583 (.A1(W16767), .A2(W27121), .ZN(O5877));
  NANDX1 G17584 (.A1(W1006), .A2(W11765), .ZN(W27130));
  NANDX1 G17585 (.A1(W4179), .A2(W12873), .ZN(W25510));
  NANDX1 G17586 (.A1(W13364), .A2(W6678), .ZN(O3924));
  NANDX1 G17587 (.A1(W15505), .A2(W19271), .ZN(W28264));
  NANDX1 G17588 (.A1(W23374), .A2(W7986), .ZN(W29958));
  NANDX1 G17589 (.A1(W26250), .A2(W24347), .ZN(W26941));
  NANDX1 G17590 (.A1(W7260), .A2(W3019), .ZN(O3436));
  NANDX1 G17591 (.A1(W23580), .A2(W6106), .ZN(O5046));
  NANDX1 G17592 (.A1(W10314), .A2(W28328), .ZN(O5121));
  NANDX1 G17593 (.A1(W4296), .A2(W10145), .ZN(O5047));
  NANDX1 G17594 (.A1(W3959), .A2(W13388), .ZN(O4425));
  NANDX1 G17595 (.A1(W11494), .A2(W29812), .ZN(W29945));
  NANDX1 G17596 (.A1(W23912), .A2(W9557), .ZN(O4538));
  NANDX1 G17597 (.A1(W23176), .A2(W29037), .ZN(O5896));
  NANDX1 G17598 (.A1(W26669), .A2(W11164), .ZN(W28275));
  NANDX1 G17599 (.A1(W18378), .A2(W10878), .ZN(O5123));
  NANDX1 G17600 (.A1(W16770), .A2(W4557), .ZN(O4427));
  NANDX1 G17601 (.A1(W16156), .A2(W22547), .ZN(W29796));
  NANDX1 G17602 (.A1(W22140), .A2(W25792), .ZN(O5048));
  NANDX1 G17603 (.A1(W17680), .A2(W4701), .ZN(O3435));
  NANDX1 G17604 (.A1(W25532), .A2(W3696), .ZN(W26945));
  NANDX1 G17605 (.A1(W26454), .A2(I1934), .ZN(O3937));
  NANDX1 G17606 (.A1(W16028), .A2(W7736), .ZN(O4537));
  NANDX1 G17607 (.A1(W16183), .A2(W4173), .ZN(W28547));
  NANDX1 G17608 (.A1(I1014), .A2(W19380), .ZN(W27124));
  NANDX1 G17609 (.A1(W9607), .A2(W9963), .ZN(W31673));
  NANDX1 G17610 (.A1(I1058), .A2(W25950), .ZN(W28576));
  NANDX1 G17611 (.A1(W995), .A2(W24576), .ZN(W31674));
  NANDX1 G17612 (.A1(W25738), .A2(W23492), .ZN(O3926));
  NANDX1 G17613 (.A1(W27968), .A2(I692), .ZN(O4546));
  NANDX1 G17614 (.A1(W24119), .A2(W5394), .ZN(O5890));
  NANDX1 G17615 (.A1(W27521), .A2(I231), .ZN(W28572));
  NANDX1 G17616 (.A1(W25375), .A2(W27684), .ZN(W28571));
  NANDX1 G17617 (.A1(W469), .A2(W11602), .ZN(W27135));
  NANDX1 G17618 (.A1(W6657), .A2(W16850), .ZN(W29954));
  NANDX1 G17619 (.A1(W11214), .A2(W18737), .ZN(W29953));
  NANDX1 G17620 (.A1(W6144), .A2(W22283), .ZN(O4541));
  NANDX1 G17621 (.A1(W6670), .A2(W19967), .ZN(W28560));
  NANDX1 G17622 (.A1(W1888), .A2(W19545), .ZN(W28559));
  NANDX1 G17623 (.A1(W10819), .A2(W19276), .ZN(O4540));
  NANDX1 G17624 (.A1(W3040), .A2(W20724), .ZN(W28271));
  NANDX1 G17625 (.A1(W5830), .A2(W1962), .ZN(W25498));
  NANDX1 G17626 (.A1(W8532), .A2(W23315), .ZN(W25532));
  NANDX1 G17627 (.A1(W25143), .A2(W5978), .ZN(W28605));
  NANDX1 G17628 (.A1(W31470), .A2(W656), .ZN(O5857));
  NANDX1 G17629 (.A1(W7748), .A2(W15896), .ZN(O3450));
  NANDX1 G17630 (.A1(W15986), .A2(W21042), .ZN(W29865));
  NANDX1 G17631 (.A1(W15290), .A2(W5397), .ZN(W26903));
  NANDX1 G17632 (.A1(W1542), .A2(W4726), .ZN(O5140));
  NANDX1 G17633 (.A1(W29891), .A2(W27251), .ZN(O5858));
  NANDX1 G17634 (.A1(W6957), .A2(W3528), .ZN(W28242));
  NANDX1 G17635 (.A1(W11448), .A2(W26769), .ZN(O4556));
  NANDX1 G17636 (.A1(W10692), .A2(W8828), .ZN(O4415));
  NANDX1 G17637 (.A1(W11348), .A2(W22265), .ZN(W29762));
  NANDX1 G17638 (.A1(W17075), .A2(W17565), .ZN(O3998));
  NANDX1 G17639 (.A1(W18040), .A2(W15305), .ZN(W28243));
  NANDX1 G17640 (.A1(I1373), .A2(W19481), .ZN(O3914));
  NANDX1 G17641 (.A1(I1671), .A2(W21148), .ZN(W25530));
  NANDX1 G17642 (.A1(W22463), .A2(W11512), .ZN(W29981));
  NANDX1 G17643 (.A1(W27329), .A2(W16215), .ZN(W31611));
  NANDX1 G17644 (.A1(W17761), .A2(W19776), .ZN(W27141));
  NANDX1 G17645 (.A1(W16913), .A2(W1053), .ZN(W28616));
  NANDX1 G17646 (.A1(I1928), .A2(W28510), .ZN(W28622));
  NANDX1 G17647 (.A1(W9583), .A2(W12157), .ZN(W27152));
  NANDX1 G17648 (.A1(W393), .A2(W26074), .ZN(O4560));
  NANDX1 G17649 (.A1(W19006), .A2(W6388), .ZN(W28620));
  NANDX1 G17650 (.A1(W21699), .A2(W15952), .ZN(O5144));
  NANDX1 G17651 (.A1(W14689), .A2(W17392), .ZN(W25541));
  NANDX1 G17652 (.A1(W25962), .A2(W4739), .ZN(W26901));
  NANDX1 G17653 (.A1(W3096), .A2(W24071), .ZN(W28617));
  NANDX1 G17654 (.A1(W8873), .A2(W10395), .ZN(O5854));
  NANDX1 G17655 (.A1(W2253), .A2(W5622), .ZN(O3915));
  NANDX1 G17656 (.A1(W14960), .A2(W23884), .ZN(O5855));
  NANDX1 G17657 (.A1(W26309), .A2(W6196), .ZN(W28614));
  NANDX1 G17658 (.A1(W21735), .A2(W577), .ZN(O5143));
  NANDX1 G17659 (.A1(W9043), .A2(W11183), .ZN(O5142));
  NANDX1 G17660 (.A1(W3963), .A2(W7702), .ZN(W25537));
  NANDX1 G17661 (.A1(W4231), .A2(W8388), .ZN(W25536));
  NANDX1 G17662 (.A1(W20138), .A2(W14345), .ZN(W27150));
  NANDX1 G17663 (.A1(W27963), .A2(W1648), .ZN(W29984));
  NANDX1 G17664 (.A1(W22921), .A2(W18733), .ZN(W29959));
  NANDX1 G17665 (.A1(W3040), .A2(W14534), .ZN(W31630));
  NANDX1 G17666 (.A1(W4661), .A2(W7161), .ZN(W26916));
  NANDX1 G17667 (.A1(W8405), .A2(W3759), .ZN(O5038));
  NANDX1 G17668 (.A1(W16191), .A2(W10539), .ZN(O4554));
  NANDX1 G17669 (.A1(W4087), .A2(W14332), .ZN(W25519));
  NANDX1 G17670 (.A1(W14049), .A2(W24066), .ZN(W29776));
  NANDX1 G17671 (.A1(W14748), .A2(W13760), .ZN(O5126));
  NANDX1 G17672 (.A1(W22127), .A2(W4227), .ZN(O5866));
  NANDX1 G17673 (.A1(W7993), .A2(W26796), .ZN(W31632));
  NANDX1 G17674 (.A1(W31525), .A2(W14340), .ZN(W31629));
  NANDX1 G17675 (.A1(W23916), .A2(W30747), .ZN(W31633));
  NANDX1 G17676 (.A1(W14781), .A2(W19022), .ZN(W25516));
  NANDX1 G17677 (.A1(W14979), .A2(W22287), .ZN(W25514));
  NANDX1 G17678 (.A1(W2846), .A2(W19413), .ZN(W27136));
  NANDX1 G17679 (.A1(W20939), .A2(W9189), .ZN(W25513));
  NANDX1 G17680 (.A1(W17671), .A2(W7547), .ZN(W31636));
  NANDX1 G17681 (.A1(W22706), .A2(W8530), .ZN(O3442));
  NANDX1 G17682 (.A1(W7926), .A2(W348), .ZN(O5868));
  NANDX1 G17683 (.A1(W26383), .A2(W22255), .ZN(W26913));
  NANDX1 G17684 (.A1(W28608), .A2(W23749), .ZN(W29765));
  NANDX1 G17685 (.A1(W16233), .A2(I48), .ZN(W28600));
  NANDX1 G17686 (.A1(W3633), .A2(W9089), .ZN(O5134));
  NANDX1 G17687 (.A1(W18534), .A2(I1523), .ZN(O5133));
  NANDX1 G17688 (.A1(W6171), .A2(W18254), .ZN(W31618));
  NANDX1 G17689 (.A1(W29428), .A2(W22044), .ZN(O5862));
  NANDX1 G17690 (.A1(W6097), .A2(W5), .ZN(W29769));
  NANDX1 G17691 (.A1(W10170), .A2(W15824), .ZN(O5036));
  NANDX1 G17692 (.A1(W6741), .A2(W6851), .ZN(W26844));
  NANDX1 G17693 (.A1(W18237), .A2(W19459), .ZN(W28598));
  NANDX1 G17694 (.A1(W22346), .A2(W5768), .ZN(W28258));
  NANDX1 G17695 (.A1(W7024), .A2(W13907), .ZN(W26914));
  NANDX1 G17696 (.A1(W3363), .A2(W22488), .ZN(W31627));
  NANDX1 G17697 (.A1(W19969), .A2(W1163), .ZN(W28260));
  NANDX1 G17698 (.A1(W4039), .A2(W23385), .ZN(O4555));
  NANDX1 G17699 (.A1(W3046), .A2(W17763), .ZN(W25524));
  NANDX1 G17700 (.A1(W16826), .A2(W14240), .ZN(W27137));
  NANDX1 G17701 (.A1(W12706), .A2(W923), .ZN(O4218));
  NANDX1 G17702 (.A1(I1224), .A2(W29586), .ZN(W30861));
  NANDX1 G17703 (.A1(W23307), .A2(W19789), .ZN(W27749));
  NANDX1 G17704 (.A1(W16036), .A2(W20216), .ZN(W26196));
  NANDX1 G17705 (.A1(W23206), .A2(W9674), .ZN(W30864));
  NANDX1 G17706 (.A1(W24289), .A2(W577), .ZN(O3674));
  NANDX1 G17707 (.A1(W27213), .A2(W11985), .ZN(W29428));
  NANDX1 G17708 (.A1(W11657), .A2(W1490), .ZN(W27750));
  NANDX1 G17709 (.A1(W16754), .A2(W2037), .ZN(W26194));
  NANDX1 G17710 (.A1(W3454), .A2(W10236), .ZN(W30445));
  NANDX1 G17711 (.A1(W675), .A2(W4504), .ZN(O3795));
  NANDX1 G17712 (.A1(W729), .A2(W2740), .ZN(W26197));
  NANDX1 G17713 (.A1(W8359), .A2(W14921), .ZN(W29432));
  NANDX1 G17714 (.A1(W26311), .A2(W21017), .ZN(O4890));
  NANDX1 G17715 (.A1(W9140), .A2(W5033), .ZN(O4219));
  NANDX1 G17716 (.A1(W9726), .A2(W592), .ZN(W26562));
  NANDX1 G17717 (.A1(W25474), .A2(W15605), .ZN(O4110));
  NANDX1 G17718 (.A1(W11873), .A2(W25359), .ZN(W27753));
  NANDX1 G17719 (.A1(W14392), .A2(W13368), .ZN(W30443));
  NANDX1 G17720 (.A1(W25118), .A2(W25042), .ZN(O3672));
  NANDX1 G17721 (.A1(W1539), .A2(W16918), .ZN(W30870));
  NANDX1 G17722 (.A1(I1384), .A2(W1829), .ZN(W27745));
  NANDX1 G17723 (.A1(W6840), .A2(W24160), .ZN(W27467));
  NANDX1 G17724 (.A1(W6267), .A2(W11237), .ZN(W27744));
  NANDX1 G17725 (.A1(W27323), .A2(W20725), .ZN(W29426));
  NANDX1 G17726 (.A1(W7417), .A2(I1342), .ZN(O5524));
  NANDX1 G17727 (.A1(W23279), .A2(W5796), .ZN(O3678));
  NANDX1 G17728 (.A1(W24705), .A2(W19259), .ZN(O5340));
  NANDX1 G17729 (.A1(W8469), .A2(W11113), .ZN(W26209));
  NANDX1 G17730 (.A1(W21150), .A2(W19453), .ZN(W30859));
  NANDX1 G17731 (.A1(W19099), .A2(W2560), .ZN(O3677));
  NANDX1 G17732 (.A1(W26848), .A2(W21911), .ZN(W29145));
  NANDX1 G17733 (.A1(W13576), .A2(W12528), .ZN(W30872));
  NANDX1 G17734 (.A1(W17060), .A2(W23407), .ZN(W26205));
  NANDX1 G17735 (.A1(W10677), .A2(I1102), .ZN(W26203));
  NANDX1 G17736 (.A1(W23936), .A2(W29663), .ZN(O5337));
  NANDX1 G17737 (.A1(I1751), .A2(W15986), .ZN(W26202));
  NANDX1 G17738 (.A1(W6178), .A2(W7620), .ZN(W27746));
  NANDX1 G17739 (.A1(W21672), .A2(W12482), .ZN(W29141));
  NANDX1 G17740 (.A1(W18387), .A2(W14300), .ZN(W27747));
  NANDX1 G17741 (.A1(W16383), .A2(W589), .ZN(W26201));
  NANDX1 G17742 (.A1(W9269), .A2(W21581), .ZN(O3675));
  NANDX1 G17743 (.A1(W9805), .A2(W27075), .ZN(W27766));
  NANDX1 G17744 (.A1(W27387), .A2(W17257), .ZN(O4758));
  NANDX1 G17745 (.A1(W27538), .A2(W6518), .ZN(W30435));
  NANDX1 G17746 (.A1(W2921), .A2(W6092), .ZN(O3667));
  NANDX1 G17747 (.A1(W27257), .A2(W17228), .ZN(W27764));
  NANDX1 G17748 (.A1(W11841), .A2(W10800), .ZN(W29125));
  NANDX1 G17749 (.A1(W13311), .A2(W11854), .ZN(O3664));
  NANDX1 G17750 (.A1(W27334), .A2(W20267), .ZN(W29441));
  NANDX1 G17751 (.A1(W29637), .A2(W9537), .ZN(W30433));
  NANDX1 G17752 (.A1(W25577), .A2(W16220), .ZN(W29442));
  NANDX1 G17753 (.A1(W5884), .A2(W10363), .ZN(O4106));
  NANDX1 G17754 (.A1(W26194), .A2(W7655), .ZN(W29440));
  NANDX1 G17755 (.A1(W13688), .A2(W18962), .ZN(W29123));
  NANDX1 G17756 (.A1(W16115), .A2(W6781), .ZN(O5539));
  NANDX1 G17757 (.A1(W25680), .A2(W22536), .ZN(W29122));
  NANDX1 G17758 (.A1(W4477), .A2(W18070), .ZN(W26174));
  NANDX1 G17759 (.A1(W28466), .A2(W573), .ZN(W29445));
  NANDX1 G17760 (.A1(W5846), .A2(W6609), .ZN(O4896));
  NANDX1 G17761 (.A1(W17265), .A2(W4943), .ZN(W26570));
  NANDX1 G17762 (.A1(W25773), .A2(W17464), .ZN(W26571));
  NANDX1 G17763 (.A1(W11397), .A2(W3847), .ZN(W27769));
  NANDX1 G17764 (.A1(W10125), .A2(W22996), .ZN(W26565));
  NANDX1 G17765 (.A1(W9687), .A2(W16331), .ZN(O5529));
  NANDX1 G17766 (.A1(W11622), .A2(W4586), .ZN(W30878));
  NANDX1 G17767 (.A1(W6626), .A2(I260), .ZN(O3671));
  NANDX1 G17768 (.A1(W10960), .A2(W14399), .ZN(O5532));
  NANDX1 G17769 (.A1(W24803), .A2(W28285), .ZN(W29132));
  NANDX1 G17770 (.A1(W539), .A2(W30260), .ZN(O5533));
  NANDX1 G17771 (.A1(W7596), .A2(W3493), .ZN(W30439));
  NANDX1 G17772 (.A1(W14090), .A2(I19), .ZN(O5534));
  NANDX1 G17773 (.A1(W1547), .A2(W20691), .ZN(W27756));
  NANDX1 G17774 (.A1(W496), .A2(W24468), .ZN(W29424));
  NANDX1 G17775 (.A1(W13131), .A2(I1507), .ZN(W27758));
  NANDX1 G17776 (.A1(W23938), .A2(W7865), .ZN(W27445));
  NANDX1 G17777 (.A1(W352), .A2(W17508), .ZN(W27759));
  NANDX1 G17778 (.A1(W5940), .A2(W19891), .ZN(O4893));
  NANDX1 G17779 (.A1(W20438), .A2(W10862), .ZN(O3669));
  NANDX1 G17780 (.A1(W6872), .A2(W5656), .ZN(O3796));
  NANDX1 G17781 (.A1(W15794), .A2(I1927), .ZN(W27444));
  NANDX1 G17782 (.A1(W11454), .A2(W22091), .ZN(W26567));
  NANDX1 G17783 (.A1(W3700), .A2(W2382), .ZN(W26185));
  NANDX1 G17784 (.A1(I457), .A2(W124), .ZN(O3689));
  NANDX1 G17785 (.A1(W3307), .A2(W17867), .ZN(O4773));
  NANDX1 G17786 (.A1(W8896), .A2(W1103), .ZN(W26248));
  NANDX1 G17787 (.A1(W27626), .A2(W2482), .ZN(O5507));
  NANDX1 G17788 (.A1(I1706), .A2(W11263), .ZN(O4209));
  NANDX1 G17789 (.A1(W3334), .A2(W21530), .ZN(W27722));
  NANDX1 G17790 (.A1(W17746), .A2(W3662), .ZN(O4876));
  NANDX1 G17791 (.A1(W14525), .A2(W7002), .ZN(O4212));
  NANDX1 G17792 (.A1(W19827), .A2(W2033), .ZN(O5351));
  NANDX1 G17793 (.A1(W8083), .A2(W15681), .ZN(W27725));
  NANDX1 G17794 (.A1(W11655), .A2(W13009), .ZN(O5349));
  NANDX1 G17795 (.A1(W22714), .A2(W931), .ZN(O4208));
  NANDX1 G17796 (.A1(W777), .A2(W7984), .ZN(W27726));
  NANDX1 G17797 (.A1(W19115), .A2(W28645), .ZN(W29164));
  NANDX1 G17798 (.A1(W21544), .A2(W8192), .ZN(O3688));
  NANDX1 G17799 (.A1(W16246), .A2(W11217), .ZN(O4881));
  NANDX1 G17800 (.A1(W1343), .A2(W17562), .ZN(O3791));
  NANDX1 G17801 (.A1(W22354), .A2(W1249), .ZN(W27728));
  NANDX1 G17802 (.A1(W22503), .A2(W8554), .ZN(O5510));
  NANDX1 G17803 (.A1(W1515), .A2(W1816), .ZN(W27730));
  NANDX1 G17804 (.A1(W14081), .A2(W17001), .ZN(W26235));
  NANDX1 G17805 (.A1(W12193), .A2(W13138), .ZN(O4119));
  NANDX1 G17806 (.A1(W25964), .A2(W9676), .ZN(W27702));
  NANDX1 G17807 (.A1(W7303), .A2(W7137), .ZN(W27493));
  NANDX1 G17808 (.A1(W20220), .A2(W26160), .ZN(W26529));
  NANDX1 G17809 (.A1(W1603), .A2(W3819), .ZN(O3785));
  NANDX1 G17810 (.A1(W2199), .A2(W22706), .ZN(O4120));
  NANDX1 G17811 (.A1(W30019), .A2(W12451), .ZN(O5505));
  NANDX1 G17812 (.A1(W6061), .A2(W25581), .ZN(W26532));
  NANDX1 G17813 (.A1(W21328), .A2(W195), .ZN(W30479));
  NANDX1 G17814 (.A1(W10938), .A2(W21122), .ZN(O4874));
  NANDX1 G17815 (.A1(W5261), .A2(W17691), .ZN(O5511));
  NANDX1 G17816 (.A1(W2641), .A2(W22398), .ZN(W26257));
  NANDX1 G17817 (.A1(W5844), .A2(W28389), .ZN(W30819));
  NANDX1 G17818 (.A1(W16953), .A2(W17470), .ZN(W27482));
  NANDX1 G17819 (.A1(W28950), .A2(W2908), .ZN(O4875));
  NANDX1 G17820 (.A1(W23171), .A2(W13239), .ZN(W26535));
  NANDX1 G17821 (.A1(W16606), .A2(W11686), .ZN(W30475));
  NANDX1 G17822 (.A1(W21080), .A2(W14599), .ZN(W29404));
  NANDX1 G17823 (.A1(W8791), .A2(W29778), .ZN(O5506));
  NANDX1 G17824 (.A1(W11006), .A2(W22059), .ZN(O3788));
  NANDX1 G17825 (.A1(W23873), .A2(I1255), .ZN(W26549));
  NANDX1 G17826 (.A1(W24317), .A2(W15981), .ZN(W29419));
  NANDX1 G17827 (.A1(W1016), .A2(W3271), .ZN(W26225));
  NANDX1 G17828 (.A1(W20223), .A2(W12761), .ZN(W26224));
  NANDX1 G17829 (.A1(W26576), .A2(W24985), .ZN(W27470));
  NANDX1 G17830 (.A1(W28107), .A2(W23574), .ZN(O4770));
  NANDX1 G17831 (.A1(W14334), .A2(W2214), .ZN(O4884));
  NANDX1 G17832 (.A1(W18272), .A2(W10201), .ZN(W30845));
  NANDX1 G17833 (.A1(W14426), .A2(W8972), .ZN(O5521));
  NANDX1 G17834 (.A1(W18821), .A2(W15047), .ZN(W26222));
  NANDX1 G17835 (.A1(I952), .A2(I370), .ZN(W30847));
  NANDX1 G17836 (.A1(I481), .A2(W1681), .ZN(O3685));
  NANDX1 G17837 (.A1(W24704), .A2(W9839), .ZN(W26550));
  NANDX1 G17838 (.A1(W27089), .A2(W2425), .ZN(O5342));
  NANDX1 G17839 (.A1(W21741), .A2(W30328), .ZN(O5522));
  NANDX1 G17840 (.A1(W17960), .A2(W4356), .ZN(O3683));
  NANDX1 G17841 (.A1(W26209), .A2(I973), .ZN(W29155));
  NANDX1 G17842 (.A1(W16706), .A2(W25105), .ZN(W26217));
  NANDX1 G17843 (.A1(W28041), .A2(W12438), .ZN(W30455));
  NANDX1 G17844 (.A1(W25321), .A2(W26507), .ZN(W30453));
  NANDX1 G17845 (.A1(W27186), .A2(W24338), .ZN(O4216));
  NANDX1 G17846 (.A1(W10918), .A2(W15499), .ZN(W29417));
  NANDX1 G17847 (.A1(W846), .A2(W18796), .ZN(O4213));
  NANDX1 G17848 (.A1(W28395), .A2(W17923), .ZN(W30830));
  NANDX1 G17849 (.A1(W13751), .A2(W8197), .ZN(W27734));
  NANDX1 G17850 (.A1(W24748), .A2(W26343), .ZN(W30464));
  NANDX1 G17851 (.A1(W3824), .A2(W28164), .ZN(W29163));
  NANDX1 G17852 (.A1(W3139), .A2(W4391), .ZN(W27735));
  NANDX1 G17853 (.A1(W15657), .A2(W16713), .ZN(O5512));
  NANDX1 G17854 (.A1(I114), .A2(W5893), .ZN(W26230));
  NANDX1 G17855 (.A1(W11008), .A2(W19077), .ZN(W29161));
  NANDX1 G17856 (.A1(W30025), .A2(W23443), .ZN(W30432));
  NANDX1 G17857 (.A1(W30090), .A2(W7727), .ZN(O5513));
  NANDX1 G17858 (.A1(I1914), .A2(I868), .ZN(W26229));
  NANDX1 G17859 (.A1(W10635), .A2(W21174), .ZN(W27736));
  NANDX1 G17860 (.A1(W1174), .A2(W27441), .ZN(O5514));
  NANDX1 G17861 (.A1(W5880), .A2(W7886), .ZN(W27473));
  NANDX1 G17862 (.A1(W11977), .A2(W23255), .ZN(W30835));
  NANDX1 G17863 (.A1(W7326), .A2(W26756), .ZN(O4883));
  NANDX1 G17864 (.A1(W4108), .A2(W15887), .ZN(O5345));
  NANDX1 G17865 (.A1(W6611), .A2(W12204), .ZN(O5344));
  NANDX1 G17866 (.A1(W9830), .A2(W24033), .ZN(O3637));
  NANDX1 G17867 (.A1(W28691), .A2(W11665), .ZN(O4741));
  NANDX1 G17868 (.A1(W27733), .A2(W20345), .ZN(O5573));
  NANDX1 G17869 (.A1(W18510), .A2(W20698), .ZN(W29473));
  NANDX1 G17870 (.A1(W18149), .A2(W16369), .ZN(O5574));
  NANDX1 G17871 (.A1(W5863), .A2(W9608), .ZN(O3640));
  NANDX1 G17872 (.A1(W9457), .A2(W9687), .ZN(O3639));
  NANDX1 G17873 (.A1(W20722), .A2(I1329), .ZN(O3638));
  NANDX1 G17874 (.A1(W6034), .A2(W23301), .ZN(W27814));
  NANDX1 G17875 (.A1(W30632), .A2(I237), .ZN(O5575));
  NANDX1 G17876 (.A1(W6802), .A2(W1100), .ZN(W27429));
  NANDX1 G17877 (.A1(W24199), .A2(I1106), .ZN(O4913));
  NANDX1 G17878 (.A1(W6576), .A2(W9772), .ZN(W29474));
  NANDX1 G17879 (.A1(W17585), .A2(W17618), .ZN(O4241));
  NANDX1 G17880 (.A1(W23853), .A2(W26973), .ZN(O4736));
  NANDX1 G17881 (.A1(W1980), .A2(W13374), .ZN(W27428));
  NANDX1 G17882 (.A1(W1358), .A2(W12659), .ZN(W27817));
  NANDX1 G17883 (.A1(W3296), .A2(W9226), .ZN(W27427));
  NANDX1 G17884 (.A1(W23099), .A2(W6649), .ZN(W27820));
  NANDX1 G17885 (.A1(W356), .A2(W11630), .ZN(O5577));
  NANDX1 G17886 (.A1(W11220), .A2(W1174), .ZN(W29084));
  NANDX1 G17887 (.A1(W23214), .A2(W29389), .ZN(W30397));
  NANDX1 G17888 (.A1(W27200), .A2(W11808), .ZN(O5318));
  NANDX1 G17889 (.A1(I753), .A2(W4467), .ZN(O4744));
  NANDX1 G17890 (.A1(W13944), .A2(W11357), .ZN(W26595));
  NANDX1 G17891 (.A1(W25778), .A2(W19248), .ZN(W26132));
  NANDX1 G17892 (.A1(W5256), .A2(W14114), .ZN(W29101));
  NANDX1 G17893 (.A1(W16399), .A2(W30710), .ZN(W30947));
  NANDX1 G17894 (.A1(W13163), .A2(W18453), .ZN(W27434));
  NANDX1 G17895 (.A1(W10883), .A2(W24900), .ZN(O4743));
  NANDX1 G17896 (.A1(W1792), .A2(W22042), .ZN(W29099));
  NANDX1 G17897 (.A1(W5074), .A2(W23156), .ZN(W27810));
  NANDX1 G17898 (.A1(W17099), .A2(W27399), .ZN(O4734));
  NANDX1 G17899 (.A1(W29594), .A2(W21471), .ZN(W30396));
  NANDX1 G17900 (.A1(W25407), .A2(W25392), .ZN(O5314));
  NANDX1 G17901 (.A1(W27601), .A2(W4264), .ZN(W29464));
  NANDX1 G17902 (.A1(W6768), .A2(W20346), .ZN(O4102));
  NANDX1 G17903 (.A1(W1905), .A2(W6182), .ZN(O5313));
  NANDX1 G17904 (.A1(W24470), .A2(W12251), .ZN(W29095));
  NANDX1 G17905 (.A1(W21638), .A2(W12461), .ZN(O5570));
  NANDX1 G17906 (.A1(W4496), .A2(W6457), .ZN(W30955));
  NANDX1 G17907 (.A1(W17168), .A2(W8808), .ZN(O5572));
  NANDX1 G17908 (.A1(W24916), .A2(I932), .ZN(W30376));
  NANDX1 G17909 (.A1(W22027), .A2(W10929), .ZN(O4727));
  NANDX1 G17910 (.A1(W18555), .A2(W10723), .ZN(W26600));
  NANDX1 G17911 (.A1(W17342), .A2(W1874), .ZN(W30974));
  NANDX1 G17912 (.A1(W18281), .A2(W23397), .ZN(W30975));
  NANDX1 G17913 (.A1(W30230), .A2(W29379), .ZN(O5582));
  NANDX1 G17914 (.A1(W21157), .A2(W22537), .ZN(O4099));
  NANDX1 G17915 (.A1(W21336), .A2(W25270), .ZN(W26602));
  NANDX1 G17916 (.A1(W9618), .A2(W4556), .ZN(W26604));
  NANDX1 G17917 (.A1(I7), .A2(W22204), .ZN(W29483));
  NANDX1 G17918 (.A1(W26015), .A2(W21916), .ZN(W30980));
  NANDX1 G17919 (.A1(W4013), .A2(I669), .ZN(W27421));
  NANDX1 G17920 (.A1(W1036), .A2(W5841), .ZN(W26605));
  NANDX1 G17921 (.A1(I1668), .A2(W22356), .ZN(O5591));
  NANDX1 G17922 (.A1(W26348), .A2(W5227), .ZN(W26606));
  NANDX1 G17923 (.A1(W26347), .A2(W24680), .ZN(O5592));
  NANDX1 G17924 (.A1(W11390), .A2(W20703), .ZN(W29066));
  NANDX1 G17925 (.A1(W18386), .A2(W26491), .ZN(W27418));
  NANDX1 G17926 (.A1(W26185), .A2(W27391), .ZN(O5303));
  NANDX1 G17927 (.A1(W19684), .A2(W7156), .ZN(W30370));
  NANDX1 G17928 (.A1(W22373), .A2(W29539), .ZN(W30993));
  NANDX1 G17929 (.A1(W24024), .A2(W20738), .ZN(O3636));
  NANDX1 G17930 (.A1(W28186), .A2(W18096), .ZN(O5307));
  NANDX1 G17931 (.A1(W27208), .A2(W25999), .ZN(O4916));
  NANDX1 G17932 (.A1(W21209), .A2(W964), .ZN(W27426));
  NANDX1 G17933 (.A1(W18399), .A2(W1526), .ZN(W27821));
  NANDX1 G17934 (.A1(W2298), .A2(W26889), .ZN(O4918));
  NANDX1 G17935 (.A1(W4433), .A2(W4248), .ZN(W26114));
  NANDX1 G17936 (.A1(W16263), .A2(W16582), .ZN(O5306));
  NANDX1 G17937 (.A1(W12059), .A2(W16642), .ZN(O3805));
  NANDX1 G17938 (.A1(I1319), .A2(W3442), .ZN(W29077));
  NANDX1 G17939 (.A1(W30115), .A2(W27397), .ZN(W30943));
  NANDX1 G17940 (.A1(W22726), .A2(W13504), .ZN(O4731));
  NANDX1 G17941 (.A1(I687), .A2(W5947), .ZN(O4730));
  NANDX1 G17942 (.A1(W6719), .A2(W12043), .ZN(W30970));
  NANDX1 G17943 (.A1(W12330), .A2(I1500), .ZN(W29074));
  NANDX1 G17944 (.A1(W1390), .A2(W25868), .ZN(O4729));
  NANDX1 G17945 (.A1(W5479), .A2(W30419), .ZN(O5581));
  NANDX1 G17946 (.A1(W8228), .A2(I1438), .ZN(W29482));
  NANDX1 G17947 (.A1(W6239), .A2(W10713), .ZN(W26108));
  NANDX1 G17948 (.A1(W17039), .A2(W19806), .ZN(W27823));
  NANDX1 G17949 (.A1(W20302), .A2(W30054), .ZN(W30917));
  NANDX1 G17950 (.A1(W17184), .A2(W12282), .ZN(W26577));
  NANDX1 G17951 (.A1(W7050), .A2(W13695), .ZN(O3658));
  NANDX1 G17952 (.A1(W24621), .A2(W9306), .ZN(W29117));
  NANDX1 G17953 (.A1(W8585), .A2(W25421), .ZN(O5547));
  NANDX1 G17954 (.A1(W18615), .A2(W26931), .ZN(O5548));
  NANDX1 G17955 (.A1(W13700), .A2(I644), .ZN(W27783));
  NANDX1 G17956 (.A1(W18332), .A2(W28938), .ZN(O4899));
  NANDX1 G17957 (.A1(W4300), .A2(W29603), .ZN(W30427));
  NANDX1 G17958 (.A1(W7436), .A2(W27895), .ZN(W29116));
  NANDX1 G17959 (.A1(W22880), .A2(W5593), .ZN(W26156));
  NANDX1 G17960 (.A1(W5668), .A2(W8193), .ZN(O4231));
  NANDX1 G17961 (.A1(W16888), .A2(W25183), .ZN(W26155));
  NANDX1 G17962 (.A1(W26461), .A2(W2454), .ZN(W27784));
  NANDX1 G17963 (.A1(W16114), .A2(W20368), .ZN(W27786));
  NANDX1 G17964 (.A1(W12176), .A2(W1511), .ZN(W30918));
  NANDX1 G17965 (.A1(W15051), .A2(W7381), .ZN(O3799));
  NANDX1 G17966 (.A1(W18872), .A2(W988), .ZN(W30425));
  NANDX1 G17967 (.A1(W21924), .A2(W22900), .ZN(W27787));
  NANDX1 G17968 (.A1(W6378), .A2(W3283), .ZN(O3800));
  NANDX1 G17969 (.A1(W9363), .A2(W16993), .ZN(W30919));
  NANDX1 G17970 (.A1(W23597), .A2(W21682), .ZN(O4226));
  NANDX1 G17971 (.A1(W8260), .A2(W23370), .ZN(O4757));
  NANDX1 G17972 (.A1(W15051), .A2(W2053), .ZN(W29447));
  NANDX1 G17973 (.A1(W10671), .A2(W6618), .ZN(W27770));
  NANDX1 G17974 (.A1(W20873), .A2(W11608), .ZN(W26572));
  NANDX1 G17975 (.A1(W13223), .A2(W17787), .ZN(O3797));
  NANDX1 G17976 (.A1(W18859), .A2(W2292), .ZN(W30431));
  NANDX1 G17977 (.A1(W18975), .A2(W1158), .ZN(W27775));
  NANDX1 G17978 (.A1(I1681), .A2(W20339), .ZN(O4898));
  NANDX1 G17979 (.A1(W14419), .A2(W16830), .ZN(W26170));
  NANDX1 G17980 (.A1(W26582), .A2(W1590), .ZN(W27788));
  NANDX1 G17981 (.A1(W3238), .A2(W14314), .ZN(O4228));
  NANDX1 G17982 (.A1(W22626), .A2(W19714), .ZN(O5330));
  NANDX1 G17983 (.A1(W8708), .A2(W7470), .ZN(O3661));
  NANDX1 G17984 (.A1(W13911), .A2(W30093), .ZN(O5543));
  NANDX1 G17985 (.A1(W6705), .A2(W23665), .ZN(W26168));
  NANDX1 G17986 (.A1(W6887), .A2(W5059), .ZN(O5544));
  NANDX1 G17987 (.A1(W21826), .A2(W29847), .ZN(O5329));
  NANDX1 G17988 (.A1(W15171), .A2(W13907), .ZN(W26165));
  NANDX1 G17989 (.A1(W15375), .A2(W9268), .ZN(W29118));
  NANDX1 G17990 (.A1(W15903), .A2(W20678), .ZN(W26136));
  NANDX1 G17991 (.A1(W19127), .A2(W14894), .ZN(W26141));
  NANDX1 G17992 (.A1(W4389), .A2(W7599), .ZN(O3646));
  NANDX1 G17993 (.A1(W4891), .A2(W2538), .ZN(W26138));
  NANDX1 G17994 (.A1(W15232), .A2(W23772), .ZN(O5559));
  NANDX1 G17995 (.A1(W6154), .A2(W11034), .ZN(W26590));
  NANDX1 G17996 (.A1(W25765), .A2(W30684), .ZN(O5561));
  NANDX1 G17997 (.A1(W15300), .A2(I1778), .ZN(O3803));
  NANDX1 G17998 (.A1(W22899), .A2(W18537), .ZN(W27437));
  NANDX1 G17999 (.A1(W19428), .A2(W10617), .ZN(W26137));
  NANDX1 G18000 (.A1(W28587), .A2(W6560), .ZN(O5562));
  NANDX1 G18001 (.A1(W16128), .A2(W13752), .ZN(O4901));
  NANDX1 G18002 (.A1(W781), .A2(W12684), .ZN(W30939));
  NANDX1 G18003 (.A1(W11731), .A2(W17986), .ZN(W27801));
  NANDX1 G18004 (.A1(W11814), .A2(W19758), .ZN(W30941));
  NANDX1 G18005 (.A1(W2789), .A2(W22799), .ZN(O4746));
  NANDX1 G18006 (.A1(W24797), .A2(W20252), .ZN(O5564));
  NANDX1 G18007 (.A1(W1592), .A2(W21203), .ZN(O4236));
  NANDX1 G18008 (.A1(W1176), .A2(W24268), .ZN(W26134));
  NANDX1 G18009 (.A1(W20433), .A2(W5179), .ZN(O4906));
  NANDX1 G18010 (.A1(W16194), .A2(W6545), .ZN(O3645));
  NANDX1 G18011 (.A1(W18487), .A2(W27077), .ZN(O5557));
  NANDX1 G18012 (.A1(W1317), .A2(W25831), .ZN(W30423));
  NANDX1 G18013 (.A1(I894), .A2(W19288), .ZN(W26582));
  NANDX1 G18014 (.A1(W14299), .A2(W15251), .ZN(O3652));
  NANDX1 G18015 (.A1(W22347), .A2(W10554), .ZN(O5554));
  NANDX1 G18016 (.A1(W8561), .A2(I892), .ZN(O5327));
  NANDX1 G18017 (.A1(W25198), .A2(W10188), .ZN(W30924));
  NANDX1 G18018 (.A1(W16407), .A2(W21987), .ZN(W30420));
  NANDX1 G18019 (.A1(W21009), .A2(W9184), .ZN(O4104));
  NANDX1 G18020 (.A1(W29381), .A2(W7503), .ZN(O5556));
  NANDX1 G18021 (.A1(W7380), .A2(W18177), .ZN(O5359));
  NANDX1 G18022 (.A1(W7390), .A2(W26034), .ZN(W26146));
  NANDX1 G18023 (.A1(I659), .A2(W27422), .ZN(O4900));
  NANDX1 G18024 (.A1(W2434), .A2(W14977), .ZN(O5558));
  NANDX1 G18025 (.A1(W26459), .A2(W23184), .ZN(O5326));
  NANDX1 G18026 (.A1(W12560), .A2(W23906), .ZN(W27798));
  NANDX1 G18027 (.A1(I1720), .A2(W19884), .ZN(O5325));
  NANDX1 G18028 (.A1(W18896), .A2(W10829), .ZN(O3801));
  NANDX1 G18029 (.A1(W30202), .A2(W506), .ZN(W30412));
  NANDX1 G18030 (.A1(W20584), .A2(W6626), .ZN(O3650));
  NANDX1 G18031 (.A1(W11829), .A2(W17650), .ZN(W30569));
  NANDX1 G18032 (.A1(W3055), .A2(W22793), .ZN(W29258));
  NANDX1 G18033 (.A1(W20294), .A2(W18446), .ZN(O5401));
  NANDX1 G18034 (.A1(W19548), .A2(I157), .ZN(W26371));
  NANDX1 G18035 (.A1(W8793), .A2(W1017), .ZN(O3762));
  NANDX1 G18036 (.A1(W4438), .A2(W8453), .ZN(W30670));
  NANDX1 G18037 (.A1(W602), .A2(W15176), .ZN(O5444));
  NANDX1 G18038 (.A1(W12423), .A2(W24220), .ZN(W30673));
  NANDX1 G18039 (.A1(W823), .A2(W21628), .ZN(O5445));
  NANDX1 G18040 (.A1(W25168), .A2(W8549), .ZN(O4807));
  NANDX1 G18041 (.A1(W21027), .A2(W16281), .ZN(O4854));
  NANDX1 G18042 (.A1(W5934), .A2(W147), .ZN(O5402));
  NANDX1 G18043 (.A1(W21087), .A2(W13783), .ZN(W26367));
  NANDX1 G18044 (.A1(W7200), .A2(W8870), .ZN(W26366));
  NANDX1 G18045 (.A1(W5383), .A2(W5850), .ZN(O4855));
  NANDX1 G18046 (.A1(W24850), .A2(W6060), .ZN(W27605));
  NANDX1 G18047 (.A1(W5178), .A2(W23896), .ZN(W29246));
  NANDX1 G18048 (.A1(W20228), .A2(W22238), .ZN(O4165));
  NANDX1 G18049 (.A1(W12977), .A2(W9215), .ZN(W30683));
  NANDX1 G18050 (.A1(W22778), .A2(W23750), .ZN(O3763));
  NANDX1 G18051 (.A1(W16893), .A2(W4228), .ZN(O3764));
  NANDX1 G18052 (.A1(W23694), .A2(W8185), .ZN(W30669));
  NANDX1 G18053 (.A1(W15152), .A2(W8643), .ZN(O3738));
  NANDX1 G18054 (.A1(W18062), .A2(W10308), .ZN(W29267));
  NANDX1 G18055 (.A1(W19387), .A2(W21750), .ZN(W30580));
  NANDX1 G18056 (.A1(W4702), .A2(W17164), .ZN(W26385));
  NANDX1 G18057 (.A1(W10392), .A2(W9024), .ZN(O4809));
  NANDX1 G18058 (.A1(W4536), .A2(W25755), .ZN(W29265));
  NANDX1 G18059 (.A1(W2585), .A2(W5181), .ZN(O4846));
  NANDX1 G18060 (.A1(W13847), .A2(W24890), .ZN(W27537));
  NANDX1 G18061 (.A1(W5128), .A2(W1369), .ZN(W30665));
  NANDX1 G18062 (.A1(W15789), .A2(W21972), .ZN(W26380));
  NANDX1 G18063 (.A1(W8297), .A2(W452), .ZN(W27529));
  NANDX1 G18064 (.A1(W21928), .A2(I428), .ZN(W29261));
  NANDX1 G18065 (.A1(W640), .A2(W6559), .ZN(W26377));
  NANDX1 G18066 (.A1(W5232), .A2(W9433), .ZN(O4162));
  NANDX1 G18067 (.A1(W26729), .A2(W9534), .ZN(W30578));
  NANDX1 G18068 (.A1(W23933), .A2(W20708), .ZN(W26376));
  NANDX1 G18069 (.A1(I134), .A2(W17601), .ZN(O4141));
  NANDX1 G18070 (.A1(W5557), .A2(W27983), .ZN(W29259));
  NANDX1 G18071 (.A1(W12924), .A2(W18252), .ZN(W26375));
  NANDX1 G18072 (.A1(W7171), .A2(I1260), .ZN(O3733));
  NANDX1 G18073 (.A1(W12035), .A2(W24225), .ZN(W27631));
  NANDX1 G18074 (.A1(I538), .A2(W3154), .ZN(O5395));
  NANDX1 G18075 (.A1(W7827), .A2(W4398), .ZN(W30707));
  NANDX1 G18076 (.A1(W22064), .A2(W89), .ZN(W27621));
  NANDX1 G18077 (.A1(W15662), .A2(W26087), .ZN(W30709));
  NANDX1 G18078 (.A1(W5616), .A2(W23123), .ZN(W29358));
  NANDX1 G18079 (.A1(W2334), .A2(W14232), .ZN(W27625));
  NANDX1 G18080 (.A1(W15810), .A2(I1748), .ZN(W29239));
  NANDX1 G18081 (.A1(W22390), .A2(W26999), .ZN(W30710));
  NANDX1 G18082 (.A1(W4613), .A2(W13533), .ZN(W27627));
  NANDX1 G18083 (.A1(W13748), .A2(W1392), .ZN(O3766));
  NANDX1 G18084 (.A1(W15616), .A2(W21662), .ZN(W27619));
  NANDX1 G18085 (.A1(W23394), .A2(W2032), .ZN(W30560));
  NANDX1 G18086 (.A1(W2560), .A2(W20732), .ZN(O3726));
  NANDX1 G18087 (.A1(W23600), .A2(W1229), .ZN(W30559));
  NANDX1 G18088 (.A1(W28306), .A2(W27726), .ZN(O5394));
  NANDX1 G18089 (.A1(I1957), .A2(W4311), .ZN(W29237));
  NANDX1 G18090 (.A1(W10795), .A2(W5371), .ZN(W26347));
  NANDX1 G18091 (.A1(W7768), .A2(W16543), .ZN(W29236));
  NANDX1 G18092 (.A1(W4278), .A2(W14699), .ZN(W30719));
  NANDX1 G18093 (.A1(W11339), .A2(W2592), .ZN(W26346));
  NANDX1 G18094 (.A1(W4745), .A2(W12407), .ZN(W29356));
  NANDX1 G18095 (.A1(W19580), .A2(W3103), .ZN(W26363));
  NANDX1 G18096 (.A1(W9546), .A2(W16474), .ZN(O3765));
  NANDX1 G18097 (.A1(W3139), .A2(W14536), .ZN(O3730));
  NANDX1 G18098 (.A1(W10873), .A2(W21238), .ZN(W29245));
  NANDX1 G18099 (.A1(W14331), .A2(W12783), .ZN(W30690));
  NANDX1 G18100 (.A1(W8757), .A2(W15274), .ZN(W30692));
  NANDX1 G18101 (.A1(W26605), .A2(W15374), .ZN(W29244));
  NANDX1 G18102 (.A1(W10180), .A2(W6807), .ZN(W27608));
  NANDX1 G18103 (.A1(W11304), .A2(W3464), .ZN(O5397));
  NANDX1 G18104 (.A1(W17278), .A2(W18178), .ZN(O3739));
  NANDX1 G18105 (.A1(W11491), .A2(W17821), .ZN(W30564));
  NANDX1 G18106 (.A1(W25740), .A2(W775), .ZN(W26469));
  NANDX1 G18107 (.A1(I622), .A2(W7649), .ZN(O3728));
  NANDX1 G18108 (.A1(W19864), .A2(W16995), .ZN(O4168));
  NANDX1 G18109 (.A1(W2947), .A2(W29152), .ZN(O5456));
  NANDX1 G18110 (.A1(W5673), .A2(W23827), .ZN(O3727));
  NANDX1 G18111 (.A1(W25427), .A2(W12763), .ZN(O5458));
  NANDX1 G18112 (.A1(W25774), .A2(W12259), .ZN(W29240));
  NANDX1 G18113 (.A1(W27164), .A2(W21001), .ZN(W27617));
  NANDX1 G18114 (.A1(W16076), .A2(W18747), .ZN(W27582));
  NANDX1 G18115 (.A1(W2049), .A2(W9079), .ZN(W29303));
  NANDX1 G18116 (.A1(W10690), .A2(W3126), .ZN(W30626));
  NANDX1 G18117 (.A1(W5139), .A2(W9402), .ZN(W26414));
  NANDX1 G18118 (.A1(W28145), .A2(W19048), .ZN(O4831));
  NANDX1 G18119 (.A1(W16836), .A2(W14784), .ZN(W26410));
  NANDX1 G18120 (.A1(W709), .A2(W27140), .ZN(W27554));
  NANDX1 G18121 (.A1(W22587), .A2(W5108), .ZN(O4832));
  NANDX1 G18122 (.A1(W16326), .A2(W6847), .ZN(W29321));
  NANDX1 G18123 (.A1(W9829), .A2(W8368), .ZN(W27553));
  NANDX1 G18124 (.A1(W3034), .A2(W19404), .ZN(W27581));
  NANDX1 G18125 (.A1(W2260), .A2(W14896), .ZN(W26415));
  NANDX1 G18126 (.A1(W16520), .A2(W7170), .ZN(O4835));
  NANDX1 G18127 (.A1(W13356), .A2(W22494), .ZN(W29326));
  NANDX1 G18128 (.A1(W5953), .A2(W8486), .ZN(W29296));
  NANDX1 G18129 (.A1(W16880), .A2(W25910), .ZN(O3757));
  NANDX1 G18130 (.A1(W1392), .A2(W20167), .ZN(W29294));
  NANDX1 G18131 (.A1(W8572), .A2(W13159), .ZN(W30594));
  NANDX1 G18132 (.A1(W12522), .A2(W24116), .ZN(W29328));
  NANDX1 G18133 (.A1(W21022), .A2(W15199), .ZN(W27586));
  NANDX1 G18134 (.A1(I519), .A2(W10807), .ZN(W27549));
  NANDX1 G18135 (.A1(W14729), .A2(W17889), .ZN(O3753));
  NANDX1 G18136 (.A1(W1675), .A2(W16959), .ZN(W26428));
  NANDX1 G18137 (.A1(W17091), .A2(W27803), .ZN(O5411));
  NANDX1 G18138 (.A1(W1117), .A2(W8646), .ZN(O4149));
  NANDX1 G18139 (.A1(I228), .A2(W13905), .ZN(W29311));
  NANDX1 G18140 (.A1(W22811), .A2(W12395), .ZN(O3750));
  NANDX1 G18141 (.A1(W1570), .A2(W21326), .ZN(O5410));
  NANDX1 G18142 (.A1(W10786), .A2(W10655), .ZN(W30612));
  NANDX1 G18143 (.A1(W18659), .A2(W20266), .ZN(W27565));
  NANDX1 G18144 (.A1(W20923), .A2(W12592), .ZN(O4829));
  NANDX1 G18145 (.A1(W10130), .A2(W25507), .ZN(W26406));
  NANDX1 G18146 (.A1(W13807), .A2(I725), .ZN(W29314));
  NANDX1 G18147 (.A1(W14588), .A2(W3370), .ZN(O3749));
  NANDX1 G18148 (.A1(W21251), .A2(W22100), .ZN(W27569));
  NANDX1 G18149 (.A1(W27234), .A2(W25517), .ZN(O4151));
  NANDX1 G18150 (.A1(W1071), .A2(W18996), .ZN(W30616));
  NANDX1 G18151 (.A1(W24465), .A2(W18039), .ZN(W26430));
  NANDX1 G18152 (.A1(W7053), .A2(W695), .ZN(W27575));
  NANDX1 G18153 (.A1(W24324), .A2(W25355), .ZN(W26420));
  NANDX1 G18154 (.A1(W22486), .A2(W12673), .ZN(W26416));
  NANDX1 G18155 (.A1(W3100), .A2(W5809), .ZN(W27544));
  NANDX1 G18156 (.A1(W16573), .A2(W10737), .ZN(W27592));
  NANDX1 G18157 (.A1(W15470), .A2(W25610), .ZN(O3745));
  NANDX1 G18158 (.A1(I34), .A2(W13164), .ZN(W30590));
  NANDX1 G18159 (.A1(W21023), .A2(W17438), .ZN(O5430));
  NANDX1 G18160 (.A1(W2376), .A2(W17533), .ZN(O5432));
  NANDX1 G18161 (.A1(W4914), .A2(W28749), .ZN(W29274));
  NANDX1 G18162 (.A1(W18281), .A2(W18652), .ZN(O4142));
  NANDX1 G18163 (.A1(W13006), .A2(W9561), .ZN(W30649));
  NANDX1 G18164 (.A1(W10954), .A2(W24574), .ZN(O5403));
  NANDX1 G18165 (.A1(W18918), .A2(W11759), .ZN(W30652));
  NANDX1 G18166 (.A1(W12724), .A2(W114), .ZN(W26449));
  NANDX1 G18167 (.A1(W24024), .A2(W1646), .ZN(W26453));
  NANDX1 G18168 (.A1(W9358), .A2(W23070), .ZN(O4160));
  NANDX1 G18169 (.A1(W20126), .A2(W8218), .ZN(W27598));
  NANDX1 G18170 (.A1(W17619), .A2(W30363), .ZN(W30659));
  NANDX1 G18171 (.A1(W7095), .A2(W264), .ZN(W26396));
  NANDX1 G18172 (.A1(W6864), .A2(W9402), .ZN(W27540));
  NANDX1 G18173 (.A1(W19530), .A2(W28193), .ZN(W29337));
  NANDX1 G18174 (.A1(W8281), .A2(W13289), .ZN(O3743));
  NANDX1 G18175 (.A1(W24412), .A2(W11311), .ZN(W27601));
  NANDX1 G18176 (.A1(W19413), .A2(W3456), .ZN(W27548));
  NANDX1 G18177 (.A1(W24469), .A2(W4133), .ZN(W30593));
  NANDX1 G18178 (.A1(I581), .A2(W14455), .ZN(W29287));
  NANDX1 G18179 (.A1(W15246), .A2(W7961), .ZN(W30636));
  NANDX1 G18180 (.A1(W7362), .A2(W5393), .ZN(W29286));
  NANDX1 G18181 (.A1(W795), .A2(W25657), .ZN(W30592));
  NANDX1 G18182 (.A1(W6103), .A2(W25733), .ZN(W26403));
  NANDX1 G18183 (.A1(W23974), .A2(W16739), .ZN(W29280));
  NANDX1 G18184 (.A1(W12127), .A2(W14470), .ZN(W26446));
  NANDX1 G18185 (.A1(W29753), .A2(W4836), .ZN(W30639));
  NANDX1 G18186 (.A1(W9683), .A2(W22598), .ZN(O5463));
  NANDX1 G18187 (.A1(W15226), .A2(W9454), .ZN(W29276));
  NANDX1 G18188 (.A1(W20026), .A2(W5880), .ZN(O5425));
  NANDX1 G18189 (.A1(W962), .A2(W23805), .ZN(W26447));
  NANDX1 G18190 (.A1(W17886), .A2(W23940), .ZN(W26402));
  NANDX1 G18191 (.A1(W8639), .A2(W7210), .ZN(W26401));
  NANDX1 G18192 (.A1(W9141), .A2(W26305), .ZN(W29335));
  NANDX1 G18193 (.A1(W20327), .A2(W14316), .ZN(W29275));
  NANDX1 G18194 (.A1(W1122), .A2(W4143), .ZN(O4158));
  NANDX1 G18195 (.A1(W14872), .A2(W14690), .ZN(O5428));
  NANDX1 G18196 (.A1(W3548), .A2(W26486), .ZN(O4784));
  NANDX1 G18197 (.A1(W24313), .A2(W18068), .ZN(W27681));
  NANDX1 G18198 (.A1(W3890), .A2(W29434), .ZN(O5484));
  NANDX1 G18199 (.A1(W20041), .A2(W21), .ZN(W27508));
  NANDX1 G18200 (.A1(W22158), .A2(I164), .ZN(O5373));
  NANDX1 G18201 (.A1(W11878), .A2(W14642), .ZN(O5486));
  NANDX1 G18202 (.A1(W9087), .A2(W3364), .ZN(W30516));
  NANDX1 G18203 (.A1(W12736), .A2(W13347), .ZN(W26509));
  NANDX1 G18204 (.A1(W23240), .A2(W3953), .ZN(W27685));
  NANDX1 G18205 (.A1(W12755), .A2(W10016), .ZN(W26510));
  NANDX1 G18206 (.A1(W25419), .A2(W24555), .ZN(O5370));
  NANDX1 G18207 (.A1(W15488), .A2(W6606), .ZN(O4866));
  NANDX1 G18208 (.A1(W3798), .A2(W8394), .ZN(O5369));
  NANDX1 G18209 (.A1(W28391), .A2(W29757), .ZN(W30509));
  NANDX1 G18210 (.A1(W26100), .A2(W21279), .ZN(O5367));
  NANDX1 G18211 (.A1(W354), .A2(W8204), .ZN(W30506));
  NANDX1 G18212 (.A1(W29660), .A2(W13388), .ZN(W30781));
  NANDX1 G18213 (.A1(W4730), .A2(W592), .ZN(W30505));
  NANDX1 G18214 (.A1(W12970), .A2(W12626), .ZN(W26511));
  NANDX1 G18215 (.A1(W27543), .A2(W19665), .ZN(O4782));
  NANDX1 G18216 (.A1(W20660), .A2(W22781), .ZN(O4126));
  NANDX1 G18217 (.A1(I390), .A2(W8736), .ZN(O3707));
  NANDX1 G18218 (.A1(W18950), .A2(W14418), .ZN(W26503));
  NANDX1 G18219 (.A1(W9932), .A2(W7692), .ZN(W27668));
  NANDX1 G18220 (.A1(W18134), .A2(W20334), .ZN(O4865));
  NANDX1 G18221 (.A1(W7884), .A2(W18994), .ZN(W27670));
  NANDX1 G18222 (.A1(W14807), .A2(W13308), .ZN(W29203));
  NANDX1 G18223 (.A1(W20967), .A2(W375), .ZN(O3708));
  NANDX1 G18224 (.A1(W15887), .A2(W23583), .ZN(W30769));
  NANDX1 G18225 (.A1(W17969), .A2(W1725), .ZN(O4187));
  NANDX1 G18226 (.A1(W10228), .A2(W9792), .ZN(W27674));
  NANDX1 G18227 (.A1(W5567), .A2(W29151), .ZN(W29389));
  NANDX1 G18228 (.A1(W5404), .A2(I1028), .ZN(W29378));
  NANDX1 G18229 (.A1(W7959), .A2(W16623), .ZN(W30526));
  NANDX1 G18230 (.A1(W13622), .A2(W2657), .ZN(O4131));
  NANDX1 G18231 (.A1(W1515), .A2(W9186), .ZN(W30522));
  NANDX1 G18232 (.A1(W9290), .A2(W21709), .ZN(W27676));
  NANDX1 G18233 (.A1(W2801), .A2(W21612), .ZN(W26294));
  NANDX1 G18234 (.A1(W15333), .A2(W11334), .ZN(W29201));
  NANDX1 G18235 (.A1(W16147), .A2(W22320), .ZN(O4130));
  NANDX1 G18236 (.A1(W18070), .A2(W9074), .ZN(W30773));
  NANDX1 G18237 (.A1(W25955), .A2(W23294), .ZN(O4201));
  NANDX1 G18238 (.A1(W7901), .A2(W23805), .ZN(O4779));
  NANDX1 G18239 (.A1(W3551), .A2(W23169), .ZN(W26522));
  NANDX1 G18240 (.A1(W9885), .A2(W12703), .ZN(W26273));
  NANDX1 G18241 (.A1(I541), .A2(W20375), .ZN(W26524));
  NANDX1 G18242 (.A1(W16817), .A2(W27569), .ZN(O4777));
  NANDX1 G18243 (.A1(W22799), .A2(W16229), .ZN(O5498));
  NANDX1 G18244 (.A1(W8404), .A2(W29406), .ZN(W30808));
  NANDX1 G18245 (.A1(W28905), .A2(W10320), .ZN(W30810));
  NANDX1 G18246 (.A1(W5050), .A2(W13227), .ZN(W26526));
  NANDX1 G18247 (.A1(W19076), .A2(W17543), .ZN(O4776));
  NANDX1 G18248 (.A1(W3506), .A2(W29036), .ZN(W30803));
  NANDX1 G18249 (.A1(W25201), .A2(W22989), .ZN(W30487));
  NANDX1 G18250 (.A1(W11946), .A2(W16894), .ZN(W29393));
  NANDX1 G18251 (.A1(W15907), .A2(W1003), .ZN(W29172));
  NANDX1 G18252 (.A1(W16644), .A2(W18671), .ZN(O5503));
  NANDX1 G18253 (.A1(W24471), .A2(W4512), .ZN(W26264));
  NANDX1 G18254 (.A1(W503), .A2(W25081), .ZN(W27701));
  NANDX1 G18255 (.A1(I1158), .A2(W6345), .ZN(O5504));
  NANDX1 G18256 (.A1(W15959), .A2(W26083), .ZN(W26263));
  NANDX1 G18257 (.A1(W5501), .A2(W3483), .ZN(O4123));
  NANDX1 G18258 (.A1(W23049), .A2(W21938), .ZN(W26520));
  NANDX1 G18259 (.A1(W16746), .A2(W26286), .ZN(O5365));
  NANDX1 G18260 (.A1(I213), .A2(W11557), .ZN(W30785));
  NANDX1 G18261 (.A1(W4484), .A2(W2229), .ZN(W26514));
  NANDX1 G18262 (.A1(W20694), .A2(W27524), .ZN(W30498));
  NANDX1 G18263 (.A1(W10736), .A2(W22043), .ZN(W30787));
  NANDX1 G18264 (.A1(W11745), .A2(W11313), .ZN(O3780));
  NANDX1 G18265 (.A1(W5135), .A2(W9648), .ZN(O5490));
  NANDX1 G18266 (.A1(W29800), .A2(W3049), .ZN(W30495));
  NANDX1 G18267 (.A1(W12589), .A2(W3692), .ZN(W30789));
  NANDX1 G18268 (.A1(W26158), .A2(W7835), .ZN(O4133));
  NANDX1 G18269 (.A1(W13969), .A2(W10892), .ZN(O3703));
  NANDX1 G18270 (.A1(W13843), .A2(W25217), .ZN(O3702));
  NANDX1 G18271 (.A1(W7758), .A2(W22174), .ZN(W30791));
  NANDX1 G18272 (.A1(W21726), .A2(W23147), .ZN(O5491));
  NANDX1 G18273 (.A1(W22307), .A2(W14994), .ZN(W29181));
  NANDX1 G18274 (.A1(W16075), .A2(W24625), .ZN(W30492));
  NANDX1 G18275 (.A1(W25970), .A2(W24540), .ZN(O3782));
  NANDX1 G18276 (.A1(W3203), .A2(W13185), .ZN(W30801));
  NANDX1 G18277 (.A1(W15624), .A2(W18826), .ZN(W29179));
  NANDX1 G18278 (.A1(W3539), .A2(W14713), .ZN(O4173));
  NANDX1 G18279 (.A1(W10321), .A2(W12877), .ZN(W27641));
  NANDX1 G18280 (.A1(W455), .A2(W16847), .ZN(W29363));
  NANDX1 G18281 (.A1(W17859), .A2(I1177), .ZN(O4137));
  NANDX1 G18282 (.A1(W19719), .A2(W8025), .ZN(O5467));
  NANDX1 G18283 (.A1(W16496), .A2(W11248), .ZN(W30733));
  NANDX1 G18284 (.A1(W16591), .A2(W20051), .ZN(W27642));
  NANDX1 G18285 (.A1(W28063), .A2(W28474), .ZN(O4859));
  NANDX1 G18286 (.A1(W15147), .A2(W3174), .ZN(O3773));
  NANDX1 G18287 (.A1(W5540), .A2(W3137), .ZN(O3718));
  NANDX1 G18288 (.A1(W17507), .A2(W15866), .ZN(O3774));
  NANDX1 G18289 (.A1(W589), .A2(W19100), .ZN(W26485));
  NANDX1 G18290 (.A1(W11805), .A2(W11280), .ZN(W30736));
  NANDX1 G18291 (.A1(W6092), .A2(I1232), .ZN(W26324));
  NANDX1 G18292 (.A1(W29525), .A2(W19148), .ZN(W30737));
  NANDX1 G18293 (.A1(W17223), .A2(W18160), .ZN(O3775));
  NANDX1 G18294 (.A1(W28780), .A2(W30530), .ZN(W30739));
  NANDX1 G18295 (.A1(W23193), .A2(W3968), .ZN(W30549));
  NANDX1 G18296 (.A1(W3035), .A2(W29482), .ZN(W30740));
  NANDX1 G18297 (.A1(W16190), .A2(W2073), .ZN(O4175));
  NANDX1 G18298 (.A1(W8035), .A2(W17386), .ZN(W26495));
  NANDX1 G18299 (.A1(W13524), .A2(W19021), .ZN(W27637));
  NANDX1 G18300 (.A1(W12556), .A2(W10361), .ZN(O3767));
  NANDX1 G18301 (.A1(W14653), .A2(W3326), .ZN(O4171));
  NANDX1 G18302 (.A1(W21717), .A2(W15513), .ZN(W27635));
  NANDX1 G18303 (.A1(W12605), .A2(W15310), .ZN(W27636));
  NANDX1 G18304 (.A1(W15216), .A2(W10297), .ZN(W26473));
  NANDX1 G18305 (.A1(W26366), .A2(W14899), .ZN(O4798));
  NANDX1 G18306 (.A1(W6541), .A2(W4467), .ZN(W29230));
  NANDX1 G18307 (.A1(W25940), .A2(W8046), .ZN(O3723));
  NANDX1 G18308 (.A1(W25597), .A2(W24241), .ZN(O5466));
  NANDX1 G18309 (.A1(W9595), .A2(W16791), .ZN(W29372));
  NANDX1 G18310 (.A1(W21451), .A2(W5986), .ZN(O3722));
  NANDX1 G18311 (.A1(W1295), .A2(W21218), .ZN(W29359));
  NANDX1 G18312 (.A1(W13255), .A2(W9448), .ZN(O4172));
  NANDX1 G18313 (.A1(W54), .A2(W7984), .ZN(W26483));
  NANDX1 G18314 (.A1(W12213), .A2(W4992), .ZN(W27640));
  NANDX1 G18315 (.A1(W19407), .A2(W26716), .ZN(O5391));
  NANDX1 G18316 (.A1(W3978), .A2(W25921), .ZN(O4793));
  NANDX1 G18317 (.A1(W17910), .A2(W20516), .ZN(W27523));
  NANDX1 G18318 (.A1(W9942), .A2(W23151), .ZN(W26328));
  NANDX1 G18319 (.A1(W21348), .A2(W11188), .ZN(O4180));
  NANDX1 G18320 (.A1(W30266), .A2(W24384), .ZN(O5477));
  NANDX1 G18321 (.A1(W12342), .A2(W3324), .ZN(O5382));
  NANDX1 G18322 (.A1(W23319), .A2(W7029), .ZN(W30534));
  NANDX1 G18323 (.A1(W26205), .A2(W17826), .ZN(W26498));
  NANDX1 G18324 (.A1(W2804), .A2(W8369), .ZN(W29208));
  NANDX1 G18325 (.A1(W6624), .A2(W13191), .ZN(W29207));
  NANDX1 G18326 (.A1(W17818), .A2(W26227), .ZN(W30533));
  NANDX1 G18327 (.A1(W1980), .A2(W4834), .ZN(W29375));
  NANDX1 G18328 (.A1(W16391), .A2(W26841), .ZN(O4179));
  NANDX1 G18329 (.A1(W22594), .A2(W6011), .ZN(W26501));
  NANDX1 G18330 (.A1(W11391), .A2(W20387), .ZN(W26302));
  NANDX1 G18331 (.A1(W13533), .A2(W843), .ZN(O4181));
  NANDX1 G18332 (.A1(W29394), .A2(W28314), .ZN(W30761));
  NANDX1 G18333 (.A1(W21522), .A2(W13635), .ZN(W27661));
  NANDX1 G18334 (.A1(W19033), .A2(W21940), .ZN(W26301));
  NANDX1 G18335 (.A1(W14190), .A2(W14598), .ZN(O4134));
  NANDX1 G18336 (.A1(W11060), .A2(W8078), .ZN(O4182));
  NANDX1 G18337 (.A1(W16265), .A2(W26695), .ZN(O5482));
  NANDX1 G18338 (.A1(W19650), .A2(W14443), .ZN(W27664));
  NANDX1 G18339 (.A1(W9102), .A2(W18301), .ZN(W30765));
  NANDX1 G18340 (.A1(W25447), .A2(W308), .ZN(W30544));
  NANDX1 G18341 (.A1(W1291), .A2(W25073), .ZN(O5470));
  NANDX1 G18342 (.A1(W7738), .A2(W17812), .ZN(W26317));
  NANDX1 G18343 (.A1(W21734), .A2(W4355), .ZN(W30743));
  NANDX1 G18344 (.A1(W8543), .A2(W18505), .ZN(O3712));
  NANDX1 G18345 (.A1(W13224), .A2(W5889), .ZN(W27647));
  NANDX1 G18346 (.A1(W955), .A2(W5385), .ZN(O3776));
  NANDX1 G18347 (.A1(W1905), .A2(W16738), .ZN(W26497));
  NANDX1 G18348 (.A1(W13941), .A2(W12114), .ZN(O4136));
  NANDX1 G18349 (.A1(W10596), .A2(W13409), .ZN(W29216));
  NANDX1 G18350 (.A1(W5549), .A2(W30042), .ZN(O5301));
  NANDX1 G18351 (.A1(W13040), .A2(W412), .ZN(W26309));
  NANDX1 G18352 (.A1(W15171), .A2(W2147), .ZN(O5474));
  NANDX1 G18353 (.A1(W19474), .A2(W3406), .ZN(W26305));
  NANDX1 G18354 (.A1(W1702), .A2(W12710), .ZN(W30540));
  NANDX1 G18355 (.A1(W22777), .A2(W605), .ZN(W26303));
  NANDX1 G18356 (.A1(I1340), .A2(W12527), .ZN(O4791));
  NANDX1 G18357 (.A1(W2358), .A2(W3193), .ZN(W27519));
  NANDX1 G18358 (.A1(W20241), .A2(W17382), .ZN(W29210));
  NANDX1 G18359 (.A1(W27118), .A2(W13126), .ZN(O4135));
  NANDX1 G18360 (.A1(W17973), .A2(W20603), .ZN(W31254));
  NANDX1 G18361 (.A1(W632), .A2(W22356), .ZN(W26729));
  NANDX1 G18362 (.A1(W3324), .A2(W6505), .ZN(O5239));
  NANDX1 G18363 (.A1(W15565), .A2(W2061), .ZN(W25874));
  NANDX1 G18364 (.A1(W25851), .A2(W4345), .ZN(W27316));
  NANDX1 G18365 (.A1(W16878), .A2(W4168), .ZN(O3559));
  NANDX1 G18366 (.A1(W4333), .A2(W6135), .ZN(W31252));
  NANDX1 G18367 (.A1(W29005), .A2(W10006), .ZN(O5236));
  NANDX1 G18368 (.A1(W3093), .A2(W18358), .ZN(W30216));
  NANDX1 G18369 (.A1(W6677), .A2(W11278), .ZN(W25871));
  NANDX1 G18370 (.A1(W320), .A2(W7155), .ZN(W28878));
  NANDX1 G18371 (.A1(W6585), .A2(W24017), .ZN(W31250));
  NANDX1 G18372 (.A1(W18326), .A2(W14213), .ZN(O4649));
  NANDX1 G18373 (.A1(I387), .A2(W16550), .ZN(O3850));
  NANDX1 G18374 (.A1(W5280), .A2(W15517), .ZN(O4647));
  NANDX1 G18375 (.A1(W6695), .A2(W1396), .ZN(O3557));
  NANDX1 G18376 (.A1(W8123), .A2(W4893), .ZN(W28015));
  NANDX1 G18377 (.A1(W5056), .A2(W12692), .ZN(W31258));
  NANDX1 G18378 (.A1(W10104), .A2(W26821), .ZN(W31259));
  NANDX1 G18379 (.A1(I910), .A2(W19839), .ZN(W26732));
  NANDX1 G18380 (.A1(W9845), .A2(W8355), .ZN(W30214));
  NANDX1 G18381 (.A1(W22678), .A2(W24479), .ZN(O5707));
  NANDX1 G18382 (.A1(W14896), .A2(W23320), .ZN(W25880));
  NANDX1 G18383 (.A1(W3511), .A2(W9262), .ZN(W30229));
  NANDX1 G18384 (.A1(W11181), .A2(W776), .ZN(W27325));
  NANDX1 G18385 (.A1(I323), .A2(W29393), .ZN(W29595));
  NANDX1 G18386 (.A1(W23324), .A2(W19188), .ZN(W31242));
  NANDX1 G18387 (.A1(W23597), .A2(W17367), .ZN(W26725));
  NANDX1 G18388 (.A1(W10065), .A2(W2260), .ZN(W27322));
  NANDX1 G18389 (.A1(W12070), .A2(W17561), .ZN(O3848));
  NANDX1 G18390 (.A1(W16745), .A2(W13013), .ZN(W30225));
  NANDX1 G18391 (.A1(W22913), .A2(W25067), .ZN(W28006));
  NANDX1 G18392 (.A1(W17253), .A2(W8717), .ZN(W29603));
  NANDX1 G18393 (.A1(W2151), .A2(W42), .ZN(O3849));
  NANDX1 G18394 (.A1(W27815), .A2(W18733), .ZN(W28007));
  NANDX1 G18395 (.A1(W12761), .A2(W25128), .ZN(O3562));
  NANDX1 G18396 (.A1(W6051), .A2(W6816), .ZN(O4311));
  NANDX1 G18397 (.A1(W25931), .A2(W10549), .ZN(W30222));
  NANDX1 G18398 (.A1(W8201), .A2(W17277), .ZN(W28010));
  NANDX1 G18399 (.A1(W4696), .A2(W3591), .ZN(W27320));
  NANDX1 G18400 (.A1(W16063), .A2(W7546), .ZN(W27318));
  NANDX1 G18401 (.A1(W1231), .A2(W25611), .ZN(W25876));
  NANDX1 G18402 (.A1(I1946), .A2(W27466), .ZN(O4972));
  NANDX1 G18403 (.A1(W12966), .A2(I248), .ZN(O4062));
  NANDX1 G18404 (.A1(W158), .A2(W28699), .ZN(O4641));
  NANDX1 G18405 (.A1(W23644), .A2(W21691), .ZN(O5713));
  NANDX1 G18406 (.A1(I52), .A2(W19706), .ZN(W30207));
  NANDX1 G18407 (.A1(W25932), .A2(W26980), .ZN(O4970));
  NANDX1 G18408 (.A1(I600), .A2(W22955), .ZN(W28860));
  NANDX1 G18409 (.A1(I170), .A2(W28153), .ZN(W28859));
  NANDX1 G18410 (.A1(W24592), .A2(W3350), .ZN(W25845));
  NANDX1 G18411 (.A1(W10050), .A2(W20758), .ZN(W28858));
  NANDX1 G18412 (.A1(W2065), .A2(W23042), .ZN(W27308));
  NANDX1 G18413 (.A1(W2587), .A2(W11261), .ZN(W26739));
  NANDX1 G18414 (.A1(W14567), .A2(W2968), .ZN(W31274));
  NANDX1 G18415 (.A1(W3149), .A2(W10756), .ZN(O4061));
  NANDX1 G18416 (.A1(W7955), .A2(W16268), .ZN(O4060));
  NANDX1 G18417 (.A1(W4704), .A2(W16926), .ZN(W28028));
  NANDX1 G18418 (.A1(W16129), .A2(W6393), .ZN(O4319));
  NANDX1 G18419 (.A1(W26980), .A2(W689), .ZN(W30202));
  NANDX1 G18420 (.A1(W15380), .A2(W5402), .ZN(O5716));
  NANDX1 G18421 (.A1(W1258), .A2(W15058), .ZN(W25840));
  NANDX1 G18422 (.A1(W25539), .A2(W5787), .ZN(W28855));
  NANDX1 G18423 (.A1(W4760), .A2(W22841), .ZN(W28865));
  NANDX1 G18424 (.A1(W20659), .A2(W27003), .ZN(O5710));
  NANDX1 G18425 (.A1(W10884), .A2(W11821), .ZN(O3851));
  NANDX1 G18426 (.A1(W20146), .A2(W22093), .ZN(W31263));
  NANDX1 G18427 (.A1(W9661), .A2(W22335), .ZN(W27314));
  NANDX1 G18428 (.A1(W23849), .A2(W22382), .ZN(O3555));
  NANDX1 G18429 (.A1(W26693), .A2(W19464), .ZN(O4645));
  NANDX1 G18430 (.A1(W8097), .A2(W2554), .ZN(W25862));
  NANDX1 G18431 (.A1(I92), .A2(W10648), .ZN(W28023));
  NANDX1 G18432 (.A1(W1187), .A2(W24357), .ZN(O4644));
  NANDX1 G18433 (.A1(W4033), .A2(W7665), .ZN(O5706));
  NANDX1 G18434 (.A1(W8696), .A2(W20880), .ZN(O4643));
  NANDX1 G18435 (.A1(W10386), .A2(W22889), .ZN(W25852));
  NANDX1 G18436 (.A1(W12457), .A2(W11182), .ZN(O4967));
  NANDX1 G18437 (.A1(W27788), .A2(W22538), .ZN(O4642));
  NANDX1 G18438 (.A1(W10779), .A2(W10089), .ZN(O5232));
  NANDX1 G18439 (.A1(W3182), .A2(W11806), .ZN(W31269));
  NANDX1 G18440 (.A1(W24165), .A2(W9856), .ZN(W28024));
  NANDX1 G18441 (.A1(W26055), .A2(W3910), .ZN(O4317));
  NANDX1 G18442 (.A1(W4093), .A2(W13499), .ZN(W25848));
  NANDX1 G18443 (.A1(W12857), .A2(W15903), .ZN(O3572));
  NANDX1 G18444 (.A1(W22870), .A2(W24582), .ZN(W30244));
  NANDX1 G18445 (.A1(W19498), .A2(W2189), .ZN(O5682));
  NANDX1 G18446 (.A1(W2049), .A2(W17871), .ZN(O5684));
  NANDX1 G18447 (.A1(W25849), .A2(W24755), .ZN(W31204));
  NANDX1 G18448 (.A1(W15118), .A2(W21044), .ZN(W29572));
  NANDX1 G18449 (.A1(W28567), .A2(W20999), .ZN(O5250));
  NANDX1 G18450 (.A1(W2203), .A2(W18354), .ZN(O4658));
  NANDX1 G18451 (.A1(W1500), .A2(W15577), .ZN(W31207));
  NANDX1 G18452 (.A1(I923), .A2(W14275), .ZN(W31208));
  NANDX1 G18453 (.A1(W17517), .A2(W20942), .ZN(W25909));
  NANDX1 G18454 (.A1(W16706), .A2(W15856), .ZN(W27972));
  NANDX1 G18455 (.A1(W5788), .A2(W15411), .ZN(W26707));
  NANDX1 G18456 (.A1(W10186), .A2(I207), .ZN(O4655));
  NANDX1 G18457 (.A1(W3401), .A2(W17350), .ZN(O3571));
  NANDX1 G18458 (.A1(W21802), .A2(W16280), .ZN(O4304));
  NANDX1 G18459 (.A1(W14194), .A2(W17789), .ZN(W26708));
  NANDX1 G18460 (.A1(W4134), .A2(W7070), .ZN(O3570));
  NANDX1 G18461 (.A1(W6983), .A2(W22733), .ZN(W25904));
  NANDX1 G18462 (.A1(W19850), .A2(W4233), .ZN(O5249));
  NANDX1 G18463 (.A1(W11509), .A2(W24194), .ZN(W27338));
  NANDX1 G18464 (.A1(W1585), .A2(W5911), .ZN(O3576));
  NANDX1 G18465 (.A1(W8774), .A2(W1937), .ZN(W30253));
  NANDX1 G18466 (.A1(W494), .A2(W21362), .ZN(W25926));
  NANDX1 G18467 (.A1(W24077), .A2(W16414), .ZN(O4955));
  NANDX1 G18468 (.A1(W17009), .A2(W2443), .ZN(O3578));
  NANDX1 G18469 (.A1(W1320), .A2(W4864), .ZN(O5254));
  NANDX1 G18470 (.A1(W18672), .A2(W2557), .ZN(W25917));
  NANDX1 G18471 (.A1(W10761), .A2(W10105), .ZN(O3838));
  NANDX1 G18472 (.A1(W7118), .A2(W22328), .ZN(O4073));
  NANDX1 G18473 (.A1(W6917), .A2(W8245), .ZN(W27968));
  NANDX1 G18474 (.A1(W2169), .A2(W2083), .ZN(O4068));
  NANDX1 G18475 (.A1(W12615), .A2(W14245), .ZN(O4664));
  NANDX1 G18476 (.A1(W28748), .A2(W4034), .ZN(O4663));
  NANDX1 G18477 (.A1(W22294), .A2(W16138), .ZN(O3574));
  NANDX1 G18478 (.A1(W18699), .A2(W26027), .ZN(W28910));
  NANDX1 G18479 (.A1(I1182), .A2(W25306), .ZN(O3573));
  NANDX1 G18480 (.A1(W21516), .A2(W25885), .ZN(O4298));
  NANDX1 G18481 (.A1(W25056), .A2(W1908), .ZN(W28907));
  NANDX1 G18482 (.A1(W26665), .A2(W22517), .ZN(O4071));
  NANDX1 G18483 (.A1(I926), .A2(W4057), .ZN(W26701));
  NANDX1 G18484 (.A1(I541), .A2(W11561), .ZN(W31235));
  NANDX1 G18485 (.A1(W4436), .A2(W16775), .ZN(O3844));
  NANDX1 G18486 (.A1(W26020), .A2(W23173), .ZN(W31225));
  NANDX1 G18487 (.A1(W12499), .A2(W17549), .ZN(W28887));
  NANDX1 G18488 (.A1(W9562), .A2(W9188), .ZN(W26719));
  NANDX1 G18489 (.A1(W26862), .A2(W2958), .ZN(W28886));
  NANDX1 G18490 (.A1(W2727), .A2(W19622), .ZN(W28885));
  NANDX1 G18491 (.A1(W2569), .A2(W24282), .ZN(W26721));
  NANDX1 G18492 (.A1(I10), .A2(W13101), .ZN(W27999));
  NANDX1 G18493 (.A1(W4702), .A2(W27830), .ZN(W28883));
  NANDX1 G18494 (.A1(W1968), .A2(W5181), .ZN(O3563));
  NANDX1 G18495 (.A1(W21329), .A2(W16868), .ZN(O5699));
  NANDX1 G18496 (.A1(W15509), .A2(W4720), .ZN(W31237));
  NANDX1 G18497 (.A1(W22641), .A2(W23371), .ZN(O5244));
  NANDX1 G18498 (.A1(W9173), .A2(W5116), .ZN(W25882));
  NANDX1 G18499 (.A1(W17681), .A2(W378), .ZN(W28000));
  NANDX1 G18500 (.A1(W19538), .A2(W13757), .ZN(O5243));
  NANDX1 G18501 (.A1(W8041), .A2(W3553), .ZN(W26722));
  NANDX1 G18502 (.A1(W11755), .A2(W4133), .ZN(O5705));
  NANDX1 G18503 (.A1(W6220), .A2(W3262), .ZN(W28002));
  NANDX1 G18504 (.A1(W26604), .A2(W3806), .ZN(O4962));
  NANDX1 G18505 (.A1(W9152), .A2(W27016), .ZN(W27329));
  NANDX1 G18506 (.A1(W2868), .A2(I1091), .ZN(W29578));
  NANDX1 G18507 (.A1(W5872), .A2(W26761), .ZN(W29579));
  NANDX1 G18508 (.A1(W2308), .A2(W12251), .ZN(W28892));
  NANDX1 G18509 (.A1(W16046), .A2(W16160), .ZN(O4957));
  NANDX1 G18510 (.A1(I1176), .A2(W22895), .ZN(O3568));
  NANDX1 G18511 (.A1(W14312), .A2(W16619), .ZN(O4307));
  NANDX1 G18512 (.A1(W4323), .A2(W11582), .ZN(W31210));
  NANDX1 G18513 (.A1(W12086), .A2(W28750), .ZN(W29582));
  NANDX1 G18514 (.A1(W23309), .A2(W17467), .ZN(W26715));
  NANDX1 G18515 (.A1(W17242), .A2(W16102), .ZN(O4059));
  NANDX1 G18516 (.A1(W24713), .A2(W8301), .ZN(W27989));
  NANDX1 G18517 (.A1(W17139), .A2(W20751), .ZN(W31212));
  NANDX1 G18518 (.A1(W14109), .A2(W25011), .ZN(O4958));
  NANDX1 G18519 (.A1(W18612), .A2(W29639), .ZN(O5693));
  NANDX1 G18520 (.A1(W24120), .A2(W11462), .ZN(W28890));
  NANDX1 G18521 (.A1(W1746), .A2(W16238), .ZN(O4960));
  NANDX1 G18522 (.A1(I1594), .A2(W18420), .ZN(W31216));
  NANDX1 G18523 (.A1(W7930), .A2(W5111), .ZN(O4066));
  NANDX1 G18524 (.A1(W8468), .A2(W20200), .ZN(W29590));
  NANDX1 G18525 (.A1(W6762), .A2(W2487), .ZN(W26777));
  NANDX1 G18526 (.A1(W5990), .A2(W15937), .ZN(W31343));
  NANDX1 G18527 (.A1(W23136), .A2(W1877), .ZN(W26775));
  NANDX1 G18528 (.A1(W21654), .A2(W7179), .ZN(O3527));
  NANDX1 G18529 (.A1(W6345), .A2(W3112), .ZN(W31345));
  NANDX1 G18530 (.A1(W8835), .A2(W19210), .ZN(O5748));
  NANDX1 G18531 (.A1(W14447), .A2(W5419), .ZN(W25778));
  NANDX1 G18532 (.A1(W2674), .A2(W14808), .ZN(W30147));
  NANDX1 G18533 (.A1(W7322), .A2(W4520), .ZN(W31348));
  NANDX1 G18534 (.A1(W24951), .A2(W19563), .ZN(W25775));
  NANDX1 G18535 (.A1(W14862), .A2(W22419), .ZN(W30146));
  NANDX1 G18536 (.A1(W20420), .A2(W5354), .ZN(O3528));
  NANDX1 G18537 (.A1(W2073), .A2(W7689), .ZN(W30145));
  NANDX1 G18538 (.A1(W2925), .A2(W22326), .ZN(O3866));
  NANDX1 G18539 (.A1(W24709), .A2(W1697), .ZN(W31351));
  NANDX1 G18540 (.A1(W27745), .A2(W10098), .ZN(W31353));
  NANDX1 G18541 (.A1(W9398), .A2(W27611), .ZN(O5201));
  NANDX1 G18542 (.A1(W23606), .A2(W11027), .ZN(O3525));
  NANDX1 G18543 (.A1(W25478), .A2(W29042), .ZN(W30140));
  NANDX1 G18544 (.A1(W14376), .A2(W20752), .ZN(W31356));
  NANDX1 G18545 (.A1(W29608), .A2(W5867), .ZN(O5751));
  NANDX1 G18546 (.A1(W14967), .A2(W3137), .ZN(O4627));
  NANDX1 G18547 (.A1(W30773), .A2(W1067), .ZN(W31331));
  NANDX1 G18548 (.A1(W5261), .A2(W17130), .ZN(O5740));
  NANDX1 G18549 (.A1(W17851), .A2(W9137), .ZN(W30166));
  NANDX1 G18550 (.A1(I1076), .A2(W3668), .ZN(O4334));
  NANDX1 G18551 (.A1(W3138), .A2(W12527), .ZN(O3864));
  NANDX1 G18552 (.A1(W14687), .A2(W17582), .ZN(W25788));
  NANDX1 G18553 (.A1(W11160), .A2(W5781), .ZN(W29644));
  NANDX1 G18554 (.A1(W6032), .A2(W15693), .ZN(W25786));
  NANDX1 G18555 (.A1(W27251), .A2(W12531), .ZN(O4335));
  NANDX1 G18556 (.A1(W8739), .A2(W17030), .ZN(O4048));
  NANDX1 G18557 (.A1(W13526), .A2(W21668), .ZN(O5206));
  NANDX1 G18558 (.A1(W24893), .A2(W636), .ZN(O5743));
  NANDX1 G18559 (.A1(W15481), .A2(W5268), .ZN(O3530));
  NANDX1 G18560 (.A1(W13549), .A2(W26010), .ZN(O4337));
  NANDX1 G18561 (.A1(I1536), .A2(W10276), .ZN(O4050));
  NANDX1 G18562 (.A1(W14522), .A2(W16265), .ZN(W28810));
  NANDX1 G18563 (.A1(W16381), .A2(W12313), .ZN(O4988));
  NANDX1 G18564 (.A1(W1513), .A2(W18561), .ZN(W30149));
  NANDX1 G18565 (.A1(W27741), .A2(W22668), .ZN(O5745));
  NANDX1 G18566 (.A1(W21466), .A2(W20096), .ZN(O4992));
  NANDX1 G18567 (.A1(W8781), .A2(W5205), .ZN(W31369));
  NANDX1 G18568 (.A1(W25514), .A2(W19272), .ZN(O4990));
  NANDX1 G18569 (.A1(W18079), .A2(W11699), .ZN(W25767));
  NANDX1 G18570 (.A1(W8510), .A2(W9941), .ZN(O3523));
  NANDX1 G18571 (.A1(W12839), .A2(W20289), .ZN(O5200));
  NANDX1 G18572 (.A1(W23071), .A2(I1208), .ZN(W30135));
  NANDX1 G18573 (.A1(W24763), .A2(W24875), .ZN(W31371));
  NANDX1 G18574 (.A1(W4520), .A2(W13254), .ZN(W28794));
  NANDX1 G18575 (.A1(W17748), .A2(W13654), .ZN(W25763));
  NANDX1 G18576 (.A1(W24342), .A2(W11217), .ZN(O3521));
  NANDX1 G18577 (.A1(W12675), .A2(W21380), .ZN(O4620));
  NANDX1 G18578 (.A1(W24231), .A2(W3365), .ZN(O5756));
  NANDX1 G18579 (.A1(W22517), .A2(W16735), .ZN(O5757));
  NANDX1 G18580 (.A1(W20355), .A2(W24125), .ZN(W29654));
  NANDX1 G18581 (.A1(W13911), .A2(W15507), .ZN(W27264));
  NANDX1 G18582 (.A1(W4097), .A2(W1636), .ZN(W25751));
  NANDX1 G18583 (.A1(W11383), .A2(W13839), .ZN(O5759));
  NANDX1 G18584 (.A1(W27427), .A2(W18403), .ZN(W30131));
  NANDX1 G18585 (.A1(W3652), .A2(W6725), .ZN(O3872));
  NANDX1 G18586 (.A1(W15653), .A2(W23223), .ZN(W31379));
  NANDX1 G18587 (.A1(I1981), .A2(W20021), .ZN(W30137));
  NANDX1 G18588 (.A1(W16202), .A2(W21168), .ZN(W26781));
  NANDX1 G18589 (.A1(W15174), .A2(W3828), .ZN(O3867));
  NANDX1 G18590 (.A1(W5222), .A2(W23655), .ZN(O5752));
  NANDX1 G18591 (.A1(W20888), .A2(W23188), .ZN(O4622));
  NANDX1 G18592 (.A1(W4194), .A2(W16597), .ZN(O3869));
  NANDX1 G18593 (.A1(W12615), .A2(W31295), .ZN(W31362));
  NANDX1 G18594 (.A1(W8295), .A2(W19373), .ZN(W30138));
  NANDX1 G18595 (.A1(W21040), .A2(W26217), .ZN(O5755));
  NANDX1 G18596 (.A1(W20985), .A2(W11346), .ZN(W28077));
  NANDX1 G18597 (.A1(W29622), .A2(W6749), .ZN(W29642));
  NANDX1 G18598 (.A1(W22150), .A2(W14887), .ZN(O4339));
  NANDX1 G18599 (.A1(W25824), .A2(W14336), .ZN(W28081));
  NANDX1 G18600 (.A1(W6679), .A2(W7915), .ZN(O4989));
  NANDX1 G18601 (.A1(W22685), .A2(W9266), .ZN(O4341));
  NANDX1 G18602 (.A1(W6918), .A2(W7709), .ZN(W28084));
  NANDX1 G18603 (.A1(I766), .A2(W20174), .ZN(W25768));
  NANDX1 G18604 (.A1(W24732), .A2(W14797), .ZN(O4343));
  NANDX1 G18605 (.A1(W18332), .A2(I597), .ZN(W27271));
  NANDX1 G18606 (.A1(W10323), .A2(W4438), .ZN(O3870));
  NANDX1 G18607 (.A1(W6292), .A2(W19844), .ZN(O5221));
  NANDX1 G18608 (.A1(W17457), .A2(W6829), .ZN(O5721));
  NANDX1 G18609 (.A1(W4521), .A2(W16727), .ZN(W25823));
  NANDX1 G18610 (.A1(W9624), .A2(W9317), .ZN(W26752));
  NANDX1 G18611 (.A1(W680), .A2(W2741), .ZN(O5225));
  NANDX1 G18612 (.A1(W19291), .A2(W9680), .ZN(W25821));
  NANDX1 G18613 (.A1(W6799), .A2(W4166), .ZN(W25819));
  NANDX1 G18614 (.A1(W19284), .A2(W18096), .ZN(W28839));
  NANDX1 G18615 (.A1(W25558), .A2(W28938), .ZN(W30188));
  NANDX1 G18616 (.A1(W13208), .A2(W3551), .ZN(O5726));
  NANDX1 G18617 (.A1(W17039), .A2(W8368), .ZN(W30187));
  NANDX1 G18618 (.A1(W10452), .A2(W11325), .ZN(W29617));
  NANDX1 G18619 (.A1(W7230), .A2(W3080), .ZN(O4056));
  NANDX1 G18620 (.A1(W25697), .A2(W1608), .ZN(W26754));
  NANDX1 G18621 (.A1(W3370), .A2(W162), .ZN(W28836));
  NANDX1 G18622 (.A1(W26167), .A2(W8913), .ZN(W28835));
  NANDX1 G18623 (.A1(W20304), .A2(W3105), .ZN(W25811));
  NANDX1 G18624 (.A1(W18245), .A2(W30739), .ZN(O5727));
  NANDX1 G18625 (.A1(I759), .A2(W6322), .ZN(W26757));
  NANDX1 G18626 (.A1(W16988), .A2(W11092), .ZN(W28833));
  NANDX1 G18627 (.A1(W3202), .A2(W9868), .ZN(W25810));
  NANDX1 G18628 (.A1(W6948), .A2(W20070), .ZN(O4636));
  NANDX1 G18629 (.A1(W20042), .A2(W30178), .ZN(W30201));
  NANDX1 G18630 (.A1(W928), .A2(W16961), .ZN(O4321));
  NANDX1 G18631 (.A1(W8422), .A2(W21117), .ZN(O4638));
  NANDX1 G18632 (.A1(W20973), .A2(W2096), .ZN(W25836));
  NANDX1 G18633 (.A1(W20757), .A2(W490), .ZN(W28853));
  NANDX1 G18634 (.A1(I539), .A2(W10118), .ZN(O3857));
  NANDX1 G18635 (.A1(W11143), .A2(W21991), .ZN(W28851));
  NANDX1 G18636 (.A1(W25052), .A2(W28090), .ZN(O4637));
  NANDX1 G18637 (.A1(W19651), .A2(W20425), .ZN(O5718));
  NANDX1 G18638 (.A1(W4888), .A2(W7022), .ZN(O5729));
  NANDX1 G18639 (.A1(W19821), .A2(W20084), .ZN(O4322));
  NANDX1 G18640 (.A1(W22494), .A2(W25432), .ZN(O4974));
  NANDX1 G18641 (.A1(W12674), .A2(I596), .ZN(O4635));
  NANDX1 G18642 (.A1(W16949), .A2(I1686), .ZN(W25833));
  NANDX1 G18643 (.A1(W696), .A2(I255), .ZN(W30197));
  NANDX1 G18644 (.A1(W25848), .A2(W14315), .ZN(O4975));
  NANDX1 G18645 (.A1(W9815), .A2(W17392), .ZN(W30195));
  NANDX1 G18646 (.A1(I839), .A2(W9823), .ZN(W28842));
  NANDX1 G18647 (.A1(W6386), .A2(W4334), .ZN(W25827));
  NANDX1 G18648 (.A1(W1117), .A2(W19603), .ZN(W30174));
  NANDX1 G18649 (.A1(W2070), .A2(W23388), .ZN(W29633));
  NANDX1 G18650 (.A1(W17212), .A2(W6080), .ZN(O4983));
  NANDX1 G18651 (.A1(W20010), .A2(W15132), .ZN(O4629));
  NANDX1 G18652 (.A1(W10521), .A2(W17586), .ZN(W29637));
  NANDX1 G18653 (.A1(W9353), .A2(W14117), .ZN(O5736));
  NANDX1 G18654 (.A1(W21131), .A2(W8417), .ZN(W30176));
  NANDX1 G18655 (.A1(W22239), .A2(W27204), .ZN(W27287));
  NANDX1 G18656 (.A1(W7010), .A2(W1322), .ZN(W31324));
  NANDX1 G18657 (.A1(W26004), .A2(W24892), .ZN(W29639));
  NANDX1 G18658 (.A1(W27239), .A2(W6388), .ZN(O4328));
  NANDX1 G18659 (.A1(W12421), .A2(W13205), .ZN(O5215));
  NANDX1 G18660 (.A1(W20561), .A2(W2790), .ZN(O5737));
  NANDX1 G18661 (.A1(W17354), .A2(W19031), .ZN(W28061));
  NANDX1 G18662 (.A1(W12634), .A2(W14590), .ZN(W25797));
  NANDX1 G18663 (.A1(I118), .A2(W17597), .ZN(W30172));
  NANDX1 G18664 (.A1(W26556), .A2(W18715), .ZN(O5213));
  NANDX1 G18665 (.A1(W5793), .A2(I1104), .ZN(W28817));
  NANDX1 G18666 (.A1(W12410), .A2(W13419), .ZN(W31328));
  NANDX1 G18667 (.A1(W261), .A2(W5508), .ZN(W31330));
  NANDX1 G18668 (.A1(W5483), .A2(W13072), .ZN(W26769));
  NANDX1 G18669 (.A1(W928), .A2(W21833), .ZN(W29628));
  NANDX1 G18670 (.A1(W29709), .A2(W27497), .ZN(O5218));
  NANDX1 G18671 (.A1(W14075), .A2(W12645), .ZN(O4055));
  NANDX1 G18672 (.A1(W28713), .A2(W6055), .ZN(O4631));
  NANDX1 G18673 (.A1(W24485), .A2(I416), .ZN(W31308));
  NANDX1 G18674 (.A1(W10327), .A2(W26028), .ZN(O4979));
  NANDX1 G18675 (.A1(W7931), .A2(W24925), .ZN(W31310));
  NANDX1 G18676 (.A1(W14788), .A2(W16524), .ZN(W31311));
  NANDX1 G18677 (.A1(W14644), .A2(W21948), .ZN(O3536));
  NANDX1 G18678 (.A1(W11583), .A2(W2696), .ZN(W27293));
  NANDX1 G18679 (.A1(W219), .A2(W921), .ZN(O4297));
  NANDX1 G18680 (.A1(W30296), .A2(W12449), .ZN(W31312));
  NANDX1 G18681 (.A1(W24738), .A2(W27938), .ZN(W30180));
  NANDX1 G18682 (.A1(W29016), .A2(W9815), .ZN(O5216));
  NANDX1 G18683 (.A1(W4821), .A2(W4345), .ZN(W31316));
  NANDX1 G18684 (.A1(W22370), .A2(W9097), .ZN(W25803));
  NANDX1 G18685 (.A1(W4694), .A2(W14292), .ZN(W31317));
  NANDX1 G18686 (.A1(W18067), .A2(W14637), .ZN(W28824));
  NANDX1 G18687 (.A1(W8513), .A2(W8862), .ZN(W27292));
  NANDX1 G18688 (.A1(W27285), .A2(W6042), .ZN(W28051));
  NANDX1 G18689 (.A1(W925), .A2(W407), .ZN(O5286));
  NANDX1 G18690 (.A1(W25337), .A2(W16892), .ZN(O4704));
  NANDX1 G18691 (.A1(W457), .A2(W25114), .ZN(O5627));
  NANDX1 G18692 (.A1(W23380), .A2(W16221), .ZN(W29016));
  NANDX1 G18693 (.A1(W22092), .A2(W13958), .ZN(W31061));
  NANDX1 G18694 (.A1(W13975), .A2(W15621), .ZN(W27867));
  NANDX1 G18695 (.A1(W7973), .A2(W22449), .ZN(O3617));
  NANDX1 G18696 (.A1(W9430), .A2(W20747), .ZN(O4927));
  NANDX1 G18697 (.A1(W9546), .A2(W17461), .ZN(W30331));
  NANDX1 G18698 (.A1(I839), .A2(W4100), .ZN(W30330));
  NANDX1 G18699 (.A1(W26843), .A2(W27239), .ZN(W30327));
  NANDX1 G18700 (.A1(W3999), .A2(W17717), .ZN(W29511));
  NANDX1 G18701 (.A1(W24010), .A2(W50), .ZN(W29010));
  NANDX1 G18702 (.A1(W24622), .A2(W24096), .ZN(W30325));
  NANDX1 G18703 (.A1(W77), .A2(W18043), .ZN(O5285));
  NANDX1 G18704 (.A1(W2058), .A2(W16073), .ZN(O4698));
  NANDX1 G18705 (.A1(W10354), .A2(W91), .ZN(W30322));
  NANDX1 G18706 (.A1(W326), .A2(W4445), .ZN(W26054));
  NANDX1 G18707 (.A1(I1437), .A2(W3575), .ZN(O4928));
  NANDX1 G18708 (.A1(W16844), .A2(W2397), .ZN(O3814));
  NANDX1 G18709 (.A1(W11357), .A2(W14425), .ZN(O4261));
  NANDX1 G18710 (.A1(W17977), .A2(W13841), .ZN(W26634));
  NANDX1 G18711 (.A1(W12521), .A2(W15218), .ZN(O4712));
  NANDX1 G18712 (.A1(W10602), .A2(W4161), .ZN(W26072));
  NANDX1 G18713 (.A1(W9329), .A2(W9481), .ZN(W31051));
  NANDX1 G18714 (.A1(W13632), .A2(W920), .ZN(W26071));
  NANDX1 G18715 (.A1(W1091), .A2(W11366), .ZN(O5294));
  NANDX1 G18716 (.A1(W18226), .A2(W30174), .ZN(O5293));
  NANDX1 G18717 (.A1(W22039), .A2(W15831), .ZN(O3618));
  NANDX1 G18718 (.A1(W16259), .A2(W19004), .ZN(O4256));
  NANDX1 G18719 (.A1(W25003), .A2(W12699), .ZN(W26633));
  NANDX1 G18720 (.A1(W9894), .A2(W4078), .ZN(W31056));
  NANDX1 G18721 (.A1(W12608), .A2(W27538), .ZN(W31068));
  NANDX1 G18722 (.A1(W7939), .A2(W1783), .ZN(O4923));
  NANDX1 G18723 (.A1(W8189), .A2(W17589), .ZN(W30341));
  NANDX1 G18724 (.A1(W16929), .A2(W19308), .ZN(W29507));
  NANDX1 G18725 (.A1(W14434), .A2(W16489), .ZN(O4708));
  NANDX1 G18726 (.A1(W16929), .A2(W14085), .ZN(W30338));
  NANDX1 G18727 (.A1(W12433), .A2(I859), .ZN(W30336));
  NANDX1 G18728 (.A1(W27800), .A2(W1757), .ZN(O4706));
  NANDX1 G18729 (.A1(W1623), .A2(W2646), .ZN(O4926));
  NANDX1 G18730 (.A1(W6533), .A2(W17488), .ZN(O4260));
  NANDX1 G18731 (.A1(W25617), .A2(W6285), .ZN(W31084));
  NANDX1 G18732 (.A1(W25437), .A2(W25789), .ZN(W26644));
  NANDX1 G18733 (.A1(W12675), .A2(W534), .ZN(O3606));
  NANDX1 G18734 (.A1(W25731), .A2(W3415), .ZN(W26645));
  NANDX1 G18735 (.A1(W15961), .A2(W19123), .ZN(W26032));
  NANDX1 G18736 (.A1(W1020), .A2(W22148), .ZN(W30316));
  NANDX1 G18737 (.A1(W2298), .A2(I1988), .ZN(W28998));
  NANDX1 G18738 (.A1(W2159), .A2(W24930), .ZN(W28996));
  NANDX1 G18739 (.A1(W8015), .A2(W21648), .ZN(O4931));
  NANDX1 G18740 (.A1(W14308), .A2(W16374), .ZN(W26031));
  NANDX1 G18741 (.A1(W3046), .A2(W7568), .ZN(W26030));
  NANDX1 G18742 (.A1(W6870), .A2(W11541), .ZN(O4264));
  NANDX1 G18743 (.A1(W10196), .A2(W23351), .ZN(W27883));
  NANDX1 G18744 (.A1(W15014), .A2(W5631), .ZN(W26028));
  NANDX1 G18745 (.A1(W11736), .A2(I844), .ZN(W30308));
  NANDX1 G18746 (.A1(W17952), .A2(W13301), .ZN(W26025));
  NANDX1 G18747 (.A1(W13132), .A2(W5015), .ZN(W28993));
  NANDX1 G18748 (.A1(W11982), .A2(W6671), .ZN(W31088));
  NANDX1 G18749 (.A1(W25852), .A2(W14856), .ZN(O3604));
  NANDX1 G18750 (.A1(W14869), .A2(W28673), .ZN(W28991));
  NANDX1 G18751 (.A1(W10172), .A2(W15143), .ZN(W27387));
  NANDX1 G18752 (.A1(W4319), .A2(W17694), .ZN(O3816));
  NANDX1 G18753 (.A1(W23499), .A2(I1914), .ZN(O4697));
  NANDX1 G18754 (.A1(W15761), .A2(W24480), .ZN(O3614));
  NANDX1 G18755 (.A1(W3123), .A2(W18853), .ZN(O4089));
  NANDX1 G18756 (.A1(W20642), .A2(W23281), .ZN(O3815));
  NANDX1 G18757 (.A1(W3336), .A2(W16150), .ZN(O5630));
  NANDX1 G18758 (.A1(W21807), .A2(W7040), .ZN(O3612));
  NANDX1 G18759 (.A1(W22179), .A2(W9408), .ZN(O4929));
  NANDX1 G18760 (.A1(W6986), .A2(I353), .ZN(O3611));
  NANDX1 G18761 (.A1(W4448), .A2(W13265), .ZN(W31073));
  NANDX1 G18762 (.A1(W26755), .A2(W16471), .ZN(W27400));
  NANDX1 G18763 (.A1(W25436), .A2(W7510), .ZN(W26642));
  NANDX1 G18764 (.A1(W23902), .A2(W8190), .ZN(O3817));
  NANDX1 G18765 (.A1(W1309), .A2(W138), .ZN(W26043));
  NANDX1 G18766 (.A1(W18110), .A2(W11195), .ZN(W29003));
  NANDX1 G18767 (.A1(W11019), .A2(W25430), .ZN(O5633));
  NANDX1 G18768 (.A1(W6787), .A2(W13001), .ZN(O3608));
  NANDX1 G18769 (.A1(W6016), .A2(W5433), .ZN(W29002));
  NANDX1 G18770 (.A1(W25110), .A2(W4280), .ZN(W26035));
  NANDX1 G18771 (.A1(W3416), .A2(W12136), .ZN(O4262));
  NANDX1 G18772 (.A1(W15068), .A2(W2327), .ZN(O4249));
  NANDX1 G18773 (.A1(W3478), .A2(I1523), .ZN(O4247));
  NANDX1 G18774 (.A1(W11416), .A2(W22425), .ZN(W27840));
  NANDX1 G18775 (.A1(W19465), .A2(I1848), .ZN(O5601));
  NANDX1 G18776 (.A1(W19057), .A2(W11267), .ZN(W26614));
  NANDX1 G18777 (.A1(W27488), .A2(W6735), .ZN(W29057));
  NANDX1 G18778 (.A1(W5832), .A2(W10992), .ZN(W26616));
  NANDX1 G18779 (.A1(W27756), .A2(W13228), .ZN(O4248));
  NANDX1 G18780 (.A1(W29539), .A2(W12359), .ZN(W31007));
  NANDX1 G18781 (.A1(W28382), .A2(W15013), .ZN(W29054));
  NANDX1 G18782 (.A1(W15424), .A2(W17359), .ZN(W26100));
  NANDX1 G18783 (.A1(W262), .A2(W12974), .ZN(W30361));
  NANDX1 G18784 (.A1(W6292), .A2(W24892), .ZN(O3628));
  NANDX1 G18785 (.A1(W4377), .A2(W23537), .ZN(O3809));
  NANDX1 G18786 (.A1(W405), .A2(W24704), .ZN(O5602));
  NANDX1 G18787 (.A1(W13832), .A2(W18180), .ZN(O4722));
  NANDX1 G18788 (.A1(W19149), .A2(W8712), .ZN(O4919));
  NANDX1 G18789 (.A1(W10728), .A2(W26780), .ZN(W31009));
  NANDX1 G18790 (.A1(W10650), .A2(W19511), .ZN(W27414));
  NANDX1 G18791 (.A1(W23755), .A2(W13135), .ZN(O3626));
  NANDX1 G18792 (.A1(W27652), .A2(I1080), .ZN(O4718));
  NANDX1 G18793 (.A1(I1033), .A2(W4145), .ZN(W27829));
  NANDX1 G18794 (.A1(W25430), .A2(W26612), .ZN(O5299));
  NANDX1 G18795 (.A1(W11819), .A2(W22587), .ZN(W30365));
  NANDX1 G18796 (.A1(W11872), .A2(W15804), .ZN(W26607));
  NANDX1 G18797 (.A1(I1978), .A2(W3890), .ZN(W29064));
  NANDX1 G18798 (.A1(W8147), .A2(W123), .ZN(O3807));
  NANDX1 G18799 (.A1(W23959), .A2(W195), .ZN(O4725));
  NANDX1 G18800 (.A1(W8359), .A2(W18963), .ZN(W27828));
  NANDX1 G18801 (.A1(W10852), .A2(W18552), .ZN(W30996));
  NANDX1 G18802 (.A1(W3029), .A2(W13088), .ZN(W29061));
  NANDX1 G18803 (.A1(W13705), .A2(W24703), .ZN(W26088));
  NANDX1 G18804 (.A1(W21688), .A2(W26111), .ZN(O5596));
  NANDX1 G18805 (.A1(W8749), .A2(I1921), .ZN(O4724));
  NANDX1 G18806 (.A1(W18133), .A2(W26659), .ZN(O5597));
  NANDX1 G18807 (.A1(W2967), .A2(W7276), .ZN(O3633));
  NANDX1 G18808 (.A1(W6447), .A2(W17343), .ZN(O5298));
  NANDX1 G18809 (.A1(W16858), .A2(W7610), .ZN(O5598));
  NANDX1 G18810 (.A1(W24197), .A2(W23331), .ZN(W26612));
  NANDX1 G18811 (.A1(W28887), .A2(W22230), .ZN(W31004));
  NANDX1 G18812 (.A1(W12866), .A2(W15446), .ZN(W29059));
  NANDX1 G18813 (.A1(W16041), .A2(W14523), .ZN(W27404));
  NANDX1 G18814 (.A1(W15549), .A2(W655), .ZN(W31031));
  NANDX1 G18815 (.A1(W3728), .A2(W28251), .ZN(O5613));
  NANDX1 G18816 (.A1(W1799), .A2(W21083), .ZN(W27406));
  NANDX1 G18817 (.A1(W17383), .A2(W24317), .ZN(O5614));
  NANDX1 G18818 (.A1(W19480), .A2(W1503), .ZN(W29037));
  NANDX1 G18819 (.A1(I1666), .A2(W5215), .ZN(W29036));
  NANDX1 G18820 (.A1(W14041), .A2(W7145), .ZN(W31042));
  NANDX1 G18821 (.A1(W25342), .A2(W616), .ZN(W26079));
  NANDX1 G18822 (.A1(W5244), .A2(W29181), .ZN(W30348));
  NANDX1 G18823 (.A1(W22425), .A2(W5772), .ZN(O4715));
  NANDX1 G18824 (.A1(I1784), .A2(W13684), .ZN(O4922));
  NANDX1 G18825 (.A1(I1490), .A2(W3376), .ZN(W29498));
  NANDX1 G18826 (.A1(W16473), .A2(W11879), .ZN(W29032));
  NANDX1 G18827 (.A1(W684), .A2(W20739), .ZN(W27857));
  NANDX1 G18828 (.A1(W6520), .A2(W26624), .ZN(O5620));
  NANDX1 G18829 (.A1(W1183), .A2(W11369), .ZN(O3622));
  NANDX1 G18830 (.A1(W10320), .A2(W4847), .ZN(W26077));
  NANDX1 G18831 (.A1(W21913), .A2(W25948), .ZN(O5624));
  NANDX1 G18832 (.A1(W9632), .A2(W19488), .ZN(W27859));
  NANDX1 G18833 (.A1(W9204), .A2(W2046), .ZN(O4092));
  NANDX1 G18834 (.A1(W25947), .A2(W24225), .ZN(O4252));
  NANDX1 G18835 (.A1(W7212), .A2(W14973), .ZN(W26087));
  NANDX1 G18836 (.A1(W4794), .A2(W6552), .ZN(O3625));
  NANDX1 G18837 (.A1(W363), .A2(W26734), .ZN(O4921));
  NANDX1 G18838 (.A1(W22882), .A2(W21056), .ZN(W31014));
  NANDX1 G18839 (.A1(W21038), .A2(W2150), .ZN(W26621));
  NANDX1 G18840 (.A1(W29432), .A2(W28960), .ZN(W31016));
  NANDX1 G18841 (.A1(W22506), .A2(W15005), .ZN(O3812));
  NANDX1 G18842 (.A1(W19133), .A2(W7578), .ZN(W31021));
  NANDX1 G18843 (.A1(W26127), .A2(W15737), .ZN(W31022));
  NANDX1 G18844 (.A1(W13581), .A2(W22923), .ZN(O3603));
  NANDX1 G18845 (.A1(W25589), .A2(W1581), .ZN(O4094));
  NANDX1 G18846 (.A1(W18097), .A2(W21110), .ZN(W26082));
  NANDX1 G18847 (.A1(W6789), .A2(W4036), .ZN(O5609));
  NANDX1 G18848 (.A1(I1749), .A2(W4154), .ZN(O3623));
  NANDX1 G18849 (.A1(W9980), .A2(W17418), .ZN(O4253));
  NANDX1 G18850 (.A1(W29722), .A2(I1287), .ZN(O5611));
  NANDX1 G18851 (.A1(W13516), .A2(W6555), .ZN(W26626));
  NANDX1 G18852 (.A1(W6760), .A2(W14655), .ZN(W27854));
  NANDX1 G18853 (.A1(W10268), .A2(W10691), .ZN(O4254));
  NANDX1 G18854 (.A1(W19930), .A2(W2774), .ZN(O4950));
  NANDX1 G18855 (.A1(I146), .A2(W14027), .ZN(O4287));
  NANDX1 G18856 (.A1(W2231), .A2(W26047), .ZN(W28931));
  NANDX1 G18857 (.A1(I344), .A2(W12045), .ZN(W25957));
  NANDX1 G18858 (.A1(W20323), .A2(W13098), .ZN(W28929));
  NANDX1 G18859 (.A1(W7881), .A2(W27119), .ZN(W31163));
  NANDX1 G18860 (.A1(W18057), .A2(W1080), .ZN(W27357));
  NANDX1 G18861 (.A1(I1523), .A2(W7053), .ZN(W27356));
  NANDX1 G18862 (.A1(I1955), .A2(W7654), .ZN(O4289));
  NANDX1 G18863 (.A1(W21504), .A2(W30538), .ZN(O5670));
  NANDX1 G18864 (.A1(W11202), .A2(W17971), .ZN(W28928));
  NANDX1 G18865 (.A1(W29560), .A2(W11173), .ZN(O5667));
  NANDX1 G18866 (.A1(W7232), .A2(W26590), .ZN(O3831));
  NANDX1 G18867 (.A1(W26668), .A2(W16673), .ZN(W26679));
  NANDX1 G18868 (.A1(W20455), .A2(W15966), .ZN(W27943));
  NANDX1 G18869 (.A1(W7969), .A2(W18861), .ZN(W31167));
  NANDX1 G18870 (.A1(W22849), .A2(W17550), .ZN(W25953));
  NANDX1 G18871 (.A1(W24524), .A2(W18799), .ZN(W27947));
  NANDX1 G18872 (.A1(W20797), .A2(W13195), .ZN(W27949));
  NANDX1 G18873 (.A1(W2844), .A2(W13854), .ZN(O4292));
  NANDX1 G18874 (.A1(W24220), .A2(W25113), .ZN(W31170));
  NANDX1 G18875 (.A1(W4989), .A2(W13948), .ZN(W31154));
  NANDX1 G18876 (.A1(W9001), .A2(W11370), .ZN(W28952));
  NANDX1 G18877 (.A1(I562), .A2(W18595), .ZN(W28950));
  NANDX1 G18878 (.A1(W25671), .A2(W22857), .ZN(W26674));
  NANDX1 G18879 (.A1(W3496), .A2(I400), .ZN(W29546));
  NANDX1 G18880 (.A1(W19343), .A2(W20681), .ZN(W28947));
  NANDX1 G18881 (.A1(W15067), .A2(W23880), .ZN(W25967));
  NANDX1 G18882 (.A1(W21585), .A2(W4), .ZN(W28946));
  NANDX1 G18883 (.A1(W7467), .A2(W3715), .ZN(O4286));
  NANDX1 G18884 (.A1(W21434), .A2(W20749), .ZN(O5665));
  NANDX1 G18885 (.A1(I1038), .A2(W21616), .ZN(W27355));
  NANDX1 G18886 (.A1(W21713), .A2(W9397), .ZN(O3829));
  NANDX1 G18887 (.A1(I1835), .A2(W27821), .ZN(W28942));
  NANDX1 G18888 (.A1(W15936), .A2(W22325), .ZN(W27361));
  NANDX1 G18889 (.A1(W9230), .A2(I647), .ZN(W27360));
  NANDX1 G18890 (.A1(W11443), .A2(W4140), .ZN(W25962));
  NANDX1 G18891 (.A1(W22377), .A2(W28219), .ZN(W31157));
  NANDX1 G18892 (.A1(W23233), .A2(W20619), .ZN(W28941));
  NANDX1 G18893 (.A1(W22985), .A2(W17879), .ZN(W25958));
  NANDX1 G18894 (.A1(W1537), .A2(W26219), .ZN(W29552));
  NANDX1 G18895 (.A1(W18365), .A2(W28734), .ZN(W31184));
  NANDX1 G18896 (.A1(W18182), .A2(W23558), .ZN(O3835));
  NANDX1 G18897 (.A1(W18652), .A2(W13942), .ZN(W31182));
  NANDX1 G18898 (.A1(W11421), .A2(W4283), .ZN(W28923));
  NANDX1 G18899 (.A1(W23436), .A2(W7717), .ZN(O4075));
  NANDX1 G18900 (.A1(W22914), .A2(W4450), .ZN(W26690));
  NANDX1 G18901 (.A1(W16172), .A2(W10373), .ZN(W30260));
  NANDX1 G18902 (.A1(W9071), .A2(W19656), .ZN(W27960));
  NANDX1 G18903 (.A1(W2410), .A2(W14821), .ZN(W28919));
  NANDX1 G18904 (.A1(W5382), .A2(W8696), .ZN(W26694));
  NANDX1 G18905 (.A1(W26791), .A2(W15995), .ZN(O5674));
  NANDX1 G18906 (.A1(W17562), .A2(W15058), .ZN(W27350));
  NANDX1 G18907 (.A1(W23591), .A2(W6363), .ZN(W25935));
  NANDX1 G18908 (.A1(W10521), .A2(W13803), .ZN(W26695));
  NANDX1 G18909 (.A1(W23550), .A2(W19516), .ZN(O4296));
  NANDX1 G18910 (.A1(W4914), .A2(W10910), .ZN(W25933));
  NANDX1 G18911 (.A1(W11519), .A2(W9390), .ZN(W25931));
  NANDX1 G18912 (.A1(W20002), .A2(W19236), .ZN(W30258));
  NANDX1 G18913 (.A1(W13862), .A2(W6330), .ZN(O5677));
  NANDX1 G18914 (.A1(W25970), .A2(W26721), .ZN(W30255));
  NANDX1 G18915 (.A1(W1150), .A2(W16505), .ZN(W28915));
  NANDX1 G18916 (.A1(I1906), .A2(W6710), .ZN(W29559));
  NANDX1 G18917 (.A1(W974), .A2(W21921), .ZN(W31172));
  NANDX1 G18918 (.A1(W2463), .A2(W21144), .ZN(W31173));
  NANDX1 G18919 (.A1(W5684), .A2(W10686), .ZN(W25950));
  NANDX1 G18920 (.A1(W26712), .A2(W16576), .ZN(O5672));
  NANDX1 G18921 (.A1(W24183), .A2(W23657), .ZN(W30268));
  NANDX1 G18922 (.A1(W4216), .A2(W6796), .ZN(W30267));
  NANDX1 G18923 (.A1(W3779), .A2(W12352), .ZN(W25948));
  NANDX1 G18924 (.A1(W26409), .A2(W27380), .ZN(W27955));
  NANDX1 G18925 (.A1(W18424), .A2(W30722), .ZN(W31177));
  NANDX1 G18926 (.A1(W6723), .A2(W25572), .ZN(O3827));
  NANDX1 G18927 (.A1(W28818), .A2(W5507), .ZN(W31179));
  NANDX1 G18928 (.A1(W11085), .A2(W8219), .ZN(O4293));
  NANDX1 G18929 (.A1(W22354), .A2(W13393), .ZN(W29560));
  NANDX1 G18930 (.A1(W5402), .A2(W29961), .ZN(O5260));
  NANDX1 G18931 (.A1(I210), .A2(W686), .ZN(W27352));
  NANDX1 G18932 (.A1(W1516), .A2(W19275), .ZN(W31180));
  NANDX1 G18933 (.A1(W19735), .A2(W1704), .ZN(O4076));
  NANDX1 G18934 (.A1(W4617), .A2(W18659), .ZN(O3585));
  NANDX1 G18935 (.A1(W21729), .A2(W8814), .ZN(W28925));
  NANDX1 G18936 (.A1(W17708), .A2(W9225), .ZN(W28980));
  NANDX1 G18937 (.A1(W12154), .A2(W21487), .ZN(O4941));
  NANDX1 G18938 (.A1(W24226), .A2(W23541), .ZN(O3601));
  NANDX1 G18939 (.A1(W21998), .A2(W22214), .ZN(W27894));
  NANDX1 G18940 (.A1(W17746), .A2(W28707), .ZN(O4693));
  NANDX1 G18941 (.A1(I1902), .A2(W29757), .ZN(W31110));
  NANDX1 G18942 (.A1(W13894), .A2(W15731), .ZN(O4692));
  NANDX1 G18943 (.A1(W13025), .A2(W4421), .ZN(W27895));
  NANDX1 G18944 (.A1(W6922), .A2(I1715), .ZN(O4082));
  NANDX1 G18945 (.A1(W21697), .A2(W9834), .ZN(W27897));
  NANDX1 G18946 (.A1(W10531), .A2(W1204), .ZN(W31111));
  NANDX1 G18947 (.A1(W24422), .A2(W18564), .ZN(W26659));
  NANDX1 G18948 (.A1(W10973), .A2(W24719), .ZN(O4687));
  NANDX1 G18949 (.A1(W2477), .A2(W28665), .ZN(W28975));
  NANDX1 G18950 (.A1(W15921), .A2(W18905), .ZN(W26001));
  NANDX1 G18951 (.A1(W21823), .A2(W10319), .ZN(W25999));
  NANDX1 G18952 (.A1(W15763), .A2(W20839), .ZN(W26665));
  NANDX1 G18953 (.A1(W17052), .A2(W25353), .ZN(O4273));
  NANDX1 G18954 (.A1(I103), .A2(W9625), .ZN(O3598));
  NANDX1 G18955 (.A1(W24431), .A2(W10787), .ZN(W30294));
  NANDX1 G18956 (.A1(W3560), .A2(W8140), .ZN(W27906));
  NANDX1 G18957 (.A1(W19782), .A2(W12602), .ZN(O5643));
  NANDX1 G18958 (.A1(W12789), .A2(W8016), .ZN(O3821));
  NANDX1 G18959 (.A1(W5603), .A2(W4835), .ZN(O4936));
  NANDX1 G18960 (.A1(W3058), .A2(W24097), .ZN(W30303));
  NANDX1 G18961 (.A1(W5207), .A2(W20153), .ZN(O4695));
  NANDX1 G18962 (.A1(W1152), .A2(W19269), .ZN(W26016));
  NANDX1 G18963 (.A1(W1448), .A2(W9815), .ZN(W31096));
  NANDX1 G18964 (.A1(W3322), .A2(I636), .ZN(W26015));
  NANDX1 G18965 (.A1(W16791), .A2(W10998), .ZN(W31098));
  NANDX1 G18966 (.A1(W28106), .A2(W5417), .ZN(O4937));
  NANDX1 G18967 (.A1(W13781), .A2(W16626), .ZN(O3597));
  NANDX1 G18968 (.A1(W21246), .A2(W4213), .ZN(O5644));
  NANDX1 G18969 (.A1(W3285), .A2(W4592), .ZN(W26011));
  NANDX1 G18970 (.A1(I1674), .A2(W29218), .ZN(W31103));
  NANDX1 G18971 (.A1(W26458), .A2(I1904), .ZN(W31104));
  NANDX1 G18972 (.A1(W12526), .A2(W19197), .ZN(W27379));
  NANDX1 G18973 (.A1(W27581), .A2(W26122), .ZN(W30298));
  NANDX1 G18974 (.A1(W21895), .A2(W3320), .ZN(W26010));
  NANDX1 G18975 (.A1(W21752), .A2(W25917), .ZN(W27374));
  NANDX1 G18976 (.A1(W21476), .A2(W20225), .ZN(O4939));
  NANDX1 G18977 (.A1(W9214), .A2(W20550), .ZN(W25972));
  NANDX1 G18978 (.A1(W11045), .A2(W20228), .ZN(O4280));
  NANDX1 G18979 (.A1(W5587), .A2(W21353), .ZN(O4681));
  NANDX1 G18980 (.A1(W8325), .A2(W2643), .ZN(W25982));
  NANDX1 G18981 (.A1(W658), .A2(W8985), .ZN(W25979));
  NANDX1 G18982 (.A1(W11488), .A2(W1942), .ZN(O5653));
  NANDX1 G18983 (.A1(W11715), .A2(W27987), .ZN(W28958));
  NANDX1 G18984 (.A1(W9342), .A2(W1344), .ZN(W27929));
  NANDX1 G18985 (.A1(W8620), .A2(I414), .ZN(W25977));
  NANDX1 G18986 (.A1(W6756), .A2(W16126), .ZN(W29544));
  NANDX1 G18987 (.A1(W21449), .A2(W9769), .ZN(O3590));
  NANDX1 G18988 (.A1(W4112), .A2(W9242), .ZN(W26669));
  NANDX1 G18989 (.A1(W10830), .A2(W21071), .ZN(W28957));
  NANDX1 G18990 (.A1(I1407), .A2(W22300), .ZN(O4284));
  NANDX1 G18991 (.A1(W29708), .A2(W30425), .ZN(W31140));
  NANDX1 G18992 (.A1(W10782), .A2(W8670), .ZN(O4080));
  NANDX1 G18993 (.A1(W2700), .A2(W4799), .ZN(W31141));
  NANDX1 G18994 (.A1(W14515), .A2(W8265), .ZN(W27934));
  NANDX1 G18995 (.A1(W26752), .A2(I154), .ZN(W31142));
  NANDX1 G18996 (.A1(W3815), .A2(W21395), .ZN(O4679));
  NANDX1 G18997 (.A1(W13733), .A2(W11286), .ZN(W28954));
  NANDX1 G18998 (.A1(W13146), .A2(W19792), .ZN(O5266));
  NANDX1 G18999 (.A1(W7826), .A2(W1741), .ZN(O3596));
  NANDX1 G19000 (.A1(W8571), .A2(W10942), .ZN(W31118));
  NANDX1 G19001 (.A1(W1305), .A2(W15257), .ZN(O5648));
  NANDX1 G19002 (.A1(W181), .A2(W11901), .ZN(W25994));
  NANDX1 G19003 (.A1(W17351), .A2(W20975), .ZN(O3595));
  NANDX1 G19004 (.A1(W14774), .A2(W16256), .ZN(O5271));
  NANDX1 G19005 (.A1(I874), .A2(W1944), .ZN(O5649));
  NANDX1 G19006 (.A1(W13573), .A2(W24038), .ZN(O5270));
  NANDX1 G19007 (.A1(W19150), .A2(W19911), .ZN(O5267));
  NANDX1 G19008 (.A1(W12199), .A2(W3653), .ZN(W29655));
  NANDX1 G19009 (.A1(W333), .A2(W25598), .ZN(O4081));
  NANDX1 G19010 (.A1(W16210), .A2(W16946), .ZN(W27920));
  NANDX1 G19011 (.A1(W21593), .A2(W11801), .ZN(W30277));
  NANDX1 G19012 (.A1(W5070), .A2(I303), .ZN(W27921));
  NANDX1 G19013 (.A1(W2976), .A2(W14477), .ZN(W26666));
  NANDX1 G19014 (.A1(W6992), .A2(W13835), .ZN(O5651));
  NANDX1 G19015 (.A1(W5120), .A2(W3065), .ZN(W27923));
  NANDX1 G19016 (.A1(W25645), .A2(W5523), .ZN(O3592));
  NANDX1 G19017 (.A1(W7145), .A2(W6721), .ZN(O4683));
  NANDX1 G19018 (.A1(W38275), .A2(W42520), .ZN(O14032));
  NANDX1 G19019 (.A1(W22599), .A2(W36605), .ZN(O14075));
  NANDX1 G19020 (.A1(W34342), .A2(W17718), .ZN(O14069));
  NANDX1 G19021 (.A1(W10960), .A2(W10827), .ZN(O14060));
  NANDX1 G19022 (.A1(W36729), .A2(W43504), .ZN(W44619));
  NANDX1 G19023 (.A1(W8462), .A2(W11627), .ZN(O14051));
  NANDX1 G19024 (.A1(W34625), .A2(W43575), .ZN(O14048));
  NANDX1 G19025 (.A1(W40080), .A2(W9832), .ZN(O14045));
  NANDX1 G19026 (.A1(W4220), .A2(W2583), .ZN(O14041));
  NANDX1 G19027 (.A1(W1721), .A2(W23174), .ZN(O14039));
  NANDX1 G19028 (.A1(W18771), .A2(W27374), .ZN(O14038));
  NANDX1 G19029 (.A1(W17035), .A2(W4842), .ZN(O14037));
  NANDX1 G19030 (.A1(W12481), .A2(W10237), .ZN(O14036));
  NANDX1 G19031 (.A1(W12692), .A2(W34725), .ZN(O14077));
  NANDX1 G19032 (.A1(W8516), .A2(W36863), .ZN(W44594));
  NANDX1 G19033 (.A1(W35155), .A2(W39359), .ZN(O14029));
  NANDX1 G19034 (.A1(W36908), .A2(W9463), .ZN(O14028));
  NANDX1 G19035 (.A1(W16609), .A2(W9128), .ZN(O14027));
  NANDX1 G19036 (.A1(W28711), .A2(W39026), .ZN(O14022));
  NANDX1 G19037 (.A1(W8592), .A2(W16255), .ZN(O14021));
  NANDX1 G19038 (.A1(W9012), .A2(W6807), .ZN(O14019));
  NANDX1 G19039 (.A1(W36327), .A2(I664), .ZN(W44567));
  NANDX1 G19040 (.A1(W6793), .A2(W22632), .ZN(O14010));
  NANDX1 G19041 (.A1(W16988), .A2(W27021), .ZN(O14007));
  NANDX1 G19042 (.A1(W11686), .A2(W17996), .ZN(O14006));
  NANDX1 G19043 (.A1(W21579), .A2(W11931), .ZN(O14101));
  NANDX1 G19044 (.A1(W22082), .A2(W16021), .ZN(O14121));
  NANDX1 G19045 (.A1(W11778), .A2(W28033), .ZN(O14120));
  NANDX1 G19046 (.A1(W41241), .A2(W39002), .ZN(W44703));
  NANDX1 G19047 (.A1(W16488), .A2(W14719), .ZN(O14115));
  NANDX1 G19048 (.A1(W11158), .A2(W33880), .ZN(W44699));
  NANDX1 G19049 (.A1(W14130), .A2(W27118), .ZN(W44697));
  NANDX1 G19050 (.A1(W39275), .A2(W10270), .ZN(O14111));
  NANDX1 G19051 (.A1(W32850), .A2(W806), .ZN(W44689));
  NANDX1 G19052 (.A1(W20737), .A2(I1659), .ZN(O14107));
  NANDX1 G19053 (.A1(W13306), .A2(W32922), .ZN(O14105));
  NANDX1 G19054 (.A1(W13145), .A2(W13268), .ZN(O14104));
  NANDX1 G19055 (.A1(W23929), .A2(W2134), .ZN(O14102));
  NANDX1 G19056 (.A1(W15801), .A2(W9811), .ZN(O14004));
  NANDX1 G19057 (.A1(W32589), .A2(W20436), .ZN(O14100));
  NANDX1 G19058 (.A1(W9409), .A2(I245), .ZN(O14097));
  NANDX1 G19059 (.A1(W30978), .A2(W11579), .ZN(O14094));
  NANDX1 G19060 (.A1(W26008), .A2(W23184), .ZN(W44666));
  NANDX1 G19061 (.A1(W16098), .A2(W19017), .ZN(W44665));
  NANDX1 G19062 (.A1(W21230), .A2(W5243), .ZN(W44662));
  NANDX1 G19063 (.A1(W21314), .A2(W4404), .ZN(O14090));
  NANDX1 G19064 (.A1(W26227), .A2(W1913), .ZN(O14083));
  NANDX1 G19065 (.A1(W14741), .A2(W32889), .ZN(O14081));
  NANDX1 G19066 (.A1(W43440), .A2(W28753), .ZN(O14080));
  NANDX1 G19067 (.A1(W34829), .A2(W38980), .ZN(O14079));
  NANDX1 G19068 (.A1(W20552), .A2(W37872), .ZN(O13914));
  NANDX1 G19069 (.A1(W29458), .A2(W16966), .ZN(O13935));
  NANDX1 G19070 (.A1(W12845), .A2(W10966), .ZN(O13933));
  NANDX1 G19071 (.A1(W10078), .A2(W12478), .ZN(O13931));
  NANDX1 G19072 (.A1(W32641), .A2(W13547), .ZN(W44469));
  NANDX1 G19073 (.A1(W7589), .A2(W10286), .ZN(O13930));
  NANDX1 G19074 (.A1(W19414), .A2(W23644), .ZN(O13928));
  NANDX1 G19075 (.A1(W33299), .A2(W7673), .ZN(O13927));
  NANDX1 G19076 (.A1(W19100), .A2(W22585), .ZN(O13924));
  NANDX1 G19077 (.A1(W26282), .A2(W44289), .ZN(O13922));
  NANDX1 G19078 (.A1(W34784), .A2(W14402), .ZN(O13921));
  NANDX1 G19079 (.A1(W15382), .A2(W21534), .ZN(W44457));
  NANDX1 G19080 (.A1(W38183), .A2(W4459), .ZN(O13917));
  NANDX1 G19081 (.A1(W8074), .A2(W36945), .ZN(O13940));
  NANDX1 G19082 (.A1(W14781), .A2(W44348), .ZN(O13913));
  NANDX1 G19083 (.A1(W41210), .A2(W13230), .ZN(O13912));
  NANDX1 G19084 (.A1(W34168), .A2(W42150), .ZN(O13905));
  NANDX1 G19085 (.A1(W41900), .A2(W1144), .ZN(O13902));
  NANDX1 G19086 (.A1(W24511), .A2(W22861), .ZN(O13898));
  NANDX1 G19087 (.A1(W37395), .A2(W4059), .ZN(O13894));
  NANDX1 G19088 (.A1(W28832), .A2(W6155), .ZN(O13892));
  NANDX1 G19089 (.A1(W36953), .A2(W21714), .ZN(O13877));
  NANDX1 G19090 (.A1(W42633), .A2(W39432), .ZN(O13874));
  NANDX1 G19091 (.A1(W22513), .A2(W34150), .ZN(O13869));
  NANDX1 G19092 (.A1(W9449), .A2(W29241), .ZN(O13867));
  NANDX1 G19093 (.A1(W2281), .A2(W26992), .ZN(O13974));
  NANDX1 G19094 (.A1(W6608), .A2(W42431), .ZN(O14003));
  NANDX1 G19095 (.A1(W25684), .A2(W44246), .ZN(O14002));
  NANDX1 G19096 (.A1(W10722), .A2(W13713), .ZN(O13999));
  NANDX1 G19097 (.A1(I1953), .A2(W20473), .ZN(O13997));
  NANDX1 G19098 (.A1(W39807), .A2(W37475), .ZN(O13995));
  NANDX1 G19099 (.A1(W26628), .A2(W2034), .ZN(O13990));
  NANDX1 G19100 (.A1(W39502), .A2(W20506), .ZN(O13989));
  NANDX1 G19101 (.A1(W30619), .A2(W11253), .ZN(O13988));
  NANDX1 G19102 (.A1(W16161), .A2(W44015), .ZN(O13979));
  NANDX1 G19103 (.A1(W14868), .A2(W3474), .ZN(O13977));
  NANDX1 G19104 (.A1(W29739), .A2(W43504), .ZN(O13976));
  NANDX1 G19105 (.A1(W36596), .A2(W31739), .ZN(O14124));
  NANDX1 G19106 (.A1(W38032), .A2(W36329), .ZN(O13973));
  NANDX1 G19107 (.A1(W1899), .A2(W42175), .ZN(O13968));
  NANDX1 G19108 (.A1(W42972), .A2(W20824), .ZN(O13961));
  NANDX1 G19109 (.A1(W3331), .A2(W37222), .ZN(O13958));
  NANDX1 G19110 (.A1(I718), .A2(W12096), .ZN(O13957));
  NANDX1 G19111 (.A1(W38468), .A2(W37115), .ZN(W44501));
  NANDX1 G19112 (.A1(W9178), .A2(I75), .ZN(W44497));
  NANDX1 G19113 (.A1(W30272), .A2(W41866), .ZN(O13949));
  NANDX1 G19114 (.A1(W16798), .A2(W33644), .ZN(O13945));
  NANDX1 G19115 (.A1(W32214), .A2(W34674), .ZN(O13944));
  NANDX1 G19116 (.A1(W34604), .A2(W11167), .ZN(O13943));
  NANDX1 G19117 (.A1(W33931), .A2(I1020), .ZN(W44926));
  NANDX1 G19118 (.A1(W14033), .A2(W30024), .ZN(O14311));
  NANDX1 G19119 (.A1(W34486), .A2(W25949), .ZN(O14310));
  NANDX1 G19120 (.A1(W29380), .A2(W38032), .ZN(W44942));
  NANDX1 G19121 (.A1(W14431), .A2(W1046), .ZN(O14308));
  NANDX1 G19122 (.A1(W32630), .A2(W42717), .ZN(W44940));
  NANDX1 G19123 (.A1(W15271), .A2(W7287), .ZN(O14307));
  NANDX1 G19124 (.A1(W11657), .A2(W11196), .ZN(O14306));
  NANDX1 G19125 (.A1(W13542), .A2(W37112), .ZN(O14305));
  NANDX1 G19126 (.A1(W28693), .A2(W34099), .ZN(O14302));
  NANDX1 G19127 (.A1(W40718), .A2(W23650), .ZN(O14299));
  NANDX1 G19128 (.A1(W21118), .A2(W7776), .ZN(O14298));
  NANDX1 G19129 (.A1(W23873), .A2(W26365), .ZN(O14296));
  NANDX1 G19130 (.A1(W1571), .A2(W11778), .ZN(O14312));
  NANDX1 G19131 (.A1(W14080), .A2(W28373), .ZN(O14294));
  NANDX1 G19132 (.A1(W44755), .A2(W23764), .ZN(O14292));
  NANDX1 G19133 (.A1(W43691), .A2(W21769), .ZN(W44922));
  NANDX1 G19134 (.A1(W26315), .A2(W31555), .ZN(O14291));
  NANDX1 G19135 (.A1(W15379), .A2(W2688), .ZN(O14288));
  NANDX1 G19136 (.A1(W36849), .A2(W44655), .ZN(W44911));
  NANDX1 G19137 (.A1(W2736), .A2(W28051), .ZN(O14281));
  NANDX1 G19138 (.A1(W5329), .A2(W25537), .ZN(O14274));
  NANDX1 G19139 (.A1(W36488), .A2(W815), .ZN(O14273));
  NANDX1 G19140 (.A1(W4112), .A2(W42200), .ZN(O14270));
  NANDX1 G19141 (.A1(W44397), .A2(W26065), .ZN(O14268));
  NANDX1 G19142 (.A1(W32403), .A2(W160), .ZN(W44988));
  NANDX1 G19143 (.A1(W15208), .A2(W28855), .ZN(O14364));
  NANDX1 G19144 (.A1(I1051), .A2(W27465), .ZN(O14363));
  NANDX1 G19145 (.A1(W41488), .A2(W22171), .ZN(O14361));
  NANDX1 G19146 (.A1(W18586), .A2(W16911), .ZN(O14360));
  NANDX1 G19147 (.A1(W4435), .A2(W28074), .ZN(O14357));
  NANDX1 G19148 (.A1(W1428), .A2(I1326), .ZN(O14356));
  NANDX1 G19149 (.A1(W15461), .A2(W13544), .ZN(O14352));
  NANDX1 G19150 (.A1(W1970), .A2(W33287), .ZN(W44995));
  NANDX1 G19151 (.A1(W497), .A2(W34506), .ZN(O14351));
  NANDX1 G19152 (.A1(W27441), .A2(W44139), .ZN(O14350));
  NANDX1 G19153 (.A1(W15655), .A2(W35198), .ZN(W44990));
  NANDX1 G19154 (.A1(W38018), .A2(W33193), .ZN(W44989));
  NANDX1 G19155 (.A1(W17407), .A2(W5676), .ZN(W44884));
  NANDX1 G19156 (.A1(W15833), .A2(W27911), .ZN(O14345));
  NANDX1 G19157 (.A1(W1853), .A2(W37923), .ZN(O14337));
  NANDX1 G19158 (.A1(W10156), .A2(W10591), .ZN(O14333));
  NANDX1 G19159 (.A1(W251), .A2(W1861), .ZN(O14332));
  NANDX1 G19160 (.A1(W2424), .A2(W19473), .ZN(O14329));
  NANDX1 G19161 (.A1(I1259), .A2(W10596), .ZN(O14319));
  NANDX1 G19162 (.A1(W14786), .A2(W2670), .ZN(O14318));
  NANDX1 G19163 (.A1(W41939), .A2(W2520), .ZN(O14317));
  NANDX1 G19164 (.A1(W39323), .A2(W5745), .ZN(W44949));
  NANDX1 G19165 (.A1(W22371), .A2(W8826), .ZN(O14313));
  NANDX1 G19166 (.A1(W35384), .A2(W36704), .ZN(W44947));
  NANDX1 G19167 (.A1(W27761), .A2(W4936), .ZN(O14166));
  NANDX1 G19168 (.A1(I712), .A2(W38738), .ZN(O14203));
  NANDX1 G19169 (.A1(W31146), .A2(W23435), .ZN(O14199));
  NANDX1 G19170 (.A1(W42042), .A2(W43517), .ZN(O14194));
  NANDX1 G19171 (.A1(W44261), .A2(W51), .ZN(O14188));
  NANDX1 G19172 (.A1(W34135), .A2(W15977), .ZN(O14184));
  NANDX1 G19173 (.A1(W42670), .A2(W16917), .ZN(O14179));
  NANDX1 G19174 (.A1(I357), .A2(W37196), .ZN(O14178));
  NANDX1 G19175 (.A1(W5496), .A2(W43622), .ZN(O14177));
  NANDX1 G19176 (.A1(W11315), .A2(W24986), .ZN(W44774));
  NANDX1 G19177 (.A1(W2303), .A2(W2158), .ZN(O14172));
  NANDX1 G19178 (.A1(W33671), .A2(W40212), .ZN(O14169));
  NANDX1 G19179 (.A1(W28668), .A2(W38256), .ZN(W44766));
  NANDX1 G19180 (.A1(W26267), .A2(W3459), .ZN(W44814));
  NANDX1 G19181 (.A1(W23654), .A2(W42099), .ZN(W44760));
  NANDX1 G19182 (.A1(W8913), .A2(W673), .ZN(O14162));
  NANDX1 G19183 (.A1(W44697), .A2(W2840), .ZN(W44755));
  NANDX1 G19184 (.A1(W40982), .A2(W44742), .ZN(O14160));
  NANDX1 G19185 (.A1(W25027), .A2(W28506), .ZN(W44748));
  NANDX1 G19186 (.A1(W914), .A2(W26132), .ZN(O14152));
  NANDX1 G19187 (.A1(W14004), .A2(W10860), .ZN(W44742));
  NANDX1 G19188 (.A1(W11758), .A2(W18544), .ZN(O14151));
  NANDX1 G19189 (.A1(W43311), .A2(W30649), .ZN(O14143));
  NANDX1 G19190 (.A1(W16509), .A2(W41988), .ZN(O14142));
  NANDX1 G19191 (.A1(W28707), .A2(W39257), .ZN(O14127));
  NANDX1 G19192 (.A1(W38046), .A2(W43679), .ZN(O14236));
  NANDX1 G19193 (.A1(W30705), .A2(W11516), .ZN(O14256));
  NANDX1 G19194 (.A1(W40374), .A2(W11275), .ZN(O14255));
  NANDX1 G19195 (.A1(W1770), .A2(W10093), .ZN(O14252));
  NANDX1 G19196 (.A1(W24799), .A2(W29486), .ZN(O14246));
  NANDX1 G19197 (.A1(W35535), .A2(W26310), .ZN(W44863));
  NANDX1 G19198 (.A1(W38744), .A2(W23933), .ZN(O14245));
  NANDX1 G19199 (.A1(W12790), .A2(W17314), .ZN(O14243));
  NANDX1 G19200 (.A1(W6369), .A2(W8736), .ZN(O14242));
  NANDX1 G19201 (.A1(W39420), .A2(W44647), .ZN(O14241));
  NANDX1 G19202 (.A1(W42245), .A2(W27135), .ZN(O14240));
  NANDX1 G19203 (.A1(W41251), .A2(W37005), .ZN(O14237));
  NANDX1 G19204 (.A1(W26348), .A2(W25779), .ZN(O13866));
  NANDX1 G19205 (.A1(W29485), .A2(W24186), .ZN(O14232));
  NANDX1 G19206 (.A1(W9912), .A2(I784), .ZN(O14230));
  NANDX1 G19207 (.A1(W1677), .A2(W28279), .ZN(O14226));
  NANDX1 G19208 (.A1(W21284), .A2(W33558), .ZN(O14225));
  NANDX1 G19209 (.A1(W35984), .A2(W26277), .ZN(O14223));
  NANDX1 G19210 (.A1(W38821), .A2(W38191), .ZN(O14222));
  NANDX1 G19211 (.A1(W27489), .A2(W24692), .ZN(O14219));
  NANDX1 G19212 (.A1(W30753), .A2(W23974), .ZN(O14218));
  NANDX1 G19213 (.A1(W10975), .A2(W6507), .ZN(O14213));
  NANDX1 G19214 (.A1(W25133), .A2(W32560), .ZN(W44821));
  NANDX1 G19215 (.A1(W43353), .A2(W11700), .ZN(O14209));
  NANDX1 G19216 (.A1(W3692), .A2(W31652), .ZN(W43981));
  NANDX1 G19217 (.A1(W4264), .A2(W2515), .ZN(O13562));
  NANDX1 G19218 (.A1(W4802), .A2(W5460), .ZN(O13561));
  NANDX1 G19219 (.A1(W21144), .A2(W2868), .ZN(O13560));
  NANDX1 G19220 (.A1(W1545), .A2(W3570), .ZN(O13558));
  NANDX1 G19221 (.A1(W28964), .A2(W38728), .ZN(W44007));
  NANDX1 G19222 (.A1(I1212), .A2(W41835), .ZN(O13553));
  NANDX1 G19223 (.A1(W40558), .A2(W34481), .ZN(O13552));
  NANDX1 G19224 (.A1(W17866), .A2(W24505), .ZN(W43999));
  NANDX1 G19225 (.A1(W1665), .A2(W5762), .ZN(O13550));
  NANDX1 G19226 (.A1(W4), .A2(W27310), .ZN(O13545));
  NANDX1 G19227 (.A1(W41616), .A2(W27470), .ZN(O13539));
  NANDX1 G19228 (.A1(W1971), .A2(W1566), .ZN(W43982));
  NANDX1 G19229 (.A1(W38711), .A2(W9479), .ZN(W44015));
  NANDX1 G19230 (.A1(W2814), .A2(W29211), .ZN(O13537));
  NANDX1 G19231 (.A1(W35189), .A2(W15424), .ZN(O13530));
  NANDX1 G19232 (.A1(W15401), .A2(I1510), .ZN(O13528));
  NANDX1 G19233 (.A1(W10754), .A2(W8445), .ZN(O13524));
  NANDX1 G19234 (.A1(W2952), .A2(W19630), .ZN(O13521));
  NANDX1 G19235 (.A1(W18561), .A2(W22983), .ZN(O13518));
  NANDX1 G19236 (.A1(W41720), .A2(W4218), .ZN(W43957));
  NANDX1 G19237 (.A1(W41820), .A2(W16439), .ZN(O13517));
  NANDX1 G19238 (.A1(W26971), .A2(W36760), .ZN(O13515));
  NANDX1 G19239 (.A1(W33553), .A2(W32565), .ZN(O13512));
  NANDX1 G19240 (.A1(W18204), .A2(W17328), .ZN(O13506));
  NANDX1 G19241 (.A1(W28579), .A2(W42252), .ZN(O13597));
  NANDX1 G19242 (.A1(W24634), .A2(W24815), .ZN(O13622));
  NANDX1 G19243 (.A1(W20007), .A2(W34057), .ZN(W44088));
  NANDX1 G19244 (.A1(W11477), .A2(W2502), .ZN(W44086));
  NANDX1 G19245 (.A1(W33887), .A2(W38090), .ZN(W44083));
  NANDX1 G19246 (.A1(W24781), .A2(W5953), .ZN(O13617));
  NANDX1 G19247 (.A1(W19561), .A2(W7728), .ZN(O13615));
  NANDX1 G19248 (.A1(W36260), .A2(W25159), .ZN(O13614));
  NANDX1 G19249 (.A1(W27765), .A2(W15845), .ZN(O13613));
  NANDX1 G19250 (.A1(W7821), .A2(W10419), .ZN(W44071));
  NANDX1 G19251 (.A1(W43765), .A2(W40133), .ZN(O13608));
  NANDX1 G19252 (.A1(W20613), .A2(W25492), .ZN(O13603));
  NANDX1 G19253 (.A1(W29782), .A2(W24059), .ZN(O13600));
  NANDX1 G19254 (.A1(W38750), .A2(W5878), .ZN(O13504));
  NANDX1 G19255 (.A1(W27872), .A2(W28419), .ZN(O13595));
  NANDX1 G19256 (.A1(W39484), .A2(W19460), .ZN(O13594));
  NANDX1 G19257 (.A1(W35053), .A2(W8267), .ZN(W44053));
  NANDX1 G19258 (.A1(W5141), .A2(W16074), .ZN(O13590));
  NANDX1 G19259 (.A1(W32665), .A2(W24169), .ZN(O13589));
  NANDX1 G19260 (.A1(W38184), .A2(I1571), .ZN(O13582));
  NANDX1 G19261 (.A1(W15727), .A2(W13089), .ZN(O13580));
  NANDX1 G19262 (.A1(W1335), .A2(W43630), .ZN(O13579));
  NANDX1 G19263 (.A1(W10584), .A2(I1826), .ZN(W44034));
  NANDX1 G19264 (.A1(W21125), .A2(W29225), .ZN(O13572));
  NANDX1 G19265 (.A1(I512), .A2(W41986), .ZN(O13565));
  NANDX1 G19266 (.A1(W7293), .A2(W35300), .ZN(W43818));
  NANDX1 G19267 (.A1(W40864), .A2(W19488), .ZN(O13436));
  NANDX1 G19268 (.A1(W42922), .A2(W26860), .ZN(O13434));
  NANDX1 G19269 (.A1(W1064), .A2(W9230), .ZN(O13431));
  NANDX1 G19270 (.A1(W3149), .A2(W87), .ZN(W43845));
  NANDX1 G19271 (.A1(W32760), .A2(W41807), .ZN(O13427));
  NANDX1 G19272 (.A1(W8772), .A2(W30443), .ZN(W43838));
  NANDX1 G19273 (.A1(W17873), .A2(W26583), .ZN(O13421));
  NANDX1 G19274 (.A1(W21563), .A2(W23816), .ZN(W43832));
  NANDX1 G19275 (.A1(W7746), .A2(W9887), .ZN(W43825));
  NANDX1 G19276 (.A1(W6155), .A2(W27719), .ZN(O13414));
  NANDX1 G19277 (.A1(W16305), .A2(W17281), .ZN(O13412));
  NANDX1 G19278 (.A1(W35433), .A2(W196), .ZN(W43819));
  NANDX1 G19279 (.A1(I272), .A2(W9756), .ZN(O13438));
  NANDX1 G19280 (.A1(W34960), .A2(W33734), .ZN(W43815));
  NANDX1 G19281 (.A1(W38300), .A2(W43532), .ZN(O13408));
  NANDX1 G19282 (.A1(W27598), .A2(W28098), .ZN(W43813));
  NANDX1 G19283 (.A1(W38670), .A2(W38632), .ZN(O13405));
  NANDX1 G19284 (.A1(W25675), .A2(W23756), .ZN(O13404));
  NANDX1 G19285 (.A1(W18974), .A2(W12675), .ZN(O13402));
  NANDX1 G19286 (.A1(I765), .A2(W19406), .ZN(O13400));
  NANDX1 G19287 (.A1(W17711), .A2(W37844), .ZN(O13399));
  NANDX1 G19288 (.A1(W29667), .A2(W9863), .ZN(O13397));
  NANDX1 G19289 (.A1(W26377), .A2(W2128), .ZN(W43798));
  NANDX1 G19290 (.A1(W41686), .A2(W23058), .ZN(O13394));
  NANDX1 G19291 (.A1(W26355), .A2(W26958), .ZN(O13480));
  NANDX1 G19292 (.A1(W1976), .A2(I1056), .ZN(O13499));
  NANDX1 G19293 (.A1(W41973), .A2(W2567), .ZN(W43932));
  NANDX1 G19294 (.A1(W7372), .A2(W13830), .ZN(O13497));
  NANDX1 G19295 (.A1(W23307), .A2(W24774), .ZN(W43930));
  NANDX1 G19296 (.A1(W8734), .A2(W34261), .ZN(O13496));
  NANDX1 G19297 (.A1(W9271), .A2(W43886), .ZN(W43928));
  NANDX1 G19298 (.A1(W23233), .A2(W34030), .ZN(O13495));
  NANDX1 G19299 (.A1(W14773), .A2(W40460), .ZN(W43926));
  NANDX1 G19300 (.A1(W36067), .A2(W43579), .ZN(O13492));
  NANDX1 G19301 (.A1(W32275), .A2(W10397), .ZN(O13488));
  NANDX1 G19302 (.A1(W32576), .A2(W12186), .ZN(O13483));
  NANDX1 G19303 (.A1(W20400), .A2(W31746), .ZN(W44091));
  NANDX1 G19304 (.A1(W23110), .A2(W23433), .ZN(O13478));
  NANDX1 G19305 (.A1(W26822), .A2(W38638), .ZN(O13470));
  NANDX1 G19306 (.A1(W22051), .A2(W27919), .ZN(O13469));
  NANDX1 G19307 (.A1(W24784), .A2(W43848), .ZN(W43884));
  NANDX1 G19308 (.A1(W27313), .A2(W639), .ZN(O13459));
  NANDX1 G19309 (.A1(I1428), .A2(W26010), .ZN(O13458));
  NANDX1 G19310 (.A1(W17379), .A2(W24505), .ZN(O13456));
  NANDX1 G19311 (.A1(W16792), .A2(W11507), .ZN(O13449));
  NANDX1 G19312 (.A1(W9447), .A2(W35449), .ZN(W43862));
  NANDX1 G19313 (.A1(I1374), .A2(W24081), .ZN(O13442));
  NANDX1 G19314 (.A1(W38181), .A2(W28545), .ZN(O13441));
  NANDX1 G19315 (.A1(W1624), .A2(W35096), .ZN(O13787));
  NANDX1 G19316 (.A1(W21286), .A2(W40976), .ZN(W44336));
  NANDX1 G19317 (.A1(W40260), .A2(W28838), .ZN(O13820));
  NANDX1 G19318 (.A1(W29773), .A2(W16273), .ZN(O13817));
  NANDX1 G19319 (.A1(W34865), .A2(W10803), .ZN(O13815));
  NANDX1 G19320 (.A1(W21076), .A2(W10515), .ZN(O13814));
  NANDX1 G19321 (.A1(W26623), .A2(W34837), .ZN(O13812));
  NANDX1 G19322 (.A1(I1350), .A2(W12303), .ZN(O13807));
  NANDX1 G19323 (.A1(W8697), .A2(W4082), .ZN(O13806));
  NANDX1 G19324 (.A1(W19130), .A2(W12101), .ZN(O13801));
  NANDX1 G19325 (.A1(W4759), .A2(W38333), .ZN(O13800));
  NANDX1 G19326 (.A1(W42063), .A2(W34540), .ZN(W44312));
  NANDX1 G19327 (.A1(W13119), .A2(W11707), .ZN(O13795));
  NANDX1 G19328 (.A1(W17065), .A2(W3709), .ZN(O13821));
  NANDX1 G19329 (.A1(W17947), .A2(W36731), .ZN(O13786));
  NANDX1 G19330 (.A1(W21152), .A2(W30692), .ZN(O13777));
  NANDX1 G19331 (.A1(W42267), .A2(W30110), .ZN(O13770));
  NANDX1 G19332 (.A1(W32174), .A2(W27152), .ZN(O13769));
  NANDX1 G19333 (.A1(W4389), .A2(W17080), .ZN(O13768));
  NANDX1 G19334 (.A1(W14249), .A2(W6493), .ZN(O13764));
  NANDX1 G19335 (.A1(W22772), .A2(W36339), .ZN(O13757));
  NANDX1 G19336 (.A1(W6214), .A2(W8660), .ZN(O13745));
  NANDX1 G19337 (.A1(W22557), .A2(W31113), .ZN(O13744));
  NANDX1 G19338 (.A1(W22778), .A2(I1524), .ZN(O13733));
  NANDX1 G19339 (.A1(W11680), .A2(W41678), .ZN(W44231));
  NANDX1 G19340 (.A1(W14091), .A2(W8973), .ZN(O13843));
  NANDX1 G19341 (.A1(W34932), .A2(W42267), .ZN(O13864));
  NANDX1 G19342 (.A1(W8421), .A2(W23644), .ZN(W44391));
  NANDX1 G19343 (.A1(W18971), .A2(W27036), .ZN(W44386));
  NANDX1 G19344 (.A1(W231), .A2(W34561), .ZN(O13860));
  NANDX1 G19345 (.A1(W37287), .A2(W40371), .ZN(W44383));
  NANDX1 G19346 (.A1(W1086), .A2(W20091), .ZN(O13857));
  NANDX1 G19347 (.A1(W31086), .A2(W3802), .ZN(O13856));
  NANDX1 G19348 (.A1(W37896), .A2(W15009), .ZN(O13854));
  NANDX1 G19349 (.A1(I1966), .A2(W42477), .ZN(O13852));
  NANDX1 G19350 (.A1(W33158), .A2(W35040), .ZN(O13851));
  NANDX1 G19351 (.A1(W36962), .A2(W3646), .ZN(O13847));
  NANDX1 G19352 (.A1(W37579), .A2(W22673), .ZN(O13846));
  NANDX1 G19353 (.A1(W39965), .A2(W27141), .ZN(O13730));
  NANDX1 G19354 (.A1(W9447), .A2(W14828), .ZN(O13842));
  NANDX1 G19355 (.A1(W15465), .A2(W36791), .ZN(O13841));
  NANDX1 G19356 (.A1(I1714), .A2(W5078), .ZN(O13838));
  NANDX1 G19357 (.A1(W41637), .A2(W21922), .ZN(O13837));
  NANDX1 G19358 (.A1(W33395), .A2(W7236), .ZN(O13834));
  NANDX1 G19359 (.A1(W18921), .A2(W35282), .ZN(O13832));
  NANDX1 G19360 (.A1(W43999), .A2(W37355), .ZN(O13828));
  NANDX1 G19361 (.A1(W40396), .A2(W32714), .ZN(O13827));
  NANDX1 G19362 (.A1(W29440), .A2(W11680), .ZN(O13826));
  NANDX1 G19363 (.A1(W24941), .A2(W6976), .ZN(O13825));
  NANDX1 G19364 (.A1(W13444), .A2(W24746), .ZN(O13824));
  NANDX1 G19365 (.A1(W32528), .A2(W1065), .ZN(O13654));
  NANDX1 G19366 (.A1(W12295), .A2(I375), .ZN(O13684));
  NANDX1 G19367 (.A1(I816), .A2(W31253), .ZN(O13681));
  NANDX1 G19368 (.A1(W3597), .A2(W43807), .ZN(W44166));
  NANDX1 G19369 (.A1(W25543), .A2(W16794), .ZN(W44163));
  NANDX1 G19370 (.A1(W10744), .A2(W29426), .ZN(O13673));
  NANDX1 G19371 (.A1(W10775), .A2(W13002), .ZN(O13670));
  NANDX1 G19372 (.A1(W12739), .A2(W13700), .ZN(O13669));
  NANDX1 G19373 (.A1(I207), .A2(W17327), .ZN(W44143));
  NANDX1 G19374 (.A1(W18789), .A2(W18568), .ZN(W44141));
  NANDX1 G19375 (.A1(W13657), .A2(W9629), .ZN(W44135));
  NANDX1 G19376 (.A1(W26801), .A2(W23533), .ZN(O13661));
  NANDX1 G19377 (.A1(W14567), .A2(W22029), .ZN(O13657));
  NANDX1 G19378 (.A1(W30109), .A2(W17089), .ZN(O13691));
  NANDX1 G19379 (.A1(W22616), .A2(W43155), .ZN(O13652));
  NANDX1 G19380 (.A1(W37493), .A2(W30001), .ZN(O13651));
  NANDX1 G19381 (.A1(W8121), .A2(W42614), .ZN(O13642));
  NANDX1 G19382 (.A1(W8211), .A2(W1450), .ZN(O13638));
  NANDX1 G19383 (.A1(W19297), .A2(W17918), .ZN(O13630));
  NANDX1 G19384 (.A1(W42958), .A2(W43488), .ZN(O13629));
  NANDX1 G19385 (.A1(W33921), .A2(W2219), .ZN(W44096));
  NANDX1 G19386 (.A1(W3029), .A2(W32048), .ZN(O13626));
  NANDX1 G19387 (.A1(W6410), .A2(W7763), .ZN(O13625));
  NANDX1 G19388 (.A1(I493), .A2(W34099), .ZN(O13624));
  NANDX1 G19389 (.A1(W24987), .A2(W25545), .ZN(W44092));
  NANDX1 G19390 (.A1(W21056), .A2(W20751), .ZN(O13710));
  NANDX1 G19391 (.A1(W25565), .A2(W7198), .ZN(O13729));
  NANDX1 G19392 (.A1(W43178), .A2(W32075), .ZN(W44225));
  NANDX1 G19393 (.A1(I937), .A2(W12059), .ZN(O13727));
  NANDX1 G19394 (.A1(W17630), .A2(W30587), .ZN(O13724));
  NANDX1 G19395 (.A1(W25418), .A2(W5795), .ZN(O13720));
  NANDX1 G19396 (.A1(W4861), .A2(W6832), .ZN(O13719));
  NANDX1 G19397 (.A1(W32112), .A2(W38987), .ZN(W44214));
  NANDX1 G19398 (.A1(W38488), .A2(W35308), .ZN(O13718));
  NANDX1 G19399 (.A1(W19446), .A2(W31328), .ZN(O13715));
  NANDX1 G19400 (.A1(W11405), .A2(W37628), .ZN(O13714));
  NANDX1 G19401 (.A1(W38881), .A2(W21753), .ZN(O13711));
  NANDX1 G19402 (.A1(W18794), .A2(W260), .ZN(O14368));
  NANDX1 G19403 (.A1(W22220), .A2(W3839), .ZN(O13709));
  NANDX1 G19404 (.A1(W37293), .A2(I746), .ZN(O13708));
  NANDX1 G19405 (.A1(W36602), .A2(W38), .ZN(O13707));
  NANDX1 G19406 (.A1(W31207), .A2(W21727), .ZN(O13705));
  NANDX1 G19407 (.A1(W7585), .A2(W34522), .ZN(O13704));
  NANDX1 G19408 (.A1(W16999), .A2(I1392), .ZN(O13703));
  NANDX1 G19409 (.A1(W22229), .A2(W11962), .ZN(O13699));
  NANDX1 G19410 (.A1(W27883), .A2(W26289), .ZN(W44185));
  NANDX1 G19411 (.A1(W11194), .A2(W5555), .ZN(O13694));
  NANDX1 G19412 (.A1(I521), .A2(W5420), .ZN(W44182));
  NANDX1 G19413 (.A1(W2045), .A2(W33782), .ZN(O13692));
  NANDX1 G19414 (.A1(W36598), .A2(W22948), .ZN(O15018));
  NANDX1 G19415 (.A1(W27283), .A2(W16236), .ZN(O15039));
  NANDX1 G19416 (.A1(I324), .A2(W43575), .ZN(O15037));
  NANDX1 G19417 (.A1(W13394), .A2(W38644), .ZN(O15036));
  NANDX1 G19418 (.A1(W31633), .A2(W10479), .ZN(W45822));
  NANDX1 G19419 (.A1(W767), .A2(W26431), .ZN(W45821));
  NANDX1 G19420 (.A1(W42707), .A2(W10), .ZN(O15035));
  NANDX1 G19421 (.A1(W32927), .A2(W43838), .ZN(O15032));
  NANDX1 G19422 (.A1(W40542), .A2(W5725), .ZN(O15031));
  NANDX1 G19423 (.A1(W7020), .A2(W20064), .ZN(O15030));
  NANDX1 G19424 (.A1(W7712), .A2(W28441), .ZN(O15029));
  NANDX1 G19425 (.A1(W12596), .A2(W18345), .ZN(O15028));
  NANDX1 G19426 (.A1(W30842), .A2(W25673), .ZN(O15024));
  NANDX1 G19427 (.A1(W32248), .A2(W32914), .ZN(O15040));
  NANDX1 G19428 (.A1(W5716), .A2(W1998), .ZN(O15013));
  NANDX1 G19429 (.A1(W32575), .A2(W8795), .ZN(W45792));
  NANDX1 G19430 (.A1(W44790), .A2(W11938), .ZN(O15010));
  NANDX1 G19431 (.A1(W28122), .A2(W24110), .ZN(O15009));
  NANDX1 G19432 (.A1(W1829), .A2(W33148), .ZN(O15008));
  NANDX1 G19433 (.A1(W20457), .A2(W2970), .ZN(W45788));
  NANDX1 G19434 (.A1(W16205), .A2(W18444), .ZN(O15004));
  NANDX1 G19435 (.A1(W11088), .A2(W34443), .ZN(O15003));
  NANDX1 G19436 (.A1(W31064), .A2(W7131), .ZN(O15001));
  NANDX1 G19437 (.A1(W14990), .A2(W9071), .ZN(W45779));
  NANDX1 G19438 (.A1(W15458), .A2(W43759), .ZN(O14994));
  NANDX1 G19439 (.A1(W20028), .A2(W32772), .ZN(O15075));
  NANDX1 G19440 (.A1(W35797), .A2(W28004), .ZN(O15108));
  NANDX1 G19441 (.A1(W19339), .A2(W23258), .ZN(O15106));
  NANDX1 G19442 (.A1(W1930), .A2(W29717), .ZN(W45907));
  NANDX1 G19443 (.A1(W18275), .A2(W7523), .ZN(O15102));
  NANDX1 G19444 (.A1(W38502), .A2(W38750), .ZN(O15101));
  NANDX1 G19445 (.A1(W22536), .A2(W11076), .ZN(W45902));
  NANDX1 G19446 (.A1(W41732), .A2(W9851), .ZN(O15098));
  NANDX1 G19447 (.A1(W24409), .A2(W8900), .ZN(O15097));
  NANDX1 G19448 (.A1(W45411), .A2(W37620), .ZN(O15093));
  NANDX1 G19449 (.A1(W38108), .A2(W37649), .ZN(O15092));
  NANDX1 G19450 (.A1(W41762), .A2(W4117), .ZN(O15090));
  NANDX1 G19451 (.A1(W16300), .A2(W37372), .ZN(O15076));
  NANDX1 G19452 (.A1(W19881), .A2(W17584), .ZN(O14993));
  NANDX1 G19453 (.A1(W26789), .A2(W30502), .ZN(O15068));
  NANDX1 G19454 (.A1(W24862), .A2(W9936), .ZN(O15066));
  NANDX1 G19455 (.A1(W34325), .A2(W8305), .ZN(W45861));
  NANDX1 G19456 (.A1(W15588), .A2(W31471), .ZN(O15064));
  NANDX1 G19457 (.A1(W5579), .A2(W11568), .ZN(W45853));
  NANDX1 G19458 (.A1(W45692), .A2(W35), .ZN(O15060));
  NANDX1 G19459 (.A1(W39346), .A2(W14473), .ZN(O15056));
  NANDX1 G19460 (.A1(W23411), .A2(W2354), .ZN(O15055));
  NANDX1 G19461 (.A1(W11974), .A2(W42540), .ZN(O15053));
  NANDX1 G19462 (.A1(W16636), .A2(W33457), .ZN(W45836));
  NANDX1 G19463 (.A1(W44662), .A2(W18650), .ZN(O15043));
  NANDX1 G19464 (.A1(W26164), .A2(W36263), .ZN(O14887));
  NANDX1 G19465 (.A1(W17026), .A2(W34730), .ZN(O14918));
  NANDX1 G19466 (.A1(W28989), .A2(W12103), .ZN(O14913));
  NANDX1 G19467 (.A1(W36673), .A2(W677), .ZN(O14911));
  NANDX1 G19468 (.A1(W19807), .A2(W12872), .ZN(O14910));
  NANDX1 G19469 (.A1(W18014), .A2(W20812), .ZN(O14909));
  NANDX1 G19470 (.A1(W8955), .A2(W28100), .ZN(O14906));
  NANDX1 G19471 (.A1(W44942), .A2(W1825), .ZN(O14905));
  NANDX1 G19472 (.A1(W37545), .A2(W2444), .ZN(O14904));
  NANDX1 G19473 (.A1(W21896), .A2(W7571), .ZN(O14903));
  NANDX1 G19474 (.A1(W24146), .A2(W12772), .ZN(W45656));
  NANDX1 G19475 (.A1(W1434), .A2(W9819), .ZN(O14893));
  NANDX1 G19476 (.A1(W22339), .A2(W21704), .ZN(O14892));
  NANDX1 G19477 (.A1(W25562), .A2(W35840), .ZN(O14922));
  NANDX1 G19478 (.A1(W42251), .A2(W18437), .ZN(O14886));
  NANDX1 G19479 (.A1(W19802), .A2(W42172), .ZN(W45639));
  NANDX1 G19480 (.A1(W31249), .A2(W17857), .ZN(O14883));
  NANDX1 G19481 (.A1(W16611), .A2(W6667), .ZN(O14882));
  NANDX1 G19482 (.A1(W31125), .A2(W34886), .ZN(O14873));
  NANDX1 G19483 (.A1(W43291), .A2(W40860), .ZN(W45625));
  NANDX1 G19484 (.A1(W30262), .A2(W1815), .ZN(O14869));
  NANDX1 G19485 (.A1(W30461), .A2(W16209), .ZN(O14867));
  NANDX1 G19486 (.A1(W14398), .A2(W39699), .ZN(O14861));
  NANDX1 G19487 (.A1(W35539), .A2(W15603), .ZN(O14860));
  NANDX1 G19488 (.A1(W41329), .A2(W987), .ZN(O14858));
  NANDX1 G19489 (.A1(W7190), .A2(W22357), .ZN(O14952));
  NANDX1 G19490 (.A1(W9680), .A2(W26911), .ZN(O14990));
  NANDX1 G19491 (.A1(W29311), .A2(W44862), .ZN(O14989));
  NANDX1 G19492 (.A1(W41343), .A2(W34211), .ZN(O14988));
  NANDX1 G19493 (.A1(W24932), .A2(W20860), .ZN(O14986));
  NANDX1 G19494 (.A1(W27153), .A2(W27846), .ZN(O14984));
  NANDX1 G19495 (.A1(W38356), .A2(W33397), .ZN(O14983));
  NANDX1 G19496 (.A1(W11795), .A2(W34736), .ZN(O14973));
  NANDX1 G19497 (.A1(W8530), .A2(W22251), .ZN(O14971));
  NANDX1 G19498 (.A1(W27968), .A2(W16699), .ZN(O14970));
  NANDX1 G19499 (.A1(W36824), .A2(W4362), .ZN(O14954));
  NANDX1 G19500 (.A1(W12273), .A2(W6159), .ZN(O14953));
  NANDX1 G19501 (.A1(W15888), .A2(W31112), .ZN(O15109));
  NANDX1 G19502 (.A1(I587), .A2(W26369), .ZN(W45718));
  NANDX1 G19503 (.A1(W2966), .A2(W20550), .ZN(O14949));
  NANDX1 G19504 (.A1(W27804), .A2(W44239), .ZN(W45715));
  NANDX1 G19505 (.A1(W25962), .A2(W10988), .ZN(O14944));
  NANDX1 G19506 (.A1(W42772), .A2(W26328), .ZN(O14940));
  NANDX1 G19507 (.A1(W5363), .A2(W19733), .ZN(O14939));
  NANDX1 G19508 (.A1(W2126), .A2(W7688), .ZN(O14938));
  NANDX1 G19509 (.A1(W10030), .A2(W33335), .ZN(O14936));
  NANDX1 G19510 (.A1(W25385), .A2(W2853), .ZN(O14930));
  NANDX1 G19511 (.A1(W37869), .A2(W3850), .ZN(O14927));
  NANDX1 G19512 (.A1(W15573), .A2(W42106), .ZN(O14925));
  NANDX1 G19513 (.A1(W19536), .A2(W28133), .ZN(O15266));
  NANDX1 G19514 (.A1(W2002), .A2(W39879), .ZN(O15297));
  NANDX1 G19515 (.A1(W25260), .A2(W44774), .ZN(O15296));
  NANDX1 G19516 (.A1(W1230), .A2(W18828), .ZN(O15293));
  NANDX1 G19517 (.A1(W22893), .A2(W22397), .ZN(O15291));
  NANDX1 G19518 (.A1(W37836), .A2(W15752), .ZN(W46135));
  NANDX1 G19519 (.A1(W20148), .A2(W45429), .ZN(O15286));
  NANDX1 G19520 (.A1(W22678), .A2(W5344), .ZN(O15284));
  NANDX1 G19521 (.A1(W45135), .A2(W42660), .ZN(O15278));
  NANDX1 G19522 (.A1(W27637), .A2(W38464), .ZN(W46124));
  NANDX1 G19523 (.A1(I1404), .A2(W33845), .ZN(O15276));
  NANDX1 G19524 (.A1(W2267), .A2(W32437), .ZN(O15270));
  NANDX1 G19525 (.A1(W27563), .A2(W46053), .ZN(W46110));
  NANDX1 G19526 (.A1(W26841), .A2(W28366), .ZN(O15300));
  NANDX1 G19527 (.A1(W21444), .A2(W4014), .ZN(O15262));
  NANDX1 G19528 (.A1(W17065), .A2(W23893), .ZN(O15260));
  NANDX1 G19529 (.A1(W27763), .A2(W30631), .ZN(O15255));
  NANDX1 G19530 (.A1(W15400), .A2(W30098), .ZN(O15254));
  NANDX1 G19531 (.A1(I1444), .A2(W43930), .ZN(O15252));
  NANDX1 G19532 (.A1(W34626), .A2(W5563), .ZN(O15251));
  NANDX1 G19533 (.A1(W73), .A2(W1641), .ZN(O15249));
  NANDX1 G19534 (.A1(W35216), .A2(W22563), .ZN(O15245));
  NANDX1 G19535 (.A1(W38650), .A2(W14962), .ZN(W46079));
  NANDX1 G19536 (.A1(W24690), .A2(W17729), .ZN(W46078));
  NANDX1 G19537 (.A1(W41171), .A2(W9654), .ZN(O15242));
  NANDX1 G19538 (.A1(W42816), .A2(W41478), .ZN(O15339));
  NANDX1 G19539 (.A1(W29789), .A2(W12221), .ZN(O15369));
  NANDX1 G19540 (.A1(W12076), .A2(W45119), .ZN(O15365));
  NANDX1 G19541 (.A1(W1740), .A2(W5855), .ZN(O15364));
  NANDX1 G19542 (.A1(I1593), .A2(W1211), .ZN(O15359));
  NANDX1 G19543 (.A1(W42324), .A2(W26272), .ZN(W46218));
  NANDX1 G19544 (.A1(W12072), .A2(W20320), .ZN(O15358));
  NANDX1 G19545 (.A1(W23877), .A2(W33425), .ZN(W46213));
  NANDX1 G19546 (.A1(I1240), .A2(I1154), .ZN(O15352));
  NANDX1 G19547 (.A1(I1008), .A2(W17561), .ZN(O15351));
  NANDX1 G19548 (.A1(W37653), .A2(W5669), .ZN(O15350));
  NANDX1 G19549 (.A1(W40066), .A2(W45033), .ZN(O15348));
  NANDX1 G19550 (.A1(W33405), .A2(I1293), .ZN(O15341));
  NANDX1 G19551 (.A1(W24329), .A2(W42717), .ZN(O15237));
  NANDX1 G19552 (.A1(W19860), .A2(I44), .ZN(O15336));
  NANDX1 G19553 (.A1(W519), .A2(W22388), .ZN(O15335));
  NANDX1 G19554 (.A1(W36233), .A2(W33771), .ZN(O15334));
  NANDX1 G19555 (.A1(I1566), .A2(W11951), .ZN(O15330));
  NANDX1 G19556 (.A1(W18069), .A2(W17778), .ZN(O15320));
  NANDX1 G19557 (.A1(W7237), .A2(W38416), .ZN(O15318));
  NANDX1 G19558 (.A1(W21287), .A2(W7133), .ZN(W46164));
  NANDX1 G19559 (.A1(W2314), .A2(W12022), .ZN(O15312));
  NANDX1 G19560 (.A1(W24596), .A2(W19329), .ZN(O15307));
  NANDX1 G19561 (.A1(W11175), .A2(W7947), .ZN(O15306));
  NANDX1 G19562 (.A1(W24238), .A2(W38135), .ZN(O15303));
  NANDX1 G19563 (.A1(W9056), .A2(W16639), .ZN(O15135));
  NANDX1 G19564 (.A1(W39646), .A2(W19286), .ZN(O15171));
  NANDX1 G19565 (.A1(W7190), .A2(W16258), .ZN(O15167));
  NANDX1 G19566 (.A1(W4777), .A2(W19565), .ZN(W45988));
  NANDX1 G19567 (.A1(W15048), .A2(W24748), .ZN(O15164));
  NANDX1 G19568 (.A1(W13231), .A2(W13777), .ZN(W45984));
  NANDX1 G19569 (.A1(W18465), .A2(W2524), .ZN(O15163));
  NANDX1 G19570 (.A1(W26668), .A2(W26100), .ZN(W45977));
  NANDX1 G19571 (.A1(W35016), .A2(W20102), .ZN(O15157));
  NANDX1 G19572 (.A1(W17273), .A2(W38180), .ZN(O15156));
  NANDX1 G19573 (.A1(W25746), .A2(W28152), .ZN(O15155));
  NANDX1 G19574 (.A1(W6197), .A2(W32867), .ZN(O15143));
  NANDX1 G19575 (.A1(W13188), .A2(W41483), .ZN(W45951));
  NANDX1 G19576 (.A1(W22931), .A2(W8248), .ZN(O15173));
  NANDX1 G19577 (.A1(W1755), .A2(W21997), .ZN(O15134));
  NANDX1 G19578 (.A1(W21693), .A2(W6050), .ZN(O15132));
  NANDX1 G19579 (.A1(W4524), .A2(I535), .ZN(O15128));
  NANDX1 G19580 (.A1(W45594), .A2(I374), .ZN(O15125));
  NANDX1 G19581 (.A1(W27744), .A2(W14582), .ZN(O15123));
  NANDX1 G19582 (.A1(W15945), .A2(W9987), .ZN(O15121));
  NANDX1 G19583 (.A1(W12417), .A2(W12953), .ZN(O15116));
  NANDX1 G19584 (.A1(W27998), .A2(W25422), .ZN(O15115));
  NANDX1 G19585 (.A1(W38807), .A2(W13277), .ZN(W45920));
  NANDX1 G19586 (.A1(W26016), .A2(W26438), .ZN(O15112));
  NANDX1 G19587 (.A1(W1961), .A2(W37158), .ZN(O15110));
  NANDX1 G19588 (.A1(W25462), .A2(W33288), .ZN(O15211));
  NANDX1 G19589 (.A1(W6546), .A2(W12677), .ZN(O15235));
  NANDX1 G19590 (.A1(W27391), .A2(W38236), .ZN(O15231));
  NANDX1 G19591 (.A1(W32511), .A2(W5997), .ZN(O15223));
  NANDX1 G19592 (.A1(W6933), .A2(W19048), .ZN(W46053));
  NANDX1 G19593 (.A1(W6321), .A2(W39757), .ZN(O15219));
  NANDX1 G19594 (.A1(W2853), .A2(W8452), .ZN(O15217));
  NANDX1 G19595 (.A1(W44031), .A2(W1168), .ZN(O15216));
  NANDX1 G19596 (.A1(W1427), .A2(W17530), .ZN(O15215));
  NANDX1 G19597 (.A1(W38965), .A2(W29521), .ZN(O15214));
  NANDX1 G19598 (.A1(W20026), .A2(W42237), .ZN(O15213));
  NANDX1 G19599 (.A1(W33557), .A2(W8974), .ZN(O15212));
  NANDX1 G19600 (.A1(W27071), .A2(W9304), .ZN(O14856));
  NANDX1 G19601 (.A1(W17612), .A2(W1771), .ZN(O15205));
  NANDX1 G19602 (.A1(W13803), .A2(I921), .ZN(O15203));
  NANDX1 G19603 (.A1(W12105), .A2(W14904), .ZN(O15201));
  NANDX1 G19604 (.A1(W25830), .A2(W25115), .ZN(O15197));
  NANDX1 G19605 (.A1(I543), .A2(W812), .ZN(O15194));
  NANDX1 G19606 (.A1(W34197), .A2(W7228), .ZN(O15191));
  NANDX1 G19607 (.A1(W18510), .A2(W31073), .ZN(O15188));
  NANDX1 G19608 (.A1(W8485), .A2(W32090), .ZN(O15185));
  NANDX1 G19609 (.A1(I722), .A2(W36709), .ZN(O15184));
  NANDX1 G19610 (.A1(W12245), .A2(W24495), .ZN(O15177));
  NANDX1 G19611 (.A1(W33687), .A2(W1991), .ZN(O15176));
  NANDX1 G19612 (.A1(W3113), .A2(W4452), .ZN(O14518));
  NANDX1 G19613 (.A1(W36341), .A2(W1171), .ZN(O14542));
  NANDX1 G19614 (.A1(W36659), .A2(W33477), .ZN(O14541));
  NANDX1 G19615 (.A1(W18801), .A2(W603), .ZN(O14539));
  NANDX1 G19616 (.A1(W387), .A2(W30444), .ZN(O14535));
  NANDX1 G19617 (.A1(W39258), .A2(W4753), .ZN(O14534));
  NANDX1 G19618 (.A1(W10713), .A2(W999), .ZN(O14533));
  NANDX1 G19619 (.A1(W19230), .A2(W10961), .ZN(W45206));
  NANDX1 G19620 (.A1(W20231), .A2(W41645), .ZN(O14528));
  NANDX1 G19621 (.A1(W19994), .A2(W25031), .ZN(O14527));
  NANDX1 G19622 (.A1(W36140), .A2(W20940), .ZN(O14523));
  NANDX1 G19623 (.A1(W3862), .A2(W42955), .ZN(O14521));
  NANDX1 G19624 (.A1(W20358), .A2(W2789), .ZN(O14519));
  NANDX1 G19625 (.A1(W14266), .A2(W40032), .ZN(O14550));
  NANDX1 G19626 (.A1(W22932), .A2(W36165), .ZN(O14517));
  NANDX1 G19627 (.A1(I1761), .A2(W32136), .ZN(O14516));
  NANDX1 G19628 (.A1(W30147), .A2(W34722), .ZN(O14513));
  NANDX1 G19629 (.A1(W16303), .A2(W32649), .ZN(O14503));
  NANDX1 G19630 (.A1(W32293), .A2(W19453), .ZN(O14501));
  NANDX1 G19631 (.A1(W9363), .A2(W23555), .ZN(O14500));
  NANDX1 G19632 (.A1(W31566), .A2(W25851), .ZN(W45171));
  NANDX1 G19633 (.A1(W24150), .A2(W33603), .ZN(O14499));
  NANDX1 G19634 (.A1(W365), .A2(W12083), .ZN(O14497));
  NANDX1 G19635 (.A1(W39728), .A2(W18951), .ZN(O14489));
  NANDX1 G19636 (.A1(W29282), .A2(W44742), .ZN(O14487));
  NANDX1 G19637 (.A1(W13190), .A2(W13646), .ZN(O14584));
  NANDX1 G19638 (.A1(W15586), .A2(W45149), .ZN(O14611));
  NANDX1 G19639 (.A1(W24578), .A2(W28907), .ZN(O14606));
  NANDX1 G19640 (.A1(W36665), .A2(W37350), .ZN(O14605));
  NANDX1 G19641 (.A1(W41229), .A2(W20449), .ZN(W45302));
  NANDX1 G19642 (.A1(W22006), .A2(W37648), .ZN(O14602));
  NANDX1 G19643 (.A1(W7155), .A2(W39914), .ZN(W45296));
  NANDX1 G19644 (.A1(W11769), .A2(I806), .ZN(O14599));
  NANDX1 G19645 (.A1(W30980), .A2(W13037), .ZN(O14597));
  NANDX1 G19646 (.A1(W21023), .A2(W14565), .ZN(O14588));
  NANDX1 G19647 (.A1(W32597), .A2(W39251), .ZN(W45281));
  NANDX1 G19648 (.A1(W12012), .A2(I274), .ZN(O14586));
  NANDX1 G19649 (.A1(W39508), .A2(W30327), .ZN(W45278));
  NANDX1 G19650 (.A1(W34050), .A2(W21999), .ZN(O14484));
  NANDX1 G19651 (.A1(W19741), .A2(W3623), .ZN(O14582));
  NANDX1 G19652 (.A1(W20272), .A2(W35803), .ZN(O14581));
  NANDX1 G19653 (.A1(W34553), .A2(W24983), .ZN(O14575));
  NANDX1 G19654 (.A1(W17541), .A2(W30919), .ZN(W45262));
  NANDX1 G19655 (.A1(W23587), .A2(W42058), .ZN(O14574));
  NANDX1 G19656 (.A1(W31686), .A2(W6985), .ZN(O14570));
  NANDX1 G19657 (.A1(W3510), .A2(W3004), .ZN(W45254));
  NANDX1 G19658 (.A1(W11980), .A2(W29809), .ZN(O14564));
  NANDX1 G19659 (.A1(W11102), .A2(W27230), .ZN(O14562));
  NANDX1 G19660 (.A1(W12946), .A2(W29250), .ZN(O14557));
  NANDX1 G19661 (.A1(W39094), .A2(W16882), .ZN(O14555));
  NANDX1 G19662 (.A1(W25277), .A2(W43516), .ZN(O14413));
  NANDX1 G19663 (.A1(W15931), .A2(W5777), .ZN(O14439));
  NANDX1 G19664 (.A1(W43432), .A2(I1993), .ZN(O14436));
  NANDX1 G19665 (.A1(W1879), .A2(W2197), .ZN(O14433));
  NANDX1 G19666 (.A1(I1104), .A2(W29441), .ZN(O14432));
  NANDX1 G19667 (.A1(W16969), .A2(W16255), .ZN(W45089));
  NANDX1 G19668 (.A1(W21630), .A2(W5130), .ZN(O14430));
  NANDX1 G19669 (.A1(W14573), .A2(W23691), .ZN(O14427));
  NANDX1 G19670 (.A1(W44864), .A2(W7702), .ZN(O14424));
  NANDX1 G19671 (.A1(W29162), .A2(W17549), .ZN(W45078));
  NANDX1 G19672 (.A1(W22161), .A2(W39234), .ZN(O14418));
  NANDX1 G19673 (.A1(W26131), .A2(W39491), .ZN(O14416));
  NANDX1 G19674 (.A1(W30345), .A2(W24424), .ZN(O14415));
  NANDX1 G19675 (.A1(W27613), .A2(W19287), .ZN(W45102));
  NANDX1 G19676 (.A1(W25447), .A2(W35662), .ZN(O14403));
  NANDX1 G19677 (.A1(W14473), .A2(W24094), .ZN(O14401));
  NANDX1 G19678 (.A1(W27418), .A2(W3007), .ZN(W45049));
  NANDX1 G19679 (.A1(W22545), .A2(W22320), .ZN(O14396));
  NANDX1 G19680 (.A1(W13919), .A2(W37257), .ZN(O14395));
  NANDX1 G19681 (.A1(W12311), .A2(W36070), .ZN(O14391));
  NANDX1 G19682 (.A1(W6834), .A2(W14416), .ZN(O14387));
  NANDX1 G19683 (.A1(W40594), .A2(W41747), .ZN(O14376));
  NANDX1 G19684 (.A1(W30540), .A2(W6424), .ZN(O14374));
  NANDX1 G19685 (.A1(W39691), .A2(W34132), .ZN(O14373));
  NANDX1 G19686 (.A1(W39466), .A2(W2276), .ZN(O14370));
  NANDX1 G19687 (.A1(W22899), .A2(W34286), .ZN(O14464));
  NANDX1 G19688 (.A1(W19396), .A2(W35087), .ZN(O14483));
  NANDX1 G19689 (.A1(W9850), .A2(W5973), .ZN(W45149));
  NANDX1 G19690 (.A1(W22277), .A2(W6145), .ZN(O14480));
  NANDX1 G19691 (.A1(W8112), .A2(W17988), .ZN(O14475));
  NANDX1 G19692 (.A1(W20941), .A2(W26726), .ZN(O14474));
  NANDX1 G19693 (.A1(W10235), .A2(W26357), .ZN(W45141));
  NANDX1 G19694 (.A1(W16862), .A2(W1533), .ZN(O14472));
  NANDX1 G19695 (.A1(W3573), .A2(W28544), .ZN(W45135));
  NANDX1 G19696 (.A1(W10904), .A2(I1915), .ZN(O14468));
  NANDX1 G19697 (.A1(W6933), .A2(W31486), .ZN(O14467));
  NANDX1 G19698 (.A1(W31312), .A2(W23372), .ZN(O14466));
  NANDX1 G19699 (.A1(W43982), .A2(W10846), .ZN(O14617));
  NANDX1 G19700 (.A1(W23546), .A2(W38785), .ZN(O14463));
  NANDX1 G19701 (.A1(W37682), .A2(W43694), .ZN(O14462));
  NANDX1 G19702 (.A1(W27897), .A2(W18201), .ZN(W45125));
  NANDX1 G19703 (.A1(W3140), .A2(W25286), .ZN(O14457));
  NANDX1 G19704 (.A1(W6275), .A2(W10026), .ZN(O14455));
  NANDX1 G19705 (.A1(W14062), .A2(W17018), .ZN(W45114));
  NANDX1 G19706 (.A1(W9597), .A2(W42363), .ZN(O14449));
  NANDX1 G19707 (.A1(W15104), .A2(W10555), .ZN(W45108));
  NANDX1 G19708 (.A1(W5392), .A2(W7910), .ZN(O14448));
  NANDX1 G19709 (.A1(W23134), .A2(W31673), .ZN(O14445));
  NANDX1 G19710 (.A1(W6921), .A2(W5768), .ZN(O14444));
  NANDX1 G19711 (.A1(W23746), .A2(W11745), .ZN(O14758));
  NANDX1 G19712 (.A1(W30068), .A2(W40281), .ZN(O14792));
  NANDX1 G19713 (.A1(W17264), .A2(W4601), .ZN(O14790));
  NANDX1 G19714 (.A1(W17764), .A2(W3667), .ZN(O14786));
  NANDX1 G19715 (.A1(I1940), .A2(W32237), .ZN(O14783));
  NANDX1 G19716 (.A1(W18543), .A2(W35691), .ZN(O14781));
  NANDX1 G19717 (.A1(W26295), .A2(W3414), .ZN(O14773));
  NANDX1 G19718 (.A1(I1494), .A2(W37331), .ZN(W45504));
  NANDX1 G19719 (.A1(W18485), .A2(W43831), .ZN(O14771));
  NANDX1 G19720 (.A1(I1536), .A2(W43786), .ZN(O14764));
  NANDX1 G19721 (.A1(W40822), .A2(W13048), .ZN(O14763));
  NANDX1 G19722 (.A1(W1814), .A2(W36975), .ZN(W45490));
  NANDX1 G19723 (.A1(W36974), .A2(W43882), .ZN(W45488));
  NANDX1 G19724 (.A1(W10146), .A2(W9079), .ZN(O14794));
  NANDX1 G19725 (.A1(W25740), .A2(W7726), .ZN(O14756));
  NANDX1 G19726 (.A1(W31104), .A2(W40175), .ZN(O14753));
  NANDX1 G19727 (.A1(W37248), .A2(W24925), .ZN(O14751));
  NANDX1 G19728 (.A1(W24223), .A2(W32280), .ZN(O14745));
  NANDX1 G19729 (.A1(W41698), .A2(W30685), .ZN(O14744));
  NANDX1 G19730 (.A1(W18690), .A2(W16546), .ZN(O14743));
  NANDX1 G19731 (.A1(W8441), .A2(W25379), .ZN(W45469));
  NANDX1 G19732 (.A1(W10254), .A2(W10336), .ZN(W45468));
  NANDX1 G19733 (.A1(W16723), .A2(W37507), .ZN(O14739));
  NANDX1 G19734 (.A1(I583), .A2(W6422), .ZN(O14737));
  NANDX1 G19735 (.A1(W18716), .A2(W30747), .ZN(W45456));
  NANDX1 G19736 (.A1(W1231), .A2(W5448), .ZN(O14832));
  NANDX1 G19737 (.A1(W35961), .A2(W12471), .ZN(O14855));
  NANDX1 G19738 (.A1(W22240), .A2(W3392), .ZN(O14849));
  NANDX1 G19739 (.A1(W7681), .A2(W6494), .ZN(O14846));
  NANDX1 G19740 (.A1(W12972), .A2(W45574), .ZN(O14843));
  NANDX1 G19741 (.A1(W36106), .A2(W11785), .ZN(O14840));
  NANDX1 G19742 (.A1(W76), .A2(W14913), .ZN(W45590));
  NANDX1 G19743 (.A1(W43843), .A2(W32135), .ZN(W45587));
  NANDX1 G19744 (.A1(W23800), .A2(W20665), .ZN(W45585));
  NANDX1 G19745 (.A1(W44132), .A2(W11415), .ZN(O14836));
  NANDX1 G19746 (.A1(W26707), .A2(W25206), .ZN(O14833));
  NANDX1 G19747 (.A1(W31888), .A2(W26849), .ZN(W45580));
  NANDX1 G19748 (.A1(W15092), .A2(W11650), .ZN(O14733));
  NANDX1 G19749 (.A1(W14628), .A2(W6636), .ZN(O14830));
  NANDX1 G19750 (.A1(W23678), .A2(W8756), .ZN(W45571));
  NANDX1 G19751 (.A1(W2276), .A2(W9739), .ZN(O14824));
  NANDX1 G19752 (.A1(W42520), .A2(W34339), .ZN(O14822));
  NANDX1 G19753 (.A1(W32425), .A2(W16877), .ZN(O14810));
  NANDX1 G19754 (.A1(W25052), .A2(W23788), .ZN(O14809));
  NANDX1 G19755 (.A1(W28576), .A2(W33988), .ZN(O14806));
  NANDX1 G19756 (.A1(W40797), .A2(W33301), .ZN(W45543));
  NANDX1 G19757 (.A1(W23628), .A2(W14105), .ZN(O14803));
  NANDX1 G19758 (.A1(W6900), .A2(W40086), .ZN(O14798));
  NANDX1 G19759 (.A1(W9918), .A2(W25804), .ZN(W45529));
  NANDX1 G19760 (.A1(W31977), .A2(W39108), .ZN(O14648));
  NANDX1 G19761 (.A1(W32114), .A2(W4110), .ZN(O14669));
  NANDX1 G19762 (.A1(W12414), .A2(W1489), .ZN(O14668));
  NANDX1 G19763 (.A1(W28066), .A2(W9158), .ZN(O14665));
  NANDX1 G19764 (.A1(I712), .A2(W31572), .ZN(O14664));
  NANDX1 G19765 (.A1(W5228), .A2(W16841), .ZN(W45371));
  NANDX1 G19766 (.A1(W12235), .A2(W17290), .ZN(O14662));
  NANDX1 G19767 (.A1(W32724), .A2(W10849), .ZN(W45365));
  NANDX1 G19768 (.A1(W22171), .A2(W1780), .ZN(W45364));
  NANDX1 G19769 (.A1(W30439), .A2(W30916), .ZN(O14656));
  NANDX1 G19770 (.A1(W22966), .A2(W1807), .ZN(O14655));
  NANDX1 G19771 (.A1(W36274), .A2(W6253), .ZN(O14650));
  NANDX1 G19772 (.A1(W6405), .A2(W23272), .ZN(O14649));
  NANDX1 G19773 (.A1(W16449), .A2(W6041), .ZN(O14671));
  NANDX1 G19774 (.A1(W34747), .A2(W1082), .ZN(O14646));
  NANDX1 G19775 (.A1(W29381), .A2(W7932), .ZN(O14644));
  NANDX1 G19776 (.A1(W27364), .A2(W21567), .ZN(O14642));
  NANDX1 G19777 (.A1(W9082), .A2(W19831), .ZN(O14638));
  NANDX1 G19778 (.A1(W22069), .A2(W6459), .ZN(O14636));
  NANDX1 G19779 (.A1(W37801), .A2(W37798), .ZN(O14635));
  NANDX1 G19780 (.A1(W10633), .A2(W41772), .ZN(O14630));
  NANDX1 G19781 (.A1(W20535), .A2(W7923), .ZN(O14628));
  NANDX1 G19782 (.A1(W20528), .A2(W41186), .ZN(O14627));
  NANDX1 G19783 (.A1(W35624), .A2(W7170), .ZN(O14626));
  NANDX1 G19784 (.A1(W36996), .A2(W41906), .ZN(O14621));
  NANDX1 G19785 (.A1(W21479), .A2(W6092), .ZN(O14704));
  NANDX1 G19786 (.A1(W42499), .A2(W15500), .ZN(O14731));
  NANDX1 G19787 (.A1(W33401), .A2(W36697), .ZN(O14730));
  NANDX1 G19788 (.A1(W23769), .A2(W18137), .ZN(O14725));
  NANDX1 G19789 (.A1(W884), .A2(W43898), .ZN(O14723));
  NANDX1 G19790 (.A1(W18858), .A2(W17529), .ZN(O14720));
  NANDX1 G19791 (.A1(W35352), .A2(W32794), .ZN(O14719));
  NANDX1 G19792 (.A1(W7828), .A2(W7963), .ZN(W45437));
  NANDX1 G19793 (.A1(W29473), .A2(W27406), .ZN(O14716));
  NANDX1 G19794 (.A1(W28699), .A2(W43819), .ZN(O14715));
  NANDX1 G19795 (.A1(W32459), .A2(W11441), .ZN(O14714));
  NANDX1 G19796 (.A1(W28700), .A2(W6807), .ZN(O14706));
  NANDX1 G19797 (.A1(W6809), .A2(W16756), .ZN(O13393));
  NANDX1 G19798 (.A1(W33437), .A2(W450), .ZN(O14698));
  NANDX1 G19799 (.A1(W14894), .A2(W12882), .ZN(W45409));
  NANDX1 G19800 (.A1(W7169), .A2(W19397), .ZN(O14689));
  NANDX1 G19801 (.A1(W32806), .A2(W42171), .ZN(O14685));
  NANDX1 G19802 (.A1(W9237), .A2(W37441), .ZN(O14684));
  NANDX1 G19803 (.A1(W43135), .A2(W7321), .ZN(O14683));
  NANDX1 G19804 (.A1(W8919), .A2(W1336), .ZN(O14680));
  NANDX1 G19805 (.A1(W32934), .A2(W2817), .ZN(W45387));
  NANDX1 G19806 (.A1(W11244), .A2(W17753), .ZN(O14674));
  NANDX1 G19807 (.A1(W16249), .A2(W8027), .ZN(W45383));
  NANDX1 G19808 (.A1(W4249), .A2(W5827), .ZN(O14672));
  NANDX1 G19809 (.A1(W21332), .A2(W21242), .ZN(O12200));
  NANDX1 G19810 (.A1(W7816), .A2(W20402), .ZN(O12225));
  NANDX1 G19811 (.A1(W29984), .A2(W12793), .ZN(O12224));
  NANDX1 G19812 (.A1(W816), .A2(W1799), .ZN(O12222));
  NANDX1 G19813 (.A1(W7555), .A2(W40752), .ZN(O12221));
  NANDX1 G19814 (.A1(W31715), .A2(W27274), .ZN(O12218));
  NANDX1 G19815 (.A1(W35800), .A2(W11073), .ZN(O12216));
  NANDX1 G19816 (.A1(W31890), .A2(W31550), .ZN(W42259));
  NANDX1 G19817 (.A1(W25587), .A2(W41397), .ZN(O12208));
  NANDX1 G19818 (.A1(W27627), .A2(W32290), .ZN(O12206));
  NANDX1 G19819 (.A1(W1333), .A2(W19061), .ZN(W42254));
  NANDX1 G19820 (.A1(W17976), .A2(W23241), .ZN(O12205));
  NANDX1 G19821 (.A1(W0), .A2(W40031), .ZN(O12204));
  NANDX1 G19822 (.A1(W11113), .A2(W2989), .ZN(O12226));
  NANDX1 G19823 (.A1(W37312), .A2(W35781), .ZN(O12199));
  NANDX1 G19824 (.A1(W2962), .A2(W3023), .ZN(W42242));
  NANDX1 G19825 (.A1(W7350), .A2(W27563), .ZN(W42239));
  NANDX1 G19826 (.A1(W29577), .A2(W13135), .ZN(W42236));
  NANDX1 G19827 (.A1(W5615), .A2(W4245), .ZN(W42233));
  NANDX1 G19828 (.A1(W4399), .A2(W35182), .ZN(O12190));
  NANDX1 G19829 (.A1(W5307), .A2(W5819), .ZN(O12189));
  NANDX1 G19830 (.A1(W9105), .A2(W22151), .ZN(W42228));
  NANDX1 G19831 (.A1(W28115), .A2(W35198), .ZN(O12188));
  NANDX1 G19832 (.A1(W30375), .A2(W37423), .ZN(O12187));
  NANDX1 G19833 (.A1(W12450), .A2(W38091), .ZN(O12185));
  NANDX1 G19834 (.A1(W33752), .A2(W22832), .ZN(W42307));
  NANDX1 G19835 (.A1(W59), .A2(W11723), .ZN(O12277));
  NANDX1 G19836 (.A1(W29346), .A2(W35664), .ZN(W42345));
  NANDX1 G19837 (.A1(W9455), .A2(W31846), .ZN(O12274));
  NANDX1 G19838 (.A1(W18731), .A2(W7804), .ZN(O12272));
  NANDX1 G19839 (.A1(W34797), .A2(W41842), .ZN(O12269));
  NANDX1 G19840 (.A1(W27153), .A2(W1589), .ZN(O12268));
  NANDX1 G19841 (.A1(W1938), .A2(I1171), .ZN(O12266));
  NANDX1 G19842 (.A1(W31372), .A2(W228), .ZN(O12260));
  NANDX1 G19843 (.A1(W35804), .A2(W33966), .ZN(O12259));
  NANDX1 G19844 (.A1(W18286), .A2(W37541), .ZN(W42317));
  NANDX1 G19845 (.A1(W25596), .A2(W17190), .ZN(O12250));
  NANDX1 G19846 (.A1(W27737), .A2(W38958), .ZN(O12246));
  NANDX1 G19847 (.A1(W32285), .A2(W34330), .ZN(O12183));
  NANDX1 G19848 (.A1(I1988), .A2(W5960), .ZN(W42306));
  NANDX1 G19849 (.A1(W3081), .A2(W27371), .ZN(W42302));
  NANDX1 G19850 (.A1(W6173), .A2(W13982), .ZN(O12243));
  NANDX1 G19851 (.A1(W25000), .A2(W21724), .ZN(W42300));
  NANDX1 G19852 (.A1(W16906), .A2(W12012), .ZN(O12241));
  NANDX1 G19853 (.A1(W32723), .A2(W20459), .ZN(W42296));
  NANDX1 G19854 (.A1(W3356), .A2(W15396), .ZN(O12240));
  NANDX1 G19855 (.A1(W18371), .A2(W22354), .ZN(O12234));
  NANDX1 G19856 (.A1(W12393), .A2(W38601), .ZN(W42288));
  NANDX1 G19857 (.A1(W30952), .A2(W16584), .ZN(O12231));
  NANDX1 G19858 (.A1(W16114), .A2(W32751), .ZN(O12228));
  NANDX1 G19859 (.A1(W401), .A2(W23932), .ZN(O12107));
  NANDX1 G19860 (.A1(W31894), .A2(W5991), .ZN(O12123));
  NANDX1 G19861 (.A1(W1953), .A2(W39688), .ZN(O12122));
  NANDX1 G19862 (.A1(W28913), .A2(W24041), .ZN(W42139));
  NANDX1 G19863 (.A1(W31423), .A2(W4956), .ZN(O12121));
  NANDX1 G19864 (.A1(W28726), .A2(W12588), .ZN(O12119));
  NANDX1 G19865 (.A1(W16272), .A2(W30194), .ZN(O12116));
  NANDX1 G19866 (.A1(W8655), .A2(W5924), .ZN(O12115));
  NANDX1 G19867 (.A1(W33503), .A2(W3851), .ZN(O12113));
  NANDX1 G19868 (.A1(W24872), .A2(W2548), .ZN(O12112));
  NANDX1 G19869 (.A1(W40009), .A2(W6078), .ZN(O12110));
  NANDX1 G19870 (.A1(I943), .A2(W23451), .ZN(O12109));
  NANDX1 G19871 (.A1(W33635), .A2(W8514), .ZN(O12108));
  NANDX1 G19872 (.A1(W30336), .A2(W9749), .ZN(O12124));
  NANDX1 G19873 (.A1(W6612), .A2(W6342), .ZN(O12105));
  NANDX1 G19874 (.A1(W12873), .A2(W14199), .ZN(O12104));
  NANDX1 G19875 (.A1(W22493), .A2(W9319), .ZN(O12102));
  NANDX1 G19876 (.A1(W40156), .A2(W21774), .ZN(O12100));
  NANDX1 G19877 (.A1(W6239), .A2(W30503), .ZN(O12099));
  NANDX1 G19878 (.A1(W22583), .A2(W20430), .ZN(W42108));
  NANDX1 G19879 (.A1(W40514), .A2(I732), .ZN(O12094));
  NANDX1 G19880 (.A1(W38907), .A2(W24122), .ZN(W42104));
  NANDX1 G19881 (.A1(W38329), .A2(W30961), .ZN(O12088));
  NANDX1 G19882 (.A1(W32368), .A2(W16357), .ZN(O12087));
  NANDX1 G19883 (.A1(W19974), .A2(W28366), .ZN(O12084));
  NANDX1 G19884 (.A1(W22066), .A2(W31661), .ZN(O12154));
  NANDX1 G19885 (.A1(W12456), .A2(W39480), .ZN(W42220));
  NANDX1 G19886 (.A1(W19399), .A2(W26482), .ZN(W42218));
  NANDX1 G19887 (.A1(W25561), .A2(W37441), .ZN(O12171));
  NANDX1 G19888 (.A1(W1763), .A2(W40348), .ZN(W42203));
  NANDX1 G19889 (.A1(W5129), .A2(W8590), .ZN(O12168));
  NANDX1 G19890 (.A1(W26422), .A2(W8043), .ZN(O12166));
  NANDX1 G19891 (.A1(W17109), .A2(W22177), .ZN(O12165));
  NANDX1 G19892 (.A1(W29358), .A2(W34531), .ZN(O12162));
  NANDX1 G19893 (.A1(W33148), .A2(W17430), .ZN(O12160));
  NANDX1 G19894 (.A1(W32083), .A2(W24066), .ZN(O12159));
  NANDX1 G19895 (.A1(W30381), .A2(W41601), .ZN(O12157));
  NANDX1 G19896 (.A1(W34957), .A2(W3400), .ZN(O12278));
  NANDX1 G19897 (.A1(W26306), .A2(W6821), .ZN(O12152));
  NANDX1 G19898 (.A1(W23907), .A2(W9223), .ZN(O12148));
  NANDX1 G19899 (.A1(W36361), .A2(W10306), .ZN(W42175));
  NANDX1 G19900 (.A1(W35142), .A2(W7672), .ZN(W42172));
  NANDX1 G19901 (.A1(W35375), .A2(I975), .ZN(W42171));
  NANDX1 G19902 (.A1(W29181), .A2(W31106), .ZN(W42164));
  NANDX1 G19903 (.A1(W19998), .A2(W3328), .ZN(O12135));
  NANDX1 G19904 (.A1(W27016), .A2(W26267), .ZN(O12134));
  NANDX1 G19905 (.A1(W30705), .A2(I361), .ZN(O12133));
  NANDX1 G19906 (.A1(W8065), .A2(W11962), .ZN(O12132));
  NANDX1 G19907 (.A1(W25055), .A2(W27004), .ZN(O12131));
  NANDX1 G19908 (.A1(W28574), .A2(W36941), .ZN(O12447));
  NANDX1 G19909 (.A1(W4818), .A2(W1126), .ZN(O12478));
  NANDX1 G19910 (.A1(W16856), .A2(W338), .ZN(O12472));
  NANDX1 G19911 (.A1(W42362), .A2(W11112), .ZN(O12470));
  NANDX1 G19912 (.A1(W32078), .A2(W13747), .ZN(O12469));
  NANDX1 G19913 (.A1(W33100), .A2(W17305), .ZN(O12468));
  NANDX1 G19914 (.A1(W37462), .A2(W27319), .ZN(O12467));
  NANDX1 G19915 (.A1(W6566), .A2(W30561), .ZN(O12464));
  NANDX1 G19916 (.A1(W37107), .A2(W4263), .ZN(O12460));
  NANDX1 G19917 (.A1(W29596), .A2(W4200), .ZN(O12459));
  NANDX1 G19918 (.A1(W2441), .A2(W6151), .ZN(W42578));
  NANDX1 G19919 (.A1(W37414), .A2(W24536), .ZN(W42573));
  NANDX1 G19920 (.A1(W5315), .A2(W6238), .ZN(O12449));
  NANDX1 G19921 (.A1(W25182), .A2(W30642), .ZN(O12482));
  NANDX1 G19922 (.A1(W8570), .A2(W13971), .ZN(O12444));
  NANDX1 G19923 (.A1(W16784), .A2(W8911), .ZN(O12437));
  NANDX1 G19924 (.A1(W21077), .A2(W7520), .ZN(O12436));
  NANDX1 G19925 (.A1(W16048), .A2(W22768), .ZN(O12434));
  NANDX1 G19926 (.A1(W24554), .A2(W6372), .ZN(O12432));
  NANDX1 G19927 (.A1(W3777), .A2(W11897), .ZN(O12428));
  NANDX1 G19928 (.A1(W21377), .A2(W37796), .ZN(O12424));
  NANDX1 G19929 (.A1(W22580), .A2(W36378), .ZN(O12423));
  NANDX1 G19930 (.A1(W21018), .A2(W40510), .ZN(W42541));
  NANDX1 G19931 (.A1(W34504), .A2(W1849), .ZN(O12421));
  NANDX1 G19932 (.A1(W39625), .A2(W36263), .ZN(O12420));
  NANDX1 G19933 (.A1(W41905), .A2(W5137), .ZN(O12504));
  NANDX1 G19934 (.A1(W1355), .A2(I1361), .ZN(O12532));
  NANDX1 G19935 (.A1(W13475), .A2(W39946), .ZN(O12531));
  NANDX1 G19936 (.A1(W11528), .A2(W36229), .ZN(O12529));
  NANDX1 G19937 (.A1(W5206), .A2(W158), .ZN(O12526));
  NANDX1 G19938 (.A1(W28129), .A2(W28103), .ZN(O12525));
  NANDX1 G19939 (.A1(W26012), .A2(W33191), .ZN(O12523));
  NANDX1 G19940 (.A1(W41170), .A2(W7018), .ZN(O12522));
  NANDX1 G19941 (.A1(W1100), .A2(W2773), .ZN(O12517));
  NANDX1 G19942 (.A1(W27360), .A2(W20387), .ZN(W42660));
  NANDX1 G19943 (.A1(W617), .A2(W17047), .ZN(O12511));
  NANDX1 G19944 (.A1(W23568), .A2(W16398), .ZN(W42653));
  NANDX1 G19945 (.A1(W26408), .A2(W9368), .ZN(O12505));
  NANDX1 G19946 (.A1(W36147), .A2(W8633), .ZN(O12413));
  NANDX1 G19947 (.A1(W3379), .A2(W39768), .ZN(O12503));
  NANDX1 G19948 (.A1(W419), .A2(W27105), .ZN(O12502));
  NANDX1 G19949 (.A1(W21608), .A2(W6693), .ZN(O12501));
  NANDX1 G19950 (.A1(W14989), .A2(W34674), .ZN(O12500));
  NANDX1 G19951 (.A1(W10646), .A2(W39031), .ZN(W42640));
  NANDX1 G19952 (.A1(W37183), .A2(W24978), .ZN(O12495));
  NANDX1 G19953 (.A1(W17091), .A2(W31408), .ZN(O12494));
  NANDX1 G19954 (.A1(W8237), .A2(W40886), .ZN(O12492));
  NANDX1 G19955 (.A1(W10936), .A2(W37975), .ZN(W42630));
  NANDX1 G19956 (.A1(W23106), .A2(W14269), .ZN(O12491));
  NANDX1 G19957 (.A1(W34106), .A2(W4716), .ZN(O12488));
  NANDX1 G19958 (.A1(W19946), .A2(W3457), .ZN(W42380));
  NANDX1 G19959 (.A1(W23671), .A2(W41945), .ZN(O12336));
  NANDX1 G19960 (.A1(W27308), .A2(W5524), .ZN(O12332));
  NANDX1 G19961 (.A1(I1569), .A2(I1575), .ZN(O12327));
  NANDX1 G19962 (.A1(W26760), .A2(W28428), .ZN(O12325));
  NANDX1 G19963 (.A1(W7058), .A2(W35591), .ZN(W42414));
  NANDX1 G19964 (.A1(W9940), .A2(W13646), .ZN(O12323));
  NANDX1 G19965 (.A1(W7819), .A2(W7733), .ZN(O12321));
  NANDX1 G19966 (.A1(W34852), .A2(W15760), .ZN(O12315));
  NANDX1 G19967 (.A1(W8966), .A2(W32832), .ZN(O12304));
  NANDX1 G19968 (.A1(W9192), .A2(W22159), .ZN(O12299));
  NANDX1 G19969 (.A1(W7973), .A2(W28941), .ZN(O12298));
  NANDX1 G19970 (.A1(W15915), .A2(W15569), .ZN(W42382));
  NANDX1 G19971 (.A1(W42064), .A2(W7978), .ZN(O12341));
  NANDX1 G19972 (.A1(W18800), .A2(W35456), .ZN(O12293));
  NANDX1 G19973 (.A1(W38089), .A2(W27504), .ZN(O12292));
  NANDX1 G19974 (.A1(W41040), .A2(W37821), .ZN(O12291));
  NANDX1 G19975 (.A1(W20301), .A2(W4456), .ZN(O12289));
  NANDX1 G19976 (.A1(W25642), .A2(W26635), .ZN(O12286));
  NANDX1 G19977 (.A1(W36501), .A2(W4268), .ZN(W42361));
  NANDX1 G19978 (.A1(W33551), .A2(W13217), .ZN(W42360));
  NANDX1 G19979 (.A1(W27753), .A2(W14893), .ZN(W42358));
  NANDX1 G19980 (.A1(W979), .A2(W41998), .ZN(O12281));
  NANDX1 G19981 (.A1(W29832), .A2(W31394), .ZN(W42352));
  NANDX1 G19982 (.A1(W16291), .A2(W25862), .ZN(W42351));
  NANDX1 G19983 (.A1(W4678), .A2(W12841), .ZN(O12374));
  NANDX1 G19984 (.A1(W25702), .A2(W29419), .ZN(O12412));
  NANDX1 G19985 (.A1(W27065), .A2(W6370), .ZN(O12409));
  NANDX1 G19986 (.A1(W38631), .A2(W10395), .ZN(W42520));
  NANDX1 G19987 (.A1(W22443), .A2(W27544), .ZN(W42515));
  NANDX1 G19988 (.A1(W34552), .A2(W12327), .ZN(O12404));
  NANDX1 G19989 (.A1(W28601), .A2(W33242), .ZN(O12403));
  NANDX1 G19990 (.A1(W28284), .A2(W33752), .ZN(O12402));
  NANDX1 G19991 (.A1(W13509), .A2(W29628), .ZN(O12391));
  NANDX1 G19992 (.A1(W12946), .A2(W31659), .ZN(O12385));
  NANDX1 G19993 (.A1(W7585), .A2(W5356), .ZN(W42490));
  NANDX1 G19994 (.A1(W36749), .A2(W3010), .ZN(O12382));
  NANDX1 G19995 (.A1(W21919), .A2(W10699), .ZN(O12083));
  NANDX1 G19996 (.A1(W6086), .A2(W35823), .ZN(W42477));
  NANDX1 G19997 (.A1(W21212), .A2(W292), .ZN(O12362));
  NANDX1 G19998 (.A1(W14915), .A2(W5584), .ZN(O12361));
  NANDX1 G19999 (.A1(W14775), .A2(W27297), .ZN(O12355));
  NANDX1 G20000 (.A1(W32131), .A2(W22689), .ZN(O12352));
  NANDX1 G20001 (.A1(W18452), .A2(W19823), .ZN(W42450));
  NANDX1 G20002 (.A1(W7998), .A2(W11556), .ZN(O12348));
  NANDX1 G20003 (.A1(W25771), .A2(W19078), .ZN(O12345));
  NANDX1 G20004 (.A1(W482), .A2(W5792), .ZN(O12343));
  NANDX1 G20005 (.A1(W3328), .A2(W18077), .ZN(O12342));
  NANDX1 G20006 (.A1(W15111), .A2(W18480), .ZN(W42439));
  NANDX1 G20007 (.A1(W16977), .A2(I1115), .ZN(O11783));
  NANDX1 G20008 (.A1(W1495), .A2(W26719), .ZN(O11813));
  NANDX1 G20009 (.A1(W22434), .A2(W667), .ZN(O11809));
  NANDX1 G20010 (.A1(W18966), .A2(W32967), .ZN(W41720));
  NANDX1 G20011 (.A1(W7686), .A2(W6729), .ZN(W41718));
  NANDX1 G20012 (.A1(W25449), .A2(W25199), .ZN(O11801));
  NANDX1 G20013 (.A1(W26236), .A2(W34949), .ZN(W41712));
  NANDX1 G20014 (.A1(W32661), .A2(W21980), .ZN(O11799));
  NANDX1 G20015 (.A1(W6924), .A2(W26621), .ZN(W41704));
  NANDX1 G20016 (.A1(W19066), .A2(W6823), .ZN(O11793));
  NANDX1 G20017 (.A1(W40310), .A2(W20966), .ZN(O11792));
  NANDX1 G20018 (.A1(W30155), .A2(I1534), .ZN(W41699));
  NANDX1 G20019 (.A1(W35386), .A2(W8588), .ZN(W41690));
  NANDX1 G20020 (.A1(W30773), .A2(W8678), .ZN(O11815));
  NANDX1 G20021 (.A1(W13819), .A2(W28692), .ZN(W41680));
  NANDX1 G20022 (.A1(W8932), .A2(W37680), .ZN(O11778));
  NANDX1 G20023 (.A1(W40568), .A2(W23724), .ZN(W41678));
  NANDX1 G20024 (.A1(W16395), .A2(W16928), .ZN(O11776));
  NANDX1 G20025 (.A1(W40532), .A2(W35659), .ZN(W41675));
  NANDX1 G20026 (.A1(W39369), .A2(W35381), .ZN(O11774));
  NANDX1 G20027 (.A1(W11333), .A2(W12171), .ZN(W41671));
  NANDX1 G20028 (.A1(W21024), .A2(W20611), .ZN(W41670));
  NANDX1 G20029 (.A1(W21357), .A2(W33536), .ZN(W41666));
  NANDX1 G20030 (.A1(W2280), .A2(W36518), .ZN(W41664));
  NANDX1 G20031 (.A1(W6133), .A2(W39684), .ZN(O11769));
  NANDX1 G20032 (.A1(W30097), .A2(W17617), .ZN(O11828));
  NANDX1 G20033 (.A1(W30054), .A2(W37472), .ZN(O11857));
  NANDX1 G20034 (.A1(W23996), .A2(W37293), .ZN(O11856));
  NANDX1 G20035 (.A1(W21792), .A2(W19910), .ZN(W41778));
  NANDX1 G20036 (.A1(W34833), .A2(W31182), .ZN(O11847));
  NANDX1 G20037 (.A1(W27277), .A2(W13136), .ZN(W41775));
  NANDX1 G20038 (.A1(W20635), .A2(W38011), .ZN(W41774));
  NANDX1 G20039 (.A1(W38993), .A2(W1535), .ZN(O11842));
  NANDX1 G20040 (.A1(W39936), .A2(W38814), .ZN(W41763));
  NANDX1 G20041 (.A1(W31934), .A2(W7836), .ZN(W41762));
  NANDX1 G20042 (.A1(W12119), .A2(W1361), .ZN(O11835));
  NANDX1 G20043 (.A1(W26461), .A2(W17754), .ZN(W41757));
  NANDX1 G20044 (.A1(W31938), .A2(W12559), .ZN(W41754));
  NANDX1 G20045 (.A1(W33063), .A2(W832), .ZN(W41661));
  NANDX1 G20046 (.A1(W33357), .A2(W22253), .ZN(O11827));
  NANDX1 G20047 (.A1(W40147), .A2(W4014), .ZN(O11826));
  NANDX1 G20048 (.A1(W37998), .A2(W29194), .ZN(W41744));
  NANDX1 G20049 (.A1(W20501), .A2(W1981), .ZN(O11824));
  NANDX1 G20050 (.A1(W23332), .A2(W30), .ZN(O11823));
  NANDX1 G20051 (.A1(W40704), .A2(W17913), .ZN(O11822));
  NANDX1 G20052 (.A1(W14309), .A2(W27954), .ZN(O11821));
  NANDX1 G20053 (.A1(W41391), .A2(W29011), .ZN(O11817));
  NANDX1 G20054 (.A1(W40243), .A2(W33558), .ZN(W41734));
  NANDX1 G20055 (.A1(W37263), .A2(W18660), .ZN(O11816));
  NANDX1 G20056 (.A1(W16814), .A2(W33225), .ZN(W41732));
  NANDX1 G20057 (.A1(W39103), .A2(W38707), .ZN(O11703));
  NANDX1 G20058 (.A1(W13409), .A2(W466), .ZN(O11718));
  NANDX1 G20059 (.A1(W18401), .A2(W41478), .ZN(O11716));
  NANDX1 G20060 (.A1(W27732), .A2(W32299), .ZN(W41589));
  NANDX1 G20061 (.A1(W4155), .A2(W27632), .ZN(O11712));
  NANDX1 G20062 (.A1(W40180), .A2(W17809), .ZN(W41587));
  NANDX1 G20063 (.A1(W19466), .A2(W17040), .ZN(O11708));
  NANDX1 G20064 (.A1(W40680), .A2(W20235), .ZN(W41582));
  NANDX1 G20065 (.A1(W40142), .A2(W41201), .ZN(O11707));
  NANDX1 G20066 (.A1(I707), .A2(W31959), .ZN(O11706));
  NANDX1 G20067 (.A1(W28479), .A2(W14259), .ZN(O11705));
  NANDX1 G20068 (.A1(W34236), .A2(W25777), .ZN(W41577));
  NANDX1 G20069 (.A1(W7179), .A2(W11772), .ZN(W41576));
  NANDX1 G20070 (.A1(W6054), .A2(W34311), .ZN(O11719));
  NANDX1 G20071 (.A1(W25466), .A2(W20055), .ZN(O11702));
  NANDX1 G20072 (.A1(W21414), .A2(W1727), .ZN(O11700));
  NANDX1 G20073 (.A1(W5409), .A2(W28487), .ZN(O11697));
  NANDX1 G20074 (.A1(W34360), .A2(I148), .ZN(O11696));
  NANDX1 G20075 (.A1(W2685), .A2(W33681), .ZN(O11690));
  NANDX1 G20076 (.A1(W7057), .A2(W9898), .ZN(O11687));
  NANDX1 G20077 (.A1(I694), .A2(W13491), .ZN(O11683));
  NANDX1 G20078 (.A1(W442), .A2(W37651), .ZN(O11681));
  NANDX1 G20079 (.A1(W7996), .A2(W3960), .ZN(O11679));
  NANDX1 G20080 (.A1(W28664), .A2(W12535), .ZN(W41543));
  NANDX1 G20081 (.A1(W35092), .A2(W9318), .ZN(O11671));
  NANDX1 G20082 (.A1(I217), .A2(W40067), .ZN(O11749));
  NANDX1 G20083 (.A1(W25208), .A2(I1014), .ZN(O11767));
  NANDX1 G20084 (.A1(W35672), .A2(W34976), .ZN(O11766));
  NANDX1 G20085 (.A1(W17822), .A2(W1118), .ZN(W41656));
  NANDX1 G20086 (.A1(W40338), .A2(W37476), .ZN(O11764));
  NANDX1 G20087 (.A1(W25769), .A2(W8674), .ZN(W41650));
  NANDX1 G20088 (.A1(W27275), .A2(W41282), .ZN(O11760));
  NANDX1 G20089 (.A1(W8390), .A2(W20289), .ZN(W41648));
  NANDX1 G20090 (.A1(W36146), .A2(W9036), .ZN(O11759));
  NANDX1 G20091 (.A1(W10295), .A2(W34762), .ZN(O11757));
  NANDX1 G20092 (.A1(W13050), .A2(W3806), .ZN(O11755));
  NANDX1 G20093 (.A1(W24960), .A2(W8173), .ZN(O11752));
  NANDX1 G20094 (.A1(W41284), .A2(W21569), .ZN(O11866));
  NANDX1 G20095 (.A1(W39922), .A2(W18512), .ZN(O11748));
  NANDX1 G20096 (.A1(W21325), .A2(W18671), .ZN(O11744));
  NANDX1 G20097 (.A1(W2237), .A2(W11118), .ZN(O11743));
  NANDX1 G20098 (.A1(I1749), .A2(W38378), .ZN(O11741));
  NANDX1 G20099 (.A1(W40526), .A2(I412), .ZN(O11740));
  NANDX1 G20100 (.A1(W33035), .A2(W22247), .ZN(O11734));
  NANDX1 G20101 (.A1(W34310), .A2(W5522), .ZN(O11731));
  NANDX1 G20102 (.A1(W6532), .A2(W27216), .ZN(W41609));
  NANDX1 G20103 (.A1(W19435), .A2(W22456), .ZN(W41607));
  NANDX1 G20104 (.A1(W26499), .A2(W35176), .ZN(O11723));
  NANDX1 G20105 (.A1(W8732), .A2(W37124), .ZN(O11721));
  NANDX1 G20106 (.A1(W13924), .A2(W33289), .ZN(W41973));
  NANDX1 G20107 (.A1(W35276), .A2(W12757), .ZN(O12008));
  NANDX1 G20108 (.A1(W40995), .A2(W27288), .ZN(W41994));
  NANDX1 G20109 (.A1(W10300), .A2(W23309), .ZN(W41992));
  NANDX1 G20110 (.A1(W11501), .A2(W34850), .ZN(O12005));
  NANDX1 G20111 (.A1(W28944), .A2(W34370), .ZN(O12004));
  NANDX1 G20112 (.A1(W13942), .A2(W24534), .ZN(O12003));
  NANDX1 G20113 (.A1(W34461), .A2(W20307), .ZN(O12002));
  NANDX1 G20114 (.A1(W31027), .A2(W6010), .ZN(O12000));
  NANDX1 G20115 (.A1(W11623), .A2(I1808), .ZN(W41981));
  NANDX1 G20116 (.A1(W7685), .A2(W20118), .ZN(W41978));
  NANDX1 G20117 (.A1(W4458), .A2(W15294), .ZN(O11996));
  NANDX1 G20118 (.A1(W16746), .A2(W34757), .ZN(W41974));
  NANDX1 G20119 (.A1(W4683), .A2(W39699), .ZN(W41997));
  NANDX1 G20120 (.A1(W14298), .A2(W38187), .ZN(O11994));
  NANDX1 G20121 (.A1(W7700), .A2(W29902), .ZN(O11990));
  NANDX1 G20122 (.A1(W16106), .A2(W15511), .ZN(O11987));
  NANDX1 G20123 (.A1(W41645), .A2(W8714), .ZN(O11986));
  NANDX1 G20124 (.A1(W8852), .A2(W30317), .ZN(O11984));
  NANDX1 G20125 (.A1(W17674), .A2(W33440), .ZN(O11983));
  NANDX1 G20126 (.A1(W14411), .A2(W29982), .ZN(O11980));
  NANDX1 G20127 (.A1(W8776), .A2(W17080), .ZN(O11979));
  NANDX1 G20128 (.A1(W9370), .A2(W29084), .ZN(W41955));
  NANDX1 G20129 (.A1(W14836), .A2(W30274), .ZN(O11978));
  NANDX1 G20130 (.A1(W17909), .A2(W7935), .ZN(O11977));
  NANDX1 G20131 (.A1(I1390), .A2(W32769), .ZN(O12044));
  NANDX1 G20132 (.A1(W11134), .A2(W27797), .ZN(O12080));
  NANDX1 G20133 (.A1(W6045), .A2(W20020), .ZN(O12072));
  NANDX1 G20134 (.A1(W24725), .A2(W13171), .ZN(O12071));
  NANDX1 G20135 (.A1(W8276), .A2(W22483), .ZN(O12069));
  NANDX1 G20136 (.A1(W16004), .A2(W23997), .ZN(O12068));
  NANDX1 G20137 (.A1(W37279), .A2(W36445), .ZN(O12067));
  NANDX1 G20138 (.A1(W25602), .A2(W4113), .ZN(W42064));
  NANDX1 G20139 (.A1(W41450), .A2(W31314), .ZN(O12056));
  NANDX1 G20140 (.A1(W20741), .A2(W13304), .ZN(O12053));
  NANDX1 G20141 (.A1(W26436), .A2(W13059), .ZN(W42049));
  NANDX1 G20142 (.A1(W4), .A2(W22493), .ZN(O12049));
  NANDX1 G20143 (.A1(W13405), .A2(W3051), .ZN(O12047));
  NANDX1 G20144 (.A1(W16403), .A2(W29714), .ZN(O11974));
  NANDX1 G20145 (.A1(W37408), .A2(W18192), .ZN(O12042));
  NANDX1 G20146 (.A1(W8615), .A2(W6655), .ZN(O12041));
  NANDX1 G20147 (.A1(I471), .A2(W30943), .ZN(O12038));
  NANDX1 G20148 (.A1(W29063), .A2(W14749), .ZN(W42033));
  NANDX1 G20149 (.A1(W25763), .A2(W2224), .ZN(W42030));
  NANDX1 G20150 (.A1(W40324), .A2(W38995), .ZN(W42029));
  NANDX1 G20151 (.A1(W22191), .A2(W32817), .ZN(O12027));
  NANDX1 G20152 (.A1(W31817), .A2(W5147), .ZN(O12020));
  NANDX1 G20153 (.A1(W801), .A2(W9638), .ZN(O12019));
  NANDX1 G20154 (.A1(W13540), .A2(W40412), .ZN(O12013));
  NANDX1 G20155 (.A1(I1445), .A2(W32372), .ZN(O12010));
  NANDX1 G20156 (.A1(W27428), .A2(W31755), .ZN(O11890));
  NANDX1 G20157 (.A1(W28993), .A2(W26593), .ZN(O11918));
  NANDX1 G20158 (.A1(W16816), .A2(W35249), .ZN(W41877));
  NANDX1 G20159 (.A1(W34309), .A2(W37929), .ZN(O11915));
  NANDX1 G20160 (.A1(W22867), .A2(W34430), .ZN(O11914));
  NANDX1 G20161 (.A1(W15818), .A2(W36758), .ZN(O11913));
  NANDX1 G20162 (.A1(W19036), .A2(W17786), .ZN(O11909));
  NANDX1 G20163 (.A1(W35711), .A2(W6625), .ZN(O11908));
  NANDX1 G20164 (.A1(W8738), .A2(W37542), .ZN(O11906));
  NANDX1 G20165 (.A1(W12698), .A2(W6141), .ZN(O11904));
  NANDX1 G20166 (.A1(W37364), .A2(W33304), .ZN(O11896));
  NANDX1 G20167 (.A1(W28591), .A2(W36745), .ZN(O11894));
  NANDX1 G20168 (.A1(W2722), .A2(W27744), .ZN(W41842));
  NANDX1 G20169 (.A1(W40938), .A2(W19709), .ZN(W41880));
  NANDX1 G20170 (.A1(W27763), .A2(I1172), .ZN(O11883));
  NANDX1 G20171 (.A1(W26661), .A2(W15018), .ZN(O11882));
  NANDX1 G20172 (.A1(W15006), .A2(W17587), .ZN(W41829));
  NANDX1 G20173 (.A1(W6755), .A2(W39059), .ZN(W41825));
  NANDX1 G20174 (.A1(W41383), .A2(W34033), .ZN(O11879));
  NANDX1 G20175 (.A1(W5542), .A2(W9100), .ZN(W41819));
  NANDX1 G20176 (.A1(W25906), .A2(W31668), .ZN(O11877));
  NANDX1 G20177 (.A1(W11281), .A2(W145), .ZN(O11873));
  NANDX1 G20178 (.A1(W26614), .A2(W38417), .ZN(O11872));
  NANDX1 G20179 (.A1(W16553), .A2(W26706), .ZN(O11867));
  NANDX1 G20180 (.A1(W30567), .A2(W36474), .ZN(W41805));
  NANDX1 G20181 (.A1(W5008), .A2(W28071), .ZN(O11956));
  NANDX1 G20182 (.A1(W26751), .A2(W39599), .ZN(O11973));
  NANDX1 G20183 (.A1(W1505), .A2(W27238), .ZN(O11970));
  NANDX1 G20184 (.A1(W797), .A2(W18797), .ZN(W41945));
  NANDX1 G20185 (.A1(W12990), .A2(W19136), .ZN(O11969));
  NANDX1 G20186 (.A1(W11251), .A2(W27023), .ZN(O11967));
  NANDX1 G20187 (.A1(W31819), .A2(W2411), .ZN(W41939));
  NANDX1 G20188 (.A1(W24093), .A2(W36279), .ZN(O11965));
  NANDX1 G20189 (.A1(W36143), .A2(W25769), .ZN(O11963));
  NANDX1 G20190 (.A1(W18985), .A2(W1642), .ZN(O11961));
  NANDX1 G20191 (.A1(W8748), .A2(W20603), .ZN(W41930));
  NANDX1 G20192 (.A1(W8997), .A2(W16185), .ZN(O11957));
  NANDX1 G20193 (.A1(W38870), .A2(W30263), .ZN(O12533));
  NANDX1 G20194 (.A1(W13499), .A2(W4709), .ZN(O11949));
  NANDX1 G20195 (.A1(W9266), .A2(W5647), .ZN(O11948));
  NANDX1 G20196 (.A1(W8387), .A2(W34248), .ZN(O11946));
  NANDX1 G20197 (.A1(W9086), .A2(W36556), .ZN(O11940));
  NANDX1 G20198 (.A1(W32606), .A2(W22937), .ZN(O11939));
  NANDX1 G20199 (.A1(W27773), .A2(W23589), .ZN(W41905));
  NANDX1 G20200 (.A1(W12904), .A2(W40587), .ZN(W41900));
  NANDX1 G20201 (.A1(W39655), .A2(W13572), .ZN(O11929));
  NANDX1 G20202 (.A1(W27865), .A2(W8598), .ZN(O11926));
  NANDX1 G20203 (.A1(W35645), .A2(W4673), .ZN(W41889));
  NANDX1 G20204 (.A1(W29166), .A2(W31247), .ZN(O11921));
  NANDX1 G20205 (.A1(W37266), .A2(W9013), .ZN(W43377));
  NANDX1 G20206 (.A1(W24526), .A2(W28795), .ZN(O13107));
  NANDX1 G20207 (.A1(W7214), .A2(W30114), .ZN(W43414));
  NANDX1 G20208 (.A1(W16505), .A2(W37174), .ZN(W43404));
  NANDX1 G20209 (.A1(W17449), .A2(I407), .ZN(W43398));
  NANDX1 G20210 (.A1(W24012), .A2(W39652), .ZN(O13094));
  NANDX1 G20211 (.A1(W42964), .A2(W34892), .ZN(O13093));
  NANDX1 G20212 (.A1(W34258), .A2(W38680), .ZN(O13092));
  NANDX1 G20213 (.A1(W5918), .A2(W2956), .ZN(O13091));
  NANDX1 G20214 (.A1(W9167), .A2(W19235), .ZN(O13090));
  NANDX1 G20215 (.A1(W43004), .A2(W17615), .ZN(O13085));
  NANDX1 G20216 (.A1(W4651), .A2(W21575), .ZN(W43380));
  NANDX1 G20217 (.A1(W271), .A2(W26671), .ZN(O13082));
  NANDX1 G20218 (.A1(W15479), .A2(W23507), .ZN(O13111));
  NANDX1 G20219 (.A1(W1894), .A2(W18028), .ZN(O13079));
  NANDX1 G20220 (.A1(W15845), .A2(W27681), .ZN(O13078));
  NANDX1 G20221 (.A1(W22846), .A2(W31110), .ZN(W43373));
  NANDX1 G20222 (.A1(W8481), .A2(W33264), .ZN(O13077));
  NANDX1 G20223 (.A1(W32819), .A2(W3816), .ZN(O13076));
  NANDX1 G20224 (.A1(W41671), .A2(W32503), .ZN(O13074));
  NANDX1 G20225 (.A1(W22988), .A2(W38986), .ZN(O13073));
  NANDX1 G20226 (.A1(W20759), .A2(W6819), .ZN(O13071));
  NANDX1 G20227 (.A1(W268), .A2(W5043), .ZN(O13070));
  NANDX1 G20228 (.A1(W28142), .A2(W15263), .ZN(O13067));
  NANDX1 G20229 (.A1(W39619), .A2(W15392), .ZN(O13064));
  NANDX1 G20230 (.A1(W11491), .A2(W11071), .ZN(O13142));
  NANDX1 G20231 (.A1(W2253), .A2(W5878), .ZN(O13165));
  NANDX1 G20232 (.A1(W33097), .A2(W30472), .ZN(O13163));
  NANDX1 G20233 (.A1(W42797), .A2(W3048), .ZN(O13162));
  NANDX1 G20234 (.A1(W9222), .A2(W21756), .ZN(O13160));
  NANDX1 G20235 (.A1(W35360), .A2(W31917), .ZN(O13159));
  NANDX1 G20236 (.A1(W35214), .A2(W37621), .ZN(O13158));
  NANDX1 G20237 (.A1(W26229), .A2(W28958), .ZN(O13155));
  NANDX1 G20238 (.A1(W39070), .A2(W31953), .ZN(O13150));
  NANDX1 G20239 (.A1(W22164), .A2(W12161), .ZN(O13149));
  NANDX1 G20240 (.A1(W43465), .A2(W35175), .ZN(O13147));
  NANDX1 G20241 (.A1(W17443), .A2(W4806), .ZN(O13144));
  NANDX1 G20242 (.A1(W2794), .A2(W20198), .ZN(W43465));
  NANDX1 G20243 (.A1(W10888), .A2(W32056), .ZN(O13062));
  NANDX1 G20244 (.A1(W1289), .A2(W5532), .ZN(O13141));
  NANDX1 G20245 (.A1(W36514), .A2(W37500), .ZN(W43453));
  NANDX1 G20246 (.A1(W8963), .A2(W4933), .ZN(O13133));
  NANDX1 G20247 (.A1(W32238), .A2(W23055), .ZN(O13129));
  NANDX1 G20248 (.A1(W4141), .A2(W34643), .ZN(W43439));
  NANDX1 G20249 (.A1(W19316), .A2(W201), .ZN(O13123));
  NANDX1 G20250 (.A1(W38852), .A2(W42673), .ZN(O13122));
  NANDX1 G20251 (.A1(W15265), .A2(W36773), .ZN(O13120));
  NANDX1 G20252 (.A1(W32743), .A2(W28428), .ZN(O13118));
  NANDX1 G20253 (.A1(W1133), .A2(W5298), .ZN(O13113));
  NANDX1 G20254 (.A1(W40806), .A2(W26813), .ZN(O13112));
  NANDX1 G20255 (.A1(W27395), .A2(W38406), .ZN(O12974));
  NANDX1 G20256 (.A1(W959), .A2(W9230), .ZN(O13002));
  NANDX1 G20257 (.A1(W32234), .A2(W25175), .ZN(O13001));
  NANDX1 G20258 (.A1(W24810), .A2(W12140), .ZN(O13000));
  NANDX1 G20259 (.A1(W30610), .A2(W9830), .ZN(O12998));
  NANDX1 G20260 (.A1(W36002), .A2(W22449), .ZN(O12996));
  NANDX1 G20261 (.A1(W15845), .A2(W29800), .ZN(W43276));
  NANDX1 G20262 (.A1(W35359), .A2(W17797), .ZN(O12990));
  NANDX1 G20263 (.A1(W20991), .A2(W22357), .ZN(O12989));
  NANDX1 G20264 (.A1(W42499), .A2(W16807), .ZN(O12988));
  NANDX1 G20265 (.A1(W4103), .A2(W27650), .ZN(O12987));
  NANDX1 G20266 (.A1(W29941), .A2(W21669), .ZN(O12984));
  NANDX1 G20267 (.A1(W23909), .A2(W31408), .ZN(O12983));
  NANDX1 G20268 (.A1(W24302), .A2(W17899), .ZN(W43288));
  NANDX1 G20269 (.A1(W31431), .A2(W42306), .ZN(O12972));
  NANDX1 G20270 (.A1(W1053), .A2(W18964), .ZN(O12971));
  NANDX1 G20271 (.A1(W26707), .A2(W7262), .ZN(O12970));
  NANDX1 G20272 (.A1(W30961), .A2(W24212), .ZN(O12966));
  NANDX1 G20273 (.A1(W21471), .A2(W5916), .ZN(O12962));
  NANDX1 G20274 (.A1(W36168), .A2(W30910), .ZN(O12961));
  NANDX1 G20275 (.A1(I788), .A2(W18168), .ZN(O12960));
  NANDX1 G20276 (.A1(W901), .A2(W16374), .ZN(W43236));
  NANDX1 G20277 (.A1(W36807), .A2(W1361), .ZN(O12957));
  NANDX1 G20278 (.A1(W7488), .A2(W10925), .ZN(O12955));
  NANDX1 G20279 (.A1(W33902), .A2(W36650), .ZN(W43232));
  NANDX1 G20280 (.A1(W9406), .A2(W21173), .ZN(O13043));
  NANDX1 G20281 (.A1(W15176), .A2(W9540), .ZN(W43353));
  NANDX1 G20282 (.A1(W29481), .A2(W30170), .ZN(O13061));
  NANDX1 G20283 (.A1(W40068), .A2(I1231), .ZN(O13059));
  NANDX1 G20284 (.A1(W17950), .A2(W13021), .ZN(O13054));
  NANDX1 G20285 (.A1(W30930), .A2(W36634), .ZN(O13053));
  NANDX1 G20286 (.A1(W33327), .A2(W22832), .ZN(O13052));
  NANDX1 G20287 (.A1(W3131), .A2(W20030), .ZN(O13051));
  NANDX1 G20288 (.A1(W11006), .A2(W41512), .ZN(O13050));
  NANDX1 G20289 (.A1(W9957), .A2(W38771), .ZN(O13048));
  NANDX1 G20290 (.A1(W38580), .A2(W12514), .ZN(O13046));
  NANDX1 G20291 (.A1(W28659), .A2(W3946), .ZN(O13044));
  NANDX1 G20292 (.A1(W31686), .A2(W598), .ZN(O13166));
  NANDX1 G20293 (.A1(W10138), .A2(W42881), .ZN(O13041));
  NANDX1 G20294 (.A1(W34091), .A2(W12119), .ZN(O13039));
  NANDX1 G20295 (.A1(W22562), .A2(W840), .ZN(O13038));
  NANDX1 G20296 (.A1(W14004), .A2(W31242), .ZN(O13036));
  NANDX1 G20297 (.A1(W28695), .A2(W20497), .ZN(O13032));
  NANDX1 G20298 (.A1(W43033), .A2(W12301), .ZN(W43319));
  NANDX1 G20299 (.A1(W18223), .A2(W25041), .ZN(O13027));
  NANDX1 G20300 (.A1(W40789), .A2(W21542), .ZN(O13020));
  NANDX1 G20301 (.A1(W40783), .A2(W13805), .ZN(O13017));
  NANDX1 G20302 (.A1(W13350), .A2(W11187), .ZN(O13014));
  NANDX1 G20303 (.A1(W37541), .A2(W36042), .ZN(O13007));
  NANDX1 G20304 (.A1(W1095), .A2(W23753), .ZN(O13313));
  NANDX1 G20305 (.A1(W8052), .A2(I1749), .ZN(O13347));
  NANDX1 G20306 (.A1(W43580), .A2(W20240), .ZN(O13343));
  NANDX1 G20307 (.A1(W27220), .A2(W15152), .ZN(W43732));
  NANDX1 G20308 (.A1(W11485), .A2(W20301), .ZN(O13342));
  NANDX1 G20309 (.A1(W30852), .A2(W29063), .ZN(O13340));
  NANDX1 G20310 (.A1(W38932), .A2(W18949), .ZN(O13339));
  NANDX1 G20311 (.A1(W19811), .A2(W1747), .ZN(O13332));
  NANDX1 G20312 (.A1(W43002), .A2(W7148), .ZN(O13331));
  NANDX1 G20313 (.A1(W23517), .A2(W12513), .ZN(O13329));
  NANDX1 G20314 (.A1(W33934), .A2(W21462), .ZN(O13324));
  NANDX1 G20315 (.A1(W15917), .A2(W13887), .ZN(W43710));
  NANDX1 G20316 (.A1(I1450), .A2(W40839), .ZN(O13317));
  NANDX1 G20317 (.A1(W13864), .A2(W11456), .ZN(O13348));
  NANDX1 G20318 (.A1(W14663), .A2(W34831), .ZN(O13312));
  NANDX1 G20319 (.A1(W18818), .A2(W27618), .ZN(O13309));
  NANDX1 G20320 (.A1(W33869), .A2(W3788), .ZN(O13306));
  NANDX1 G20321 (.A1(I1544), .A2(W42122), .ZN(O13305));
  NANDX1 G20322 (.A1(W28327), .A2(W6675), .ZN(W43684));
  NANDX1 G20323 (.A1(W27438), .A2(I677), .ZN(W43681));
  NANDX1 G20324 (.A1(W9903), .A2(W15022), .ZN(O13295));
  NANDX1 G20325 (.A1(W34448), .A2(W1541), .ZN(O13293));
  NANDX1 G20326 (.A1(W26540), .A2(W16297), .ZN(O13291));
  NANDX1 G20327 (.A1(W17278), .A2(W33577), .ZN(O13290));
  NANDX1 G20328 (.A1(W15744), .A2(W42778), .ZN(O13288));
  NANDX1 G20329 (.A1(W38493), .A2(I36), .ZN(O13367));
  NANDX1 G20330 (.A1(W25600), .A2(W29303), .ZN(O13391));
  NANDX1 G20331 (.A1(W5738), .A2(W21968), .ZN(O13390));
  NANDX1 G20332 (.A1(W29265), .A2(W43678), .ZN(W43786));
  NANDX1 G20333 (.A1(W38403), .A2(W19128), .ZN(O13380));
  NANDX1 G20334 (.A1(W1316), .A2(W1572), .ZN(O13378));
  NANDX1 G20335 (.A1(W26512), .A2(W12612), .ZN(O13377));
  NANDX1 G20336 (.A1(W35353), .A2(W24897), .ZN(O13374));
  NANDX1 G20337 (.A1(W14687), .A2(W36092), .ZN(O13373));
  NANDX1 G20338 (.A1(W42499), .A2(W2087), .ZN(O13372));
  NANDX1 G20339 (.A1(W36661), .A2(W2535), .ZN(O13368));
  NANDX1 G20340 (.A1(W13385), .A2(W42366), .ZN(W43766));
  NANDX1 G20341 (.A1(W30214), .A2(W35903), .ZN(W43765));
  NANDX1 G20342 (.A1(W6868), .A2(W41149), .ZN(W43652));
  NANDX1 G20343 (.A1(W33832), .A2(W613), .ZN(O13364));
  NANDX1 G20344 (.A1(W6868), .A2(W16201), .ZN(W43757));
  NANDX1 G20345 (.A1(W31908), .A2(W15957), .ZN(W43755));
  NANDX1 G20346 (.A1(W28405), .A2(W42739), .ZN(O13358));
  NANDX1 G20347 (.A1(W28484), .A2(W36605), .ZN(W43750));
  NANDX1 G20348 (.A1(W32379), .A2(W1883), .ZN(O13356));
  NANDX1 G20349 (.A1(W3911), .A2(W41015), .ZN(O13355));
  NANDX1 G20350 (.A1(W4220), .A2(W25944), .ZN(O13354));
  NANDX1 G20351 (.A1(W14341), .A2(W36070), .ZN(O13353));
  NANDX1 G20352 (.A1(W22345), .A2(W11149), .ZN(O13350));
  NANDX1 G20353 (.A1(W10310), .A2(W39289), .ZN(O13349));
  NANDX1 G20354 (.A1(W35800), .A2(W22731), .ZN(O13192));
  NANDX1 G20355 (.A1(W34995), .A2(W11688), .ZN(O13222));
  NANDX1 G20356 (.A1(W26565), .A2(W10283), .ZN(O13218));
  NANDX1 G20357 (.A1(W31096), .A2(W9298), .ZN(W43557));
  NANDX1 G20358 (.A1(W4021), .A2(W12222), .ZN(W43556));
  NANDX1 G20359 (.A1(W24288), .A2(W26796), .ZN(W43555));
  NANDX1 G20360 (.A1(W10182), .A2(W22925), .ZN(O13212));
  NANDX1 G20361 (.A1(W7718), .A2(W34986), .ZN(O13206));
  NANDX1 G20362 (.A1(W13012), .A2(W25189), .ZN(W43542));
  NANDX1 G20363 (.A1(W807), .A2(W20258), .ZN(O13201));
  NANDX1 G20364 (.A1(W31279), .A2(W13880), .ZN(W43538));
  NANDX1 G20365 (.A1(W19582), .A2(W6553), .ZN(O13200));
  NANDX1 G20366 (.A1(W27859), .A2(W39310), .ZN(O13194));
  NANDX1 G20367 (.A1(W41772), .A2(W10191), .ZN(O13223));
  NANDX1 G20368 (.A1(W19137), .A2(W25541), .ZN(O13191));
  NANDX1 G20369 (.A1(W12453), .A2(W7260), .ZN(O13184));
  NANDX1 G20370 (.A1(W41393), .A2(W22066), .ZN(W43511));
  NANDX1 G20371 (.A1(W18392), .A2(W17537), .ZN(O13183));
  NANDX1 G20372 (.A1(W5530), .A2(W36955), .ZN(O13178));
  NANDX1 G20373 (.A1(W27337), .A2(W28473), .ZN(O13177));
  NANDX1 G20374 (.A1(W32033), .A2(W34859), .ZN(O13176));
  NANDX1 G20375 (.A1(W17287), .A2(W9917), .ZN(O13175));
  NANDX1 G20376 (.A1(W37453), .A2(W10359), .ZN(O13174));
  NANDX1 G20377 (.A1(W41164), .A2(W39459), .ZN(O13168));
  NANDX1 G20378 (.A1(W2976), .A2(W7929), .ZN(W43492));
  NANDX1 G20379 (.A1(W12628), .A2(W29299), .ZN(W43618));
  NANDX1 G20380 (.A1(W6486), .A2(W39652), .ZN(O13283));
  NANDX1 G20381 (.A1(W14914), .A2(W8832), .ZN(O13281));
  NANDX1 G20382 (.A1(W10821), .A2(I1442), .ZN(W43645));
  NANDX1 G20383 (.A1(W22162), .A2(W2135), .ZN(W43643));
  NANDX1 G20384 (.A1(W5311), .A2(W6664), .ZN(O13277));
  NANDX1 G20385 (.A1(W24311), .A2(W27719), .ZN(W43637));
  NANDX1 G20386 (.A1(W22252), .A2(W26071), .ZN(W43635));
  NANDX1 G20387 (.A1(W39233), .A2(W18513), .ZN(W43631));
  NANDX1 G20388 (.A1(W27735), .A2(W34302), .ZN(W43630));
  NANDX1 G20389 (.A1(W13783), .A2(W18428), .ZN(O13269));
  NANDX1 G20390 (.A1(W29637), .A2(W32247), .ZN(O13266));
  NANDX1 G20391 (.A1(W41110), .A2(W17652), .ZN(O12949));
  NANDX1 G20392 (.A1(W4496), .A2(W42822), .ZN(O13258));
  NANDX1 G20393 (.A1(W25627), .A2(W25115), .ZN(O13257));
  NANDX1 G20394 (.A1(W25490), .A2(W28862), .ZN(O13247));
  NANDX1 G20395 (.A1(W10609), .A2(W38115), .ZN(O13245));
  NANDX1 G20396 (.A1(W1794), .A2(W12829), .ZN(O13243));
  NANDX1 G20397 (.A1(W19613), .A2(W31288), .ZN(O13238));
  NANDX1 G20398 (.A1(W30610), .A2(W9907), .ZN(O13237));
  NANDX1 G20399 (.A1(W14511), .A2(W14335), .ZN(O13236));
  NANDX1 G20400 (.A1(W3783), .A2(W4611), .ZN(O13234));
  NANDX1 G20401 (.A1(W21670), .A2(W18830), .ZN(O13228));
  NANDX1 G20402 (.A1(W9087), .A2(W37932), .ZN(O13226));
  NANDX1 G20403 (.A1(W35415), .A2(W9869), .ZN(W42838));
  NANDX1 G20404 (.A1(W33121), .A2(W1196), .ZN(O12674));
  NANDX1 G20405 (.A1(W21340), .A2(W4968), .ZN(O12670));
  NANDX1 G20406 (.A1(W34702), .A2(W28833), .ZN(W42857));
  NANDX1 G20407 (.A1(W37883), .A2(W3299), .ZN(O12664));
  NANDX1 G20408 (.A1(W38252), .A2(W7423), .ZN(O12663));
  NANDX1 G20409 (.A1(W26035), .A2(W38132), .ZN(O12662));
  NANDX1 G20410 (.A1(W6772), .A2(W1158), .ZN(O12661));
  NANDX1 G20411 (.A1(W6407), .A2(W4715), .ZN(O12660));
  NANDX1 G20412 (.A1(W16492), .A2(W35016), .ZN(O12657));
  NANDX1 G20413 (.A1(W6768), .A2(W40423), .ZN(O12656));
  NANDX1 G20414 (.A1(W1072), .A2(W20497), .ZN(O12655));
  NANDX1 G20415 (.A1(W37643), .A2(W39877), .ZN(O12652));
  NANDX1 G20416 (.A1(W4943), .A2(W3247), .ZN(O12678));
  NANDX1 G20417 (.A1(W4784), .A2(W11517), .ZN(O12651));
  NANDX1 G20418 (.A1(W9344), .A2(W24958), .ZN(O12650));
  NANDX1 G20419 (.A1(W37592), .A2(W33280), .ZN(O12646));
  NANDX1 G20420 (.A1(W9929), .A2(W1213), .ZN(O12644));
  NANDX1 G20421 (.A1(W33198), .A2(W36650), .ZN(O12642));
  NANDX1 G20422 (.A1(W17398), .A2(I437), .ZN(O12641));
  NANDX1 G20423 (.A1(W15410), .A2(W39870), .ZN(W42823));
  NANDX1 G20424 (.A1(W11758), .A2(W12644), .ZN(W42822));
  NANDX1 G20425 (.A1(W16724), .A2(W17975), .ZN(O12639));
  NANDX1 G20426 (.A1(W26784), .A2(W15275), .ZN(O12635));
  NANDX1 G20427 (.A1(W25839), .A2(W18278), .ZN(O12633));
  NANDX1 G20428 (.A1(W9566), .A2(W10711), .ZN(W42893));
  NANDX1 G20429 (.A1(W20839), .A2(I1389), .ZN(O12720));
  NANDX1 G20430 (.A1(W314), .A2(W34379), .ZN(O12719));
  NANDX1 G20431 (.A1(W18379), .A2(W36418), .ZN(W42928));
  NANDX1 G20432 (.A1(W14825), .A2(W30439), .ZN(O12715));
  NANDX1 G20433 (.A1(W460), .A2(W33698), .ZN(W42922));
  NANDX1 G20434 (.A1(W3346), .A2(W33221), .ZN(O12703));
  NANDX1 G20435 (.A1(W9590), .A2(W18244), .ZN(W42908));
  NANDX1 G20436 (.A1(W30253), .A2(W26010), .ZN(O12700));
  NANDX1 G20437 (.A1(W33386), .A2(W9226), .ZN(O12696));
  NANDX1 G20438 (.A1(I683), .A2(W33021), .ZN(W42901));
  NANDX1 G20439 (.A1(W31506), .A2(W28587), .ZN(W42900));
  NANDX1 G20440 (.A1(W2409), .A2(W13317), .ZN(O12694));
  NANDX1 G20441 (.A1(W16406), .A2(W10226), .ZN(O12630));
  NANDX1 G20442 (.A1(W26232), .A2(W29900), .ZN(W42891));
  NANDX1 G20443 (.A1(W22425), .A2(W10351), .ZN(W42890));
  NANDX1 G20444 (.A1(W13034), .A2(W36989), .ZN(O12689));
  NANDX1 G20445 (.A1(W1310), .A2(W25445), .ZN(O12688));
  NANDX1 G20446 (.A1(W24439), .A2(W1978), .ZN(O12686));
  NANDX1 G20447 (.A1(W7121), .A2(W31288), .ZN(O12685));
  NANDX1 G20448 (.A1(W13788), .A2(W41106), .ZN(O12684));
  NANDX1 G20449 (.A1(W3251), .A2(W42372), .ZN(W42881));
  NANDX1 G20450 (.A1(W38061), .A2(W27266), .ZN(O12683));
  NANDX1 G20451 (.A1(W28730), .A2(W34672), .ZN(O12682));
  NANDX1 G20452 (.A1(W39933), .A2(W11746), .ZN(O12680));
  NANDX1 G20453 (.A1(W16705), .A2(W7071), .ZN(O12562));
  NANDX1 G20454 (.A1(W4504), .A2(W2745), .ZN(O12586));
  NANDX1 G20455 (.A1(W763), .A2(W37625), .ZN(O12581));
  NANDX1 G20456 (.A1(W10013), .A2(W40008), .ZN(O12578));
  NANDX1 G20457 (.A1(W13589), .A2(W28820), .ZN(W42739));
  NANDX1 G20458 (.A1(W15370), .A2(W18348), .ZN(O12577));
  NANDX1 G20459 (.A1(W11108), .A2(W23589), .ZN(O12576));
  NANDX1 G20460 (.A1(W42673), .A2(W10426), .ZN(O12575));
  NANDX1 G20461 (.A1(W6622), .A2(W24937), .ZN(O12573));
  NANDX1 G20462 (.A1(W41855), .A2(W10572), .ZN(W42731));
  NANDX1 G20463 (.A1(W40952), .A2(W30524), .ZN(O12572));
  NANDX1 G20464 (.A1(W1671), .A2(W24892), .ZN(O12571));
  NANDX1 G20465 (.A1(W10589), .A2(W22610), .ZN(O12570));
  NANDX1 G20466 (.A1(W2924), .A2(W26844), .ZN(O12587));
  NANDX1 G20467 (.A1(W30176), .A2(W37188), .ZN(W42717));
  NANDX1 G20468 (.A1(W30806), .A2(W38637), .ZN(O12554));
  NANDX1 G20469 (.A1(W4075), .A2(W29965), .ZN(W42707));
  NANDX1 G20470 (.A1(W23577), .A2(W15425), .ZN(O12552));
  NANDX1 G20471 (.A1(W289), .A2(W38688), .ZN(O12550));
  NANDX1 G20472 (.A1(W17266), .A2(W1600), .ZN(W42699));
  NANDX1 G20473 (.A1(W40737), .A2(W8010), .ZN(O12544));
  NANDX1 G20474 (.A1(W34078), .A2(W28024), .ZN(O12541));
  NANDX1 G20475 (.A1(W32366), .A2(W5338), .ZN(O12540));
  NANDX1 G20476 (.A1(W31254), .A2(W6445), .ZN(O12539));
  NANDX1 G20477 (.A1(W7997), .A2(W30025), .ZN(O12534));
  NANDX1 G20478 (.A1(W39186), .A2(W1874), .ZN(O12608));
  NANDX1 G20479 (.A1(W26474), .A2(W19471), .ZN(O12626));
  NANDX1 G20480 (.A1(W38172), .A2(W34047), .ZN(W42805));
  NANDX1 G20481 (.A1(W32281), .A2(W5210), .ZN(O12620));
  NANDX1 G20482 (.A1(W16507), .A2(W32240), .ZN(O12619));
  NANDX1 G20483 (.A1(W15817), .A2(W21754), .ZN(W42797));
  NANDX1 G20484 (.A1(W33518), .A2(W25949), .ZN(W42791));
  NANDX1 G20485 (.A1(W30808), .A2(W10435), .ZN(W42790));
  NANDX1 G20486 (.A1(W25901), .A2(W38435), .ZN(O12614));
  NANDX1 G20487 (.A1(W22831), .A2(W29099), .ZN(O12613));
  NANDX1 G20488 (.A1(W17833), .A2(W32859), .ZN(W42786));
  NANDX1 G20489 (.A1(W29265), .A2(W24073), .ZN(O12612));
  NANDX1 G20490 (.A1(W21595), .A2(W22805), .ZN(O12725));
  NANDX1 G20491 (.A1(W22121), .A2(I798), .ZN(W42778));
  NANDX1 G20492 (.A1(W32796), .A2(W16741), .ZN(O12606));
  NANDX1 G20493 (.A1(W37395), .A2(W37136), .ZN(O12603));
  NANDX1 G20494 (.A1(W18143), .A2(W7772), .ZN(O12602));
  NANDX1 G20495 (.A1(W6171), .A2(W42218), .ZN(O12601));
  NANDX1 G20496 (.A1(W3542), .A2(W6264), .ZN(O12600));
  NANDX1 G20497 (.A1(W38601), .A2(W1391), .ZN(O12596));
  NANDX1 G20498 (.A1(W15932), .A2(W33444), .ZN(O12595));
  NANDX1 G20499 (.A1(W16464), .A2(W9345), .ZN(O12591));
  NANDX1 G20500 (.A1(W30716), .A2(W15709), .ZN(W42754));
  NANDX1 G20501 (.A1(I1175), .A2(W11834), .ZN(O12589));
  NANDX1 G20502 (.A1(W7008), .A2(W22730), .ZN(O12857));
  NANDX1 G20503 (.A1(W14183), .A2(W38627), .ZN(O12886));
  NANDX1 G20504 (.A1(W28938), .A2(W6491), .ZN(O12884));
  NANDX1 G20505 (.A1(W2404), .A2(W27322), .ZN(O12881));
  NANDX1 G20506 (.A1(W15155), .A2(W18470), .ZN(W43142));
  NANDX1 G20507 (.A1(W23062), .A2(W13507), .ZN(O12880));
  NANDX1 G20508 (.A1(W12860), .A2(W28072), .ZN(O12873));
  NANDX1 G20509 (.A1(W22953), .A2(W34093), .ZN(O12869));
  NANDX1 G20510 (.A1(W12555), .A2(W8803), .ZN(W43122));
  NANDX1 G20511 (.A1(W16431), .A2(W17718), .ZN(O12866));
  NANDX1 G20512 (.A1(W41114), .A2(W9193), .ZN(W43119));
  NANDX1 G20513 (.A1(W12691), .A2(W22114), .ZN(O12865));
  NANDX1 G20514 (.A1(W15413), .A2(W3430), .ZN(O12862));
  NANDX1 G20515 (.A1(W1011), .A2(W31168), .ZN(O12890));
  NANDX1 G20516 (.A1(W38876), .A2(W56), .ZN(O12856));
  NANDX1 G20517 (.A1(W42452), .A2(W31934), .ZN(O12855));
  NANDX1 G20518 (.A1(W6940), .A2(W1222), .ZN(W43103));
  NANDX1 G20519 (.A1(W23927), .A2(W23783), .ZN(W43100));
  NANDX1 G20520 (.A1(W32155), .A2(W38421), .ZN(O12848));
  NANDX1 G20521 (.A1(W28576), .A2(W28934), .ZN(O12845));
  NANDX1 G20522 (.A1(W35429), .A2(W17579), .ZN(O12844));
  NANDX1 G20523 (.A1(W36240), .A2(W16824), .ZN(O12842));
  NANDX1 G20524 (.A1(W41012), .A2(I1220), .ZN(O12838));
  NANDX1 G20525 (.A1(W13981), .A2(W36989), .ZN(O12837));
  NANDX1 G20526 (.A1(W40721), .A2(W25297), .ZN(O12833));
  NANDX1 G20527 (.A1(W22448), .A2(W33429), .ZN(W43186));
  NANDX1 G20528 (.A1(W16281), .A2(W8139), .ZN(O12947));
  NANDX1 G20529 (.A1(W12079), .A2(W7337), .ZN(O12943));
  NANDX1 G20530 (.A1(W9786), .A2(W3121), .ZN(W43216));
  NANDX1 G20531 (.A1(W6549), .A2(W15507), .ZN(O12941));
  NANDX1 G20532 (.A1(W26647), .A2(W39980), .ZN(O12940));
  NANDX1 G20533 (.A1(W14089), .A2(W22594), .ZN(O12937));
  NANDX1 G20534 (.A1(W41661), .A2(W1265), .ZN(W43208));
  NANDX1 G20535 (.A1(W34808), .A2(W6966), .ZN(W43205));
  NANDX1 G20536 (.A1(W42146), .A2(W6134), .ZN(O12933));
  NANDX1 G20537 (.A1(W35881), .A2(W18748), .ZN(O12932));
  NANDX1 G20538 (.A1(W12063), .A2(W3459), .ZN(O12919));
  NANDX1 G20539 (.A1(W38477), .A2(W12341), .ZN(W43075));
  NANDX1 G20540 (.A1(W8286), .A2(W15532), .ZN(O12917));
  NANDX1 G20541 (.A1(W42770), .A2(W13066), .ZN(O12916));
  NANDX1 G20542 (.A1(I594), .A2(W38133), .ZN(O12911));
  NANDX1 G20543 (.A1(W41203), .A2(W37506), .ZN(W43176));
  NANDX1 G20544 (.A1(W31307), .A2(W31903), .ZN(O12907));
  NANDX1 G20545 (.A1(W28070), .A2(W2118), .ZN(O12905));
  NANDX1 G20546 (.A1(W19313), .A2(W29936), .ZN(O12904));
  NANDX1 G20547 (.A1(W9884), .A2(W2021), .ZN(O12902));
  NANDX1 G20548 (.A1(W38745), .A2(I1331), .ZN(O12901));
  NANDX1 G20549 (.A1(W14189), .A2(W32351), .ZN(O12898));
  NANDX1 G20550 (.A1(W20135), .A2(W31338), .ZN(O12895));
  NANDX1 G20551 (.A1(W38776), .A2(W21499), .ZN(W42979));
  NANDX1 G20552 (.A1(W16461), .A2(W3427), .ZN(O12779));
  NANDX1 G20553 (.A1(W38004), .A2(W18129), .ZN(O12778));
  NANDX1 G20554 (.A1(W16155), .A2(W22072), .ZN(O12775));
  NANDX1 G20555 (.A1(W29408), .A2(W35033), .ZN(O12771));
  NANDX1 G20556 (.A1(W25683), .A2(W34972), .ZN(O12770));
  NANDX1 G20557 (.A1(W11902), .A2(W40466), .ZN(O12769));
  NANDX1 G20558 (.A1(W32491), .A2(W21222), .ZN(O12767));
  NANDX1 G20559 (.A1(W26681), .A2(W4760), .ZN(O12766));
  NANDX1 G20560 (.A1(W4923), .A2(W24818), .ZN(O12764));
  NANDX1 G20561 (.A1(W3298), .A2(W10755), .ZN(W42983));
  NANDX1 G20562 (.A1(W1161), .A2(W35629), .ZN(O12758));
  NANDX1 G20563 (.A1(W40502), .A2(W35824), .ZN(W42981));
  NANDX1 G20564 (.A1(W42363), .A2(W478), .ZN(O12780));
  NANDX1 G20565 (.A1(W1335), .A2(W35035), .ZN(W42976));
  NANDX1 G20566 (.A1(W34593), .A2(W39161), .ZN(O12746));
  NANDX1 G20567 (.A1(W12582), .A2(W27599), .ZN(O12743));
  NANDX1 G20568 (.A1(W13739), .A2(W18164), .ZN(O12742));
  NANDX1 G20569 (.A1(W22131), .A2(W42032), .ZN(O12741));
  NANDX1 G20570 (.A1(W41680), .A2(W42327), .ZN(W42958));
  NANDX1 G20571 (.A1(W21256), .A2(W18745), .ZN(O12738));
  NANDX1 G20572 (.A1(W8965), .A2(W18187), .ZN(O12737));
  NANDX1 G20573 (.A1(W35198), .A2(W42220), .ZN(O12733));
  NANDX1 G20574 (.A1(W21372), .A2(W15006), .ZN(O12730));
  NANDX1 G20575 (.A1(W40866), .A2(W14995), .ZN(O12728));
  NANDX1 G20576 (.A1(W3251), .A2(W10562), .ZN(O12808));
  NANDX1 G20577 (.A1(W20068), .A2(W614), .ZN(O12832));
  NANDX1 G20578 (.A1(W1048), .A2(W34768), .ZN(O12831));
  NANDX1 G20579 (.A1(W16293), .A2(W14434), .ZN(O12828));
  NANDX1 G20580 (.A1(W24710), .A2(W7068), .ZN(O12826));
  NANDX1 G20581 (.A1(W2843), .A2(W7906), .ZN(O12824));
  NANDX1 G20582 (.A1(W12715), .A2(W6175), .ZN(O12820));
  NANDX1 G20583 (.A1(W40225), .A2(W18930), .ZN(O12818));
  NANDX1 G20584 (.A1(W26138), .A2(W3693), .ZN(O12815));
  NANDX1 G20585 (.A1(W5931), .A2(W15002), .ZN(W43054));
  NANDX1 G20586 (.A1(W29036), .A2(W24815), .ZN(W43051));
  NANDX1 G20587 (.A1(W4358), .A2(W12519), .ZN(O12811));
  NANDX1 G20588 (.A1(W29280), .A2(W3006), .ZN(O15374));
  NANDX1 G20589 (.A1(W3982), .A2(W4911), .ZN(O12804));
  NANDX1 G20590 (.A1(W34302), .A2(W14509), .ZN(O12803));
  NANDX1 G20591 (.A1(W35448), .A2(W42311), .ZN(O12797));
  NANDX1 G20592 (.A1(W8878), .A2(W13162), .ZN(O12796));
  NANDX1 G20593 (.A1(W6177), .A2(W38185), .ZN(W43025));
  NANDX1 G20594 (.A1(W16960), .A2(W36978), .ZN(W43022));
  NANDX1 G20595 (.A1(W4983), .A2(W17642), .ZN(O12788));
  NANDX1 G20596 (.A1(W37979), .A2(W14984), .ZN(O12786));
  NANDX1 G20597 (.A1(W150), .A2(W39025), .ZN(O12785));
  NANDX1 G20598 (.A1(W33612), .A2(W23061), .ZN(W43017));
  NANDX1 G20599 (.A1(W11525), .A2(W37564), .ZN(O12783));
  NANDX1 G20600 (.A1(W36672), .A2(W46432), .ZN(O18230));
  NANDX1 G20601 (.A1(W14679), .A2(W24627), .ZN(O18265));
  NANDX1 G20602 (.A1(W5744), .A2(W33668), .ZN(O18263));
  NANDX1 G20603 (.A1(W35321), .A2(W48790), .ZN(O18254));
  NANDX1 G20604 (.A1(W30428), .A2(W18061), .ZN(O18253));
  NANDX1 G20605 (.A1(W17054), .A2(W48899), .ZN(O18247));
  NANDX1 G20606 (.A1(W41160), .A2(W12873), .ZN(W49437));
  NANDX1 G20607 (.A1(W37208), .A2(W31318), .ZN(O18241));
  NANDX1 G20608 (.A1(W348), .A2(W45281), .ZN(W49433));
  NANDX1 G20609 (.A1(W24651), .A2(I1681), .ZN(O18238));
  NANDX1 G20610 (.A1(W4544), .A2(W31252), .ZN(O18235));
  NANDX1 G20611 (.A1(W35160), .A2(W45111), .ZN(O18232));
  NANDX1 G20612 (.A1(W7514), .A2(W16627), .ZN(O18231));
  NANDX1 G20613 (.A1(W18719), .A2(W13768), .ZN(O18270));
  NANDX1 G20614 (.A1(W29521), .A2(W10082), .ZN(O18219));
  NANDX1 G20615 (.A1(W28296), .A2(W4267), .ZN(O18214));
  NANDX1 G20616 (.A1(W39312), .A2(W35138), .ZN(O18213));
  NANDX1 G20617 (.A1(W5364), .A2(W3659), .ZN(O18210));
  NANDX1 G20618 (.A1(W12908), .A2(W35373), .ZN(O18206));
  NANDX1 G20619 (.A1(W18977), .A2(W34594), .ZN(O18203));
  NANDX1 G20620 (.A1(W3500), .A2(W12244), .ZN(O18201));
  NANDX1 G20621 (.A1(W35787), .A2(W2986), .ZN(O18195));
  NANDX1 G20622 (.A1(W17961), .A2(W22220), .ZN(O18194));
  NANDX1 G20623 (.A1(W9371), .A2(W8944), .ZN(O18193));
  NANDX1 G20624 (.A1(W28234), .A2(W33563), .ZN(O18189));
  NANDX1 G20625 (.A1(W27244), .A2(W40296), .ZN(O18304));
  NANDX1 G20626 (.A1(W18129), .A2(W46486), .ZN(O18338));
  NANDX1 G20627 (.A1(W48556), .A2(W19607), .ZN(O18335));
  NANDX1 G20628 (.A1(W9811), .A2(W32321), .ZN(O18334));
  NANDX1 G20629 (.A1(W8455), .A2(W1694), .ZN(O18332));
  NANDX1 G20630 (.A1(W27202), .A2(W31274), .ZN(O18331));
  NANDX1 G20631 (.A1(W9116), .A2(W34050), .ZN(W49527));
  NANDX1 G20632 (.A1(W10803), .A2(W24949), .ZN(O18327));
  NANDX1 G20633 (.A1(W11703), .A2(W38992), .ZN(O18323));
  NANDX1 G20634 (.A1(W11580), .A2(W26346), .ZN(O18319));
  NANDX1 G20635 (.A1(W18019), .A2(W32962), .ZN(O18309));
  NANDX1 G20636 (.A1(W38398), .A2(W31318), .ZN(O18308));
  NANDX1 G20637 (.A1(W48256), .A2(W21006), .ZN(O18307));
  NANDX1 G20638 (.A1(W43122), .A2(W48074), .ZN(O18188));
  NANDX1 G20639 (.A1(W7780), .A2(W6978), .ZN(O18303));
  NANDX1 G20640 (.A1(W22135), .A2(W4551), .ZN(O18298));
  NANDX1 G20641 (.A1(W23028), .A2(W28824), .ZN(O18293));
  NANDX1 G20642 (.A1(W14607), .A2(W9358), .ZN(O18292));
  NANDX1 G20643 (.A1(W14802), .A2(W6941), .ZN(O18291));
  NANDX1 G20644 (.A1(W21699), .A2(W14034), .ZN(O18288));
  NANDX1 G20645 (.A1(W6233), .A2(W26866), .ZN(O18286));
  NANDX1 G20646 (.A1(W1368), .A2(W25974), .ZN(O18282));
  NANDX1 G20647 (.A1(W10473), .A2(W333), .ZN(O18281));
  NANDX1 G20648 (.A1(I579), .A2(W24082), .ZN(O18279));
  NANDX1 G20649 (.A1(W30900), .A2(I1000), .ZN(O18273));
  NANDX1 G20650 (.A1(W8356), .A2(W33279), .ZN(O18105));
  NANDX1 G20651 (.A1(W10193), .A2(W18296), .ZN(O18143));
  NANDX1 G20652 (.A1(W34659), .A2(W17465), .ZN(O18141));
  NANDX1 G20653 (.A1(W6104), .A2(W4278), .ZN(O18138));
  NANDX1 G20654 (.A1(W34387), .A2(W33079), .ZN(O18132));
  NANDX1 G20655 (.A1(W37642), .A2(W11931), .ZN(O18131));
  NANDX1 G20656 (.A1(W16240), .A2(I1450), .ZN(O18128));
  NANDX1 G20657 (.A1(W44182), .A2(I748), .ZN(O18126));
  NANDX1 G20658 (.A1(W35634), .A2(W32203), .ZN(O18122));
  NANDX1 G20659 (.A1(W24128), .A2(W27060), .ZN(O18120));
  NANDX1 G20660 (.A1(W22275), .A2(W25413), .ZN(O18115));
  NANDX1 G20661 (.A1(W35194), .A2(W14093), .ZN(O18114));
  NANDX1 G20662 (.A1(W42351), .A2(W26025), .ZN(O18111));
  NANDX1 G20663 (.A1(W29274), .A2(W11560), .ZN(O18144));
  NANDX1 G20664 (.A1(W20630), .A2(W24685), .ZN(O18104));
  NANDX1 G20665 (.A1(W43896), .A2(W48437), .ZN(O18092));
  NANDX1 G20666 (.A1(W43462), .A2(W45980), .ZN(W49276));
  NANDX1 G20667 (.A1(W34008), .A2(W4832), .ZN(O18088));
  NANDX1 G20668 (.A1(W7189), .A2(W28177), .ZN(O18078));
  NANDX1 G20669 (.A1(W34959), .A2(W30581), .ZN(O18075));
  NANDX1 G20670 (.A1(W15233), .A2(W17957), .ZN(O18074));
  NANDX1 G20671 (.A1(W2417), .A2(W24975), .ZN(O18073));
  NANDX1 G20672 (.A1(W40128), .A2(W23021), .ZN(O18062));
  NANDX1 G20673 (.A1(W19013), .A2(W13828), .ZN(O18057));
  NANDX1 G20674 (.A1(W24284), .A2(W506), .ZN(O18056));
  NANDX1 G20675 (.A1(W42307), .A2(W2214), .ZN(O18165));
  NANDX1 G20676 (.A1(W37455), .A2(W48664), .ZN(W49379));
  NANDX1 G20677 (.A1(W2493), .A2(W2849), .ZN(O18182));
  NANDX1 G20678 (.A1(W17623), .A2(W28491), .ZN(O18180));
  NANDX1 G20679 (.A1(W16488), .A2(W27139), .ZN(W49368));
  NANDX1 G20680 (.A1(W45569), .A2(W10722), .ZN(O18177));
  NANDX1 G20681 (.A1(W39660), .A2(W44077), .ZN(O18175));
  NANDX1 G20682 (.A1(W24461), .A2(W46660), .ZN(O18174));
  NANDX1 G20683 (.A1(W10806), .A2(W36630), .ZN(O18172));
  NANDX1 G20684 (.A1(W33968), .A2(W11936), .ZN(O18171));
  NANDX1 G20685 (.A1(W16760), .A2(W24031), .ZN(O18167));
  NANDX1 G20686 (.A1(W47120), .A2(W17695), .ZN(O18166));
  NANDX1 G20687 (.A1(W36175), .A2(W34339), .ZN(O18340));
  NANDX1 G20688 (.A1(W14563), .A2(W46218), .ZN(O18160));
  NANDX1 G20689 (.A1(W12998), .A2(I1576), .ZN(O18159));
  NANDX1 G20690 (.A1(W16977), .A2(W7411), .ZN(O18157));
  NANDX1 G20691 (.A1(W18575), .A2(W23273), .ZN(O18154));
  NANDX1 G20692 (.A1(W4776), .A2(W7948), .ZN(W49341));
  NANDX1 G20693 (.A1(W47559), .A2(W14154), .ZN(O18152));
  NANDX1 G20694 (.A1(W46079), .A2(W16781), .ZN(O18151));
  NANDX1 G20695 (.A1(W28588), .A2(W22745), .ZN(O18150));
  NANDX1 G20696 (.A1(W27217), .A2(W1751), .ZN(O18148));
  NANDX1 G20697 (.A1(W29913), .A2(W37245), .ZN(O18147));
  NANDX1 G20698 (.A1(W41673), .A2(W18487), .ZN(O18145));
  NANDX1 G20699 (.A1(W38230), .A2(W27100), .ZN(O18516));
  NANDX1 G20700 (.A1(W7271), .A2(W25541), .ZN(O18536));
  NANDX1 G20701 (.A1(W4595), .A2(W32970), .ZN(O18535));
  NANDX1 G20702 (.A1(W38370), .A2(W44007), .ZN(O18534));
  NANDX1 G20703 (.A1(W8268), .A2(W3789), .ZN(O18531));
  NANDX1 G20704 (.A1(W16098), .A2(W1862), .ZN(O18530));
  NANDX1 G20705 (.A1(W35478), .A2(W34530), .ZN(O18529));
  NANDX1 G20706 (.A1(W14644), .A2(W5769), .ZN(O18525));
  NANDX1 G20707 (.A1(W6021), .A2(W22596), .ZN(O18524));
  NANDX1 G20708 (.A1(W41856), .A2(W17816), .ZN(O18521));
  NANDX1 G20709 (.A1(W18850), .A2(W5582), .ZN(O18520));
  NANDX1 G20710 (.A1(I1014), .A2(W3807), .ZN(O18518));
  NANDX1 G20711 (.A1(W27027), .A2(W20098), .ZN(O18517));
  NANDX1 G20712 (.A1(W19383), .A2(W35602), .ZN(O18537));
  NANDX1 G20713 (.A1(W39484), .A2(W20993), .ZN(O18515));
  NANDX1 G20714 (.A1(W1591), .A2(W41930), .ZN(O18514));
  NANDX1 G20715 (.A1(W18460), .A2(W38025), .ZN(O18512));
  NANDX1 G20716 (.A1(W12648), .A2(W47565), .ZN(O18508));
  NANDX1 G20717 (.A1(W49379), .A2(W79), .ZN(O18500));
  NANDX1 G20718 (.A1(W46708), .A2(W22786), .ZN(O18498));
  NANDX1 G20719 (.A1(W48254), .A2(W15533), .ZN(O18497));
  NANDX1 G20720 (.A1(I1800), .A2(W46107), .ZN(O18495));
  NANDX1 G20721 (.A1(W2795), .A2(W28541), .ZN(W49687));
  NANDX1 G20722 (.A1(W1011), .A2(W11639), .ZN(O18477));
  NANDX1 G20723 (.A1(W13546), .A2(W33193), .ZN(O18476));
  NANDX1 G20724 (.A1(W48395), .A2(W33929), .ZN(O18596));
  NANDX1 G20725 (.A1(W32388), .A2(W17987), .ZN(O18618));
  NANDX1 G20726 (.A1(W21826), .A2(W24839), .ZN(O18617));
  NANDX1 G20727 (.A1(W31557), .A2(W41665), .ZN(O18614));
  NANDX1 G20728 (.A1(W26228), .A2(W3986), .ZN(O18613));
  NANDX1 G20729 (.A1(W3466), .A2(W22077), .ZN(O18611));
  NANDX1 G20730 (.A1(W34260), .A2(W30663), .ZN(O18609));
  NANDX1 G20731 (.A1(W21600), .A2(W28604), .ZN(O18608));
  NANDX1 G20732 (.A1(W44397), .A2(W33060), .ZN(W49816));
  NANDX1 G20733 (.A1(W31536), .A2(W18489), .ZN(O18601));
  NANDX1 G20734 (.A1(W17956), .A2(W4928), .ZN(O18600));
  NANDX1 G20735 (.A1(W37374), .A2(W18610), .ZN(O18599));
  NANDX1 G20736 (.A1(W16994), .A2(W8522), .ZN(O18597));
  NANDX1 G20737 (.A1(W38781), .A2(W14275), .ZN(O18475));
  NANDX1 G20738 (.A1(W14240), .A2(W42358), .ZN(O18589));
  NANDX1 G20739 (.A1(W21376), .A2(W24078), .ZN(O18588));
  NANDX1 G20740 (.A1(W2642), .A2(W7562), .ZN(O18575));
  NANDX1 G20741 (.A1(W3770), .A2(I417), .ZN(O18574));
  NANDX1 G20742 (.A1(W19647), .A2(W19497), .ZN(O18568));
  NANDX1 G20743 (.A1(W48231), .A2(W25461), .ZN(O18563));
  NANDX1 G20744 (.A1(W7968), .A2(W18231), .ZN(O18550));
  NANDX1 G20745 (.A1(W41216), .A2(W4247), .ZN(O18548));
  NANDX1 G20746 (.A1(W2765), .A2(W5589), .ZN(O18546));
  NANDX1 G20747 (.A1(W38540), .A2(W37016), .ZN(O18544));
  NANDX1 G20748 (.A1(W44542), .A2(W40134), .ZN(O18541));
  NANDX1 G20749 (.A1(W884), .A2(W37840), .ZN(O18374));
  NANDX1 G20750 (.A1(W45102), .A2(W40315), .ZN(O18415));
  NANDX1 G20751 (.A1(W39958), .A2(W4479), .ZN(O18414));
  NANDX1 G20752 (.A1(W15186), .A2(W42983), .ZN(O18411));
  NANDX1 G20753 (.A1(W25945), .A2(W27754), .ZN(O18409));
  NANDX1 G20754 (.A1(W25881), .A2(W28646), .ZN(O18405));
  NANDX1 G20755 (.A1(W10289), .A2(W46638), .ZN(O18404));
  NANDX1 G20756 (.A1(W35329), .A2(W24327), .ZN(O18390));
  NANDX1 G20757 (.A1(W8238), .A2(W9858), .ZN(O18389));
  NANDX1 G20758 (.A1(W44950), .A2(W30945), .ZN(O18388));
  NANDX1 G20759 (.A1(W41403), .A2(W28649), .ZN(O18384));
  NANDX1 G20760 (.A1(W46411), .A2(W3694), .ZN(O18380));
  NANDX1 G20761 (.A1(W19057), .A2(W46480), .ZN(O18376));
  NANDX1 G20762 (.A1(W26542), .A2(W33966), .ZN(O18417));
  NANDX1 G20763 (.A1(W6720), .A2(W47611), .ZN(W49570));
  NANDX1 G20764 (.A1(W4416), .A2(W32123), .ZN(O18366));
  NANDX1 G20765 (.A1(W47665), .A2(W44359), .ZN(O18365));
  NANDX1 G20766 (.A1(W29995), .A2(W15809), .ZN(O18359));
  NANDX1 G20767 (.A1(W27579), .A2(W21810), .ZN(O18358));
  NANDX1 G20768 (.A1(W43958), .A2(W48777), .ZN(O18357));
  NANDX1 G20769 (.A1(W563), .A2(W37837), .ZN(O18356));
  NANDX1 G20770 (.A1(W28175), .A2(W17200), .ZN(O18353));
  NANDX1 G20771 (.A1(W16198), .A2(W17458), .ZN(O18351));
  NANDX1 G20772 (.A1(W15045), .A2(W31559), .ZN(O18349));
  NANDX1 G20773 (.A1(W6459), .A2(W40048), .ZN(O18342));
  NANDX1 G20774 (.A1(W3657), .A2(W33590), .ZN(O18452));
  NANDX1 G20775 (.A1(W14548), .A2(W12187), .ZN(O18471));
  NANDX1 G20776 (.A1(W20899), .A2(W21207), .ZN(O18469));
  NANDX1 G20777 (.A1(W17937), .A2(W19762), .ZN(O18467));
  NANDX1 G20778 (.A1(W48803), .A2(W47993), .ZN(O18466));
  NANDX1 G20779 (.A1(W38281), .A2(W16961), .ZN(O18463));
  NANDX1 G20780 (.A1(W49634), .A2(I1146), .ZN(O18462));
  NANDX1 G20781 (.A1(W30856), .A2(W29654), .ZN(W49668));
  NANDX1 G20782 (.A1(W434), .A2(W49078), .ZN(O18458));
  NANDX1 G20783 (.A1(W31345), .A2(W731), .ZN(O18457));
  NANDX1 G20784 (.A1(W17848), .A2(W26930), .ZN(W49660));
  NANDX1 G20785 (.A1(W48976), .A2(W46029), .ZN(O18454));
  NANDX1 G20786 (.A1(W14858), .A2(W41154), .ZN(O18052));
  NANDX1 G20787 (.A1(W936), .A2(W34213), .ZN(O18450));
  NANDX1 G20788 (.A1(W3162), .A2(W19089), .ZN(O18448));
  NANDX1 G20789 (.A1(W19878), .A2(W47386), .ZN(O18440));
  NANDX1 G20790 (.A1(I1204), .A2(W41620), .ZN(O18435));
  NANDX1 G20791 (.A1(W41030), .A2(W39053), .ZN(O18430));
  NANDX1 G20792 (.A1(W26537), .A2(W3519), .ZN(W49634));
  NANDX1 G20793 (.A1(I410), .A2(W4163), .ZN(O18429));
  NANDX1 G20794 (.A1(W21286), .A2(W35023), .ZN(O18428));
  NANDX1 G20795 (.A1(W35160), .A2(W22073), .ZN(O18426));
  NANDX1 G20796 (.A1(W30492), .A2(W8551), .ZN(O18424));
  NANDX1 G20797 (.A1(W3350), .A2(W11187), .ZN(O18418));
  NANDX1 G20798 (.A1(W18419), .A2(W17890), .ZN(O17661));
  NANDX1 G20799 (.A1(W39968), .A2(W30197), .ZN(O17698));
  NANDX1 G20800 (.A1(W13985), .A2(W15483), .ZN(O17696));
  NANDX1 G20801 (.A1(W41463), .A2(W7168), .ZN(W48848));
  NANDX1 G20802 (.A1(W41198), .A2(W13132), .ZN(O17692));
  NANDX1 G20803 (.A1(W10696), .A2(W30684), .ZN(O17687));
  NANDX1 G20804 (.A1(W48145), .A2(W31443), .ZN(O17685));
  NANDX1 G20805 (.A1(W47158), .A2(W44150), .ZN(W48836));
  NANDX1 G20806 (.A1(W9147), .A2(W4053), .ZN(O17679));
  NANDX1 G20807 (.A1(W13150), .A2(W17208), .ZN(O17673));
  NANDX1 G20808 (.A1(W44742), .A2(W24812), .ZN(O17671));
  NANDX1 G20809 (.A1(W21880), .A2(I1848), .ZN(O17670));
  NANDX1 G20810 (.A1(W44989), .A2(W39279), .ZN(O17665));
  NANDX1 G20811 (.A1(W21401), .A2(W12034), .ZN(O17706));
  NANDX1 G20812 (.A1(W7219), .A2(W30151), .ZN(O17655));
  NANDX1 G20813 (.A1(W19424), .A2(W43917), .ZN(W48803));
  NANDX1 G20814 (.A1(W23856), .A2(W5634), .ZN(O17651));
  NANDX1 G20815 (.A1(W32568), .A2(W37763), .ZN(W48790));
  NANDX1 G20816 (.A1(W34127), .A2(W675), .ZN(O17638));
  NANDX1 G20817 (.A1(W12593), .A2(W30167), .ZN(O17636));
  NANDX1 G20818 (.A1(W48670), .A2(W17511), .ZN(O17635));
  NANDX1 G20819 (.A1(W28453), .A2(W45821), .ZN(O17634));
  NANDX1 G20820 (.A1(W21754), .A2(W29922), .ZN(W48777));
  NANDX1 G20821 (.A1(W178), .A2(W24467), .ZN(O17630));
  NANDX1 G20822 (.A1(W27293), .A2(W20923), .ZN(O17626));
  NANDX1 G20823 (.A1(W1829), .A2(W46776), .ZN(O17752));
  NANDX1 G20824 (.A1(W18425), .A2(W11867), .ZN(O17777));
  NANDX1 G20825 (.A1(W46641), .A2(W261), .ZN(W48936));
  NANDX1 G20826 (.A1(W39312), .A2(W8079), .ZN(O17769));
  NANDX1 G20827 (.A1(W26082), .A2(W16845), .ZN(O17766));
  NANDX1 G20828 (.A1(W15473), .A2(W24732), .ZN(O17765));
  NANDX1 G20829 (.A1(W32289), .A2(W38369), .ZN(O17763));
  NANDX1 G20830 (.A1(W41678), .A2(W17086), .ZN(O17760));
  NANDX1 G20831 (.A1(W1583), .A2(W8347), .ZN(W48915));
  NANDX1 G20832 (.A1(W23233), .A2(W27476), .ZN(O17756));
  NANDX1 G20833 (.A1(I635), .A2(W22048), .ZN(O17755));
  NANDX1 G20834 (.A1(W35491), .A2(W1877), .ZN(O17754));
  NANDX1 G20835 (.A1(W14491), .A2(W48602), .ZN(O17753));
  NANDX1 G20836 (.A1(W27795), .A2(W17982), .ZN(O17618));
  NANDX1 G20837 (.A1(W37514), .A2(W12682), .ZN(W48908));
  NANDX1 G20838 (.A1(W39666), .A2(W12756), .ZN(O17747));
  NANDX1 G20839 (.A1(I492), .A2(W19793), .ZN(O17745));
  NANDX1 G20840 (.A1(W11501), .A2(W48775), .ZN(W48899));
  NANDX1 G20841 (.A1(W26194), .A2(W6446), .ZN(O17741));
  NANDX1 G20842 (.A1(W2024), .A2(W45858), .ZN(O17736));
  NANDX1 G20843 (.A1(W7624), .A2(W33383), .ZN(O17729));
  NANDX1 G20844 (.A1(W37233), .A2(W45296), .ZN(O17727));
  NANDX1 G20845 (.A1(W36309), .A2(W5058), .ZN(O17725));
  NANDX1 G20846 (.A1(W31176), .A2(W46848), .ZN(O17719));
  NANDX1 G20847 (.A1(W18862), .A2(W9355), .ZN(O17715));
  NANDX1 G20848 (.A1(W11526), .A2(W41383), .ZN(O17528));
  NANDX1 G20849 (.A1(I435), .A2(W44922), .ZN(O17553));
  NANDX1 G20850 (.A1(W36911), .A2(W16531), .ZN(O17551));
  NANDX1 G20851 (.A1(W32365), .A2(W40575), .ZN(O17549));
  NANDX1 G20852 (.A1(W31311), .A2(W43203), .ZN(O17548));
  NANDX1 G20853 (.A1(W7029), .A2(W5633), .ZN(O17545));
  NANDX1 G20854 (.A1(W21048), .A2(W9920), .ZN(O17543));
  NANDX1 G20855 (.A1(I1769), .A2(W39816), .ZN(O17542));
  NANDX1 G20856 (.A1(W18630), .A2(W2562), .ZN(O17541));
  NANDX1 G20857 (.A1(W31142), .A2(W46378), .ZN(O17537));
  NANDX1 G20858 (.A1(W37524), .A2(W35065), .ZN(O17535));
  NANDX1 G20859 (.A1(W38675), .A2(W32919), .ZN(W48669));
  NANDX1 G20860 (.A1(W42450), .A2(W8869), .ZN(W48664));
  NANDX1 G20861 (.A1(W8799), .A2(W23201), .ZN(O17554));
  NANDX1 G20862 (.A1(W28760), .A2(W39736), .ZN(O17527));
  NANDX1 G20863 (.A1(W28471), .A2(W2385), .ZN(O17523));
  NANDX1 G20864 (.A1(W30857), .A2(W1967), .ZN(O17522));
  NANDX1 G20865 (.A1(W48148), .A2(W4287), .ZN(O17519));
  NANDX1 G20866 (.A1(W18158), .A2(W38055), .ZN(O17514));
  NANDX1 G20867 (.A1(W37966), .A2(W3110), .ZN(O17505));
  NANDX1 G20868 (.A1(W32101), .A2(W36867), .ZN(O17500));
  NANDX1 G20869 (.A1(W27733), .A2(W3605), .ZN(O17499));
  NANDX1 G20870 (.A1(W46415), .A2(W7399), .ZN(O17497));
  NANDX1 G20871 (.A1(W41577), .A2(W17841), .ZN(O17496));
  NANDX1 G20872 (.A1(W33087), .A2(W26243), .ZN(O17491));
  NANDX1 G20873 (.A1(W30164), .A2(W11877), .ZN(O17584));
  NANDX1 G20874 (.A1(W23350), .A2(W26376), .ZN(O17615));
  NANDX1 G20875 (.A1(W29189), .A2(W12770), .ZN(O17613));
  NANDX1 G20876 (.A1(W47278), .A2(W9741), .ZN(O17609));
  NANDX1 G20877 (.A1(W10522), .A2(W10373), .ZN(O17608));
  NANDX1 G20878 (.A1(W7778), .A2(W28174), .ZN(O17607));
  NANDX1 G20879 (.A1(I1903), .A2(W27239), .ZN(O17603));
  NANDX1 G20880 (.A1(W33624), .A2(W4018), .ZN(O17601));
  NANDX1 G20881 (.A1(W17591), .A2(W42106), .ZN(W48739));
  NANDX1 G20882 (.A1(W14058), .A2(W20949), .ZN(O17592));
  NANDX1 G20883 (.A1(W16729), .A2(W8023), .ZN(O17588));
  NANDX1 G20884 (.A1(W18858), .A2(W37738), .ZN(O17587));
  NANDX1 G20885 (.A1(W18691), .A2(W18104), .ZN(O17778));
  NANDX1 G20886 (.A1(W21036), .A2(W27009), .ZN(O17582));
  NANDX1 G20887 (.A1(W32984), .A2(W2399), .ZN(O17581));
  NANDX1 G20888 (.A1(W18897), .A2(W5263), .ZN(W48717));
  NANDX1 G20889 (.A1(W21620), .A2(W16121), .ZN(O17575));
  NANDX1 G20890 (.A1(W20337), .A2(W23758), .ZN(O17574));
  NANDX1 G20891 (.A1(W37464), .A2(W48114), .ZN(O17573));
  NANDX1 G20892 (.A1(W23465), .A2(W28751), .ZN(O17571));
  NANDX1 G20893 (.A1(W17498), .A2(W44159), .ZN(W48706));
  NANDX1 G20894 (.A1(W24408), .A2(W4658), .ZN(O17561));
  NANDX1 G20895 (.A1(W41694), .A2(W6292), .ZN(W48695));
  NANDX1 G20896 (.A1(W27934), .A2(W15431), .ZN(O17556));
  NANDX1 G20897 (.A1(W6548), .A2(W37460), .ZN(O17939));
  NANDX1 G20898 (.A1(W27867), .A2(W46733), .ZN(O17979));
  NANDX1 G20899 (.A1(W43757), .A2(W32485), .ZN(O17978));
  NANDX1 G20900 (.A1(W17163), .A2(W47266), .ZN(O17975));
  NANDX1 G20901 (.A1(W46531), .A2(W43398), .ZN(O17972));
  NANDX1 G20902 (.A1(W39460), .A2(W33855), .ZN(O17963));
  NANDX1 G20903 (.A1(W23036), .A2(W15406), .ZN(O17962));
  NANDX1 G20904 (.A1(W30120), .A2(I142), .ZN(O17958));
  NANDX1 G20905 (.A1(W40674), .A2(W18175), .ZN(O17954));
  NANDX1 G20906 (.A1(W2525), .A2(W5168), .ZN(O17953));
  NANDX1 G20907 (.A1(W30207), .A2(W8253), .ZN(O17950));
  NANDX1 G20908 (.A1(W36162), .A2(W8416), .ZN(O17946));
  NANDX1 G20909 (.A1(W39403), .A2(W4214), .ZN(O17944));
  NANDX1 G20910 (.A1(W43695), .A2(W46512), .ZN(O17984));
  NANDX1 G20911 (.A1(W10698), .A2(W41022), .ZN(O17937));
  NANDX1 G20912 (.A1(W42605), .A2(W47404), .ZN(O17933));
  NANDX1 G20913 (.A1(W33151), .A2(W10913), .ZN(O17932));
  NANDX1 G20914 (.A1(W17340), .A2(W19148), .ZN(O17931));
  NANDX1 G20915 (.A1(W7617), .A2(W34589), .ZN(O17928));
  NANDX1 G20916 (.A1(W40799), .A2(W23357), .ZN(O17926));
  NANDX1 G20917 (.A1(W839), .A2(W26707), .ZN(O17922));
  NANDX1 G20918 (.A1(W35019), .A2(W19034), .ZN(O17920));
  NANDX1 G20919 (.A1(W4881), .A2(W13708), .ZN(O17919));
  NANDX1 G20920 (.A1(W12969), .A2(W11297), .ZN(W49087));
  NANDX1 G20921 (.A1(W20125), .A2(W30743), .ZN(W49086));
  NANDX1 G20922 (.A1(W38689), .A2(W9396), .ZN(O18016));
  NANDX1 G20923 (.A1(W6615), .A2(W44999), .ZN(W49234));
  NANDX1 G20924 (.A1(W46860), .A2(W38951), .ZN(O18051));
  NANDX1 G20925 (.A1(W33364), .A2(W45364), .ZN(O18049));
  NANDX1 G20926 (.A1(W36347), .A2(W27074), .ZN(O18048));
  NANDX1 G20927 (.A1(W44864), .A2(I128), .ZN(O18038));
  NANDX1 G20928 (.A1(W44364), .A2(W29056), .ZN(O18037));
  NANDX1 G20929 (.A1(W7622), .A2(W3646), .ZN(O18036));
  NANDX1 G20930 (.A1(W29171), .A2(W33485), .ZN(O18034));
  NANDX1 G20931 (.A1(W22926), .A2(W29417), .ZN(O18032));
  NANDX1 G20932 (.A1(W634), .A2(W22561), .ZN(O18026));
  NANDX1 G20933 (.A1(W46769), .A2(W46313), .ZN(O18025));
  NANDX1 G20934 (.A1(W24378), .A2(W5973), .ZN(O18023));
  NANDX1 G20935 (.A1(W36299), .A2(W28129), .ZN(O17913));
  NANDX1 G20936 (.A1(W40881), .A2(W1945), .ZN(O18015));
  NANDX1 G20937 (.A1(W42019), .A2(W45922), .ZN(O18014));
  NANDX1 G20938 (.A1(W2512), .A2(W26299), .ZN(W49190));
  NANDX1 G20939 (.A1(W45533), .A2(W18994), .ZN(O18003));
  NANDX1 G20940 (.A1(W27982), .A2(W37294), .ZN(O18001));
  NANDX1 G20941 (.A1(W19750), .A2(W47516), .ZN(O17999));
  NANDX1 G20942 (.A1(W13907), .A2(I878), .ZN(O17997));
  NANDX1 G20943 (.A1(W14148), .A2(W47854), .ZN(O17996));
  NANDX1 G20944 (.A1(W18103), .A2(W15505), .ZN(O17993));
  NANDX1 G20945 (.A1(W20149), .A2(W10081), .ZN(O17992));
  NANDX1 G20946 (.A1(W29731), .A2(W5638), .ZN(O17989));
  NANDX1 G20947 (.A1(W30133), .A2(W2775), .ZN(O17812));
  NANDX1 G20948 (.A1(W42838), .A2(W37081), .ZN(O17858));
  NANDX1 G20949 (.A1(W41804), .A2(W5469), .ZN(O17853));
  NANDX1 G20950 (.A1(W12776), .A2(W46786), .ZN(O17851));
  NANDX1 G20951 (.A1(I503), .A2(W3774), .ZN(O17846));
  NANDX1 G20952 (.A1(W1365), .A2(W10116), .ZN(O17842));
  NANDX1 G20953 (.A1(W42300), .A2(W29723), .ZN(O17839));
  NANDX1 G20954 (.A1(W9073), .A2(W27775), .ZN(O17836));
  NANDX1 G20955 (.A1(W9242), .A2(W25755), .ZN(O17828));
  NANDX1 G20956 (.A1(W24200), .A2(W20752), .ZN(O17821));
  NANDX1 G20957 (.A1(W3824), .A2(W16407), .ZN(O17818));
  NANDX1 G20958 (.A1(W48459), .A2(W37736), .ZN(O17817));
  NANDX1 G20959 (.A1(W27528), .A2(W18416), .ZN(O17816));
  NANDX1 G20960 (.A1(W10599), .A2(W41473), .ZN(O17862));
  NANDX1 G20961 (.A1(W24042), .A2(W697), .ZN(O17808));
  NANDX1 G20962 (.A1(W5124), .A2(W29362), .ZN(O17806));
  NANDX1 G20963 (.A1(W16010), .A2(W35341), .ZN(O17804));
  NANDX1 G20964 (.A1(W22452), .A2(W36067), .ZN(O17802));
  NANDX1 G20965 (.A1(W21445), .A2(W21601), .ZN(W48963));
  NANDX1 G20966 (.A1(W4178), .A2(W7581), .ZN(O17801));
  NANDX1 G20967 (.A1(W11506), .A2(W37256), .ZN(O17800));
  NANDX1 G20968 (.A1(W13586), .A2(W30424), .ZN(W48958));
  NANDX1 G20969 (.A1(W21389), .A2(W18701), .ZN(O17791));
  NANDX1 G20970 (.A1(W9162), .A2(W40696), .ZN(O17788));
  NANDX1 G20971 (.A1(W13933), .A2(W19188), .ZN(O17780));
  NANDX1 G20972 (.A1(W44775), .A2(W33748), .ZN(O17892));
  NANDX1 G20973 (.A1(W40267), .A2(W7564), .ZN(O17912));
  NANDX1 G20974 (.A1(W44086), .A2(W32345), .ZN(O17911));
  NANDX1 G20975 (.A1(W34952), .A2(W10317), .ZN(O17910));
  NANDX1 G20976 (.A1(W23196), .A2(W12846), .ZN(O17909));
  NANDX1 G20977 (.A1(W40712), .A2(W44092), .ZN(O17907));
  NANDX1 G20978 (.A1(W28886), .A2(W20526), .ZN(O17906));
  NANDX1 G20979 (.A1(W10459), .A2(W7981), .ZN(O17905));
  NANDX1 G20980 (.A1(W43864), .A2(W44388), .ZN(O17902));
  NANDX1 G20981 (.A1(W16855), .A2(W20723), .ZN(O17901));
  NANDX1 G20982 (.A1(W35782), .A2(W37023), .ZN(O17900));
  NANDX1 G20983 (.A1(W46812), .A2(W3585), .ZN(W49068));
  NANDX1 G20984 (.A1(W19293), .A2(W33308), .ZN(W49839));
  NANDX1 G20985 (.A1(W45322), .A2(W16293), .ZN(O17889));
  NANDX1 G20986 (.A1(W41009), .A2(W43746), .ZN(O17888));
  NANDX1 G20987 (.A1(W24897), .A2(W4126), .ZN(O17887));
  NANDX1 G20988 (.A1(W12746), .A2(W25440), .ZN(O17886));
  NANDX1 G20989 (.A1(W15776), .A2(W21071), .ZN(O17881));
  NANDX1 G20990 (.A1(I269), .A2(W42228), .ZN(O17880));
  NANDX1 G20991 (.A1(W46227), .A2(W16603), .ZN(O17875));
  NANDX1 G20992 (.A1(W4027), .A2(W48540), .ZN(O17874));
  NANDX1 G20993 (.A1(W37822), .A2(W18916), .ZN(O17871));
  NANDX1 G20994 (.A1(W20865), .A2(W36142), .ZN(O17867));
  NANDX1 G20995 (.A1(W46999), .A2(W46764), .ZN(O17865));
  NANDX1 G20996 (.A1(W7968), .A2(W34206), .ZN(O19354));
  NANDX1 G20997 (.A1(W43093), .A2(W10208), .ZN(O19388));
  NANDX1 G20998 (.A1(W43119), .A2(W21642), .ZN(O19385));
  NANDX1 G20999 (.A1(W40990), .A2(W22351), .ZN(O19382));
  NANDX1 G21000 (.A1(W34948), .A2(W50072), .ZN(O19378));
  NANDX1 G21001 (.A1(W14236), .A2(I366), .ZN(O19374));
  NANDX1 G21002 (.A1(W21141), .A2(W46707), .ZN(O19372));
  NANDX1 G21003 (.A1(W3338), .A2(W30070), .ZN(O19367));
  NANDX1 G21004 (.A1(W5823), .A2(W9034), .ZN(O19365));
  NANDX1 G21005 (.A1(W39042), .A2(W32755), .ZN(O19363));
  NANDX1 G21006 (.A1(W30733), .A2(W13870), .ZN(O19359));
  NANDX1 G21007 (.A1(W40875), .A2(W10575), .ZN(O19358));
  NANDX1 G21008 (.A1(W16347), .A2(W10924), .ZN(O19357));
  NANDX1 G21009 (.A1(W37541), .A2(W38043), .ZN(O19392));
  NANDX1 G21010 (.A1(W1208), .A2(W1520), .ZN(O19351));
  NANDX1 G21011 (.A1(W19419), .A2(W5946), .ZN(O19350));
  NANDX1 G21012 (.A1(W24557), .A2(W9598), .ZN(O19349));
  NANDX1 G21013 (.A1(W49368), .A2(W44993), .ZN(O19348));
  NANDX1 G21014 (.A1(W8208), .A2(W8978), .ZN(O19347));
  NANDX1 G21015 (.A1(W2693), .A2(W1910), .ZN(O19341));
  NANDX1 G21016 (.A1(W993), .A2(W26675), .ZN(W50563));
  NANDX1 G21017 (.A1(W26879), .A2(W44990), .ZN(O19324));
  NANDX1 G21018 (.A1(W45264), .A2(W42033), .ZN(O19323));
  NANDX1 G21019 (.A1(W41454), .A2(W16083), .ZN(O19322));
  NANDX1 G21020 (.A1(W41104), .A2(W2025), .ZN(O19318));
  NANDX1 G21021 (.A1(W47296), .A2(W12708), .ZN(O19423));
  NANDX1 G21022 (.A1(W33515), .A2(W38752), .ZN(O19478));
  NANDX1 G21023 (.A1(W36640), .A2(W17391), .ZN(O19473));
  NANDX1 G21024 (.A1(W50410), .A2(W22988), .ZN(O19472));
  NANDX1 G21025 (.A1(W32504), .A2(W12083), .ZN(O19470));
  NANDX1 G21026 (.A1(W2290), .A2(W37099), .ZN(O19460));
  NANDX1 G21027 (.A1(W36144), .A2(W2875), .ZN(O19458));
  NANDX1 G21028 (.A1(W39427), .A2(W26987), .ZN(O19450));
  NANDX1 G21029 (.A1(W12991), .A2(W42857), .ZN(O19444));
  NANDX1 G21030 (.A1(W34481), .A2(W19250), .ZN(O19439));
  NANDX1 G21031 (.A1(W9985), .A2(W9492), .ZN(O19436));
  NANDX1 G21032 (.A1(W14357), .A2(W34858), .ZN(O19430));
  NANDX1 G21033 (.A1(W36021), .A2(W33714), .ZN(O19426));
  NANDX1 G21034 (.A1(W41076), .A2(W14317), .ZN(O19316));
  NANDX1 G21035 (.A1(W41380), .A2(I764), .ZN(O19421));
  NANDX1 G21036 (.A1(W50250), .A2(W11748), .ZN(O19420));
  NANDX1 G21037 (.A1(W14961), .A2(W18667), .ZN(O19416));
  NANDX1 G21038 (.A1(W43756), .A2(W829), .ZN(O19414));
  NANDX1 G21039 (.A1(W20400), .A2(W44391), .ZN(O19413));
  NANDX1 G21040 (.A1(W2171), .A2(W16836), .ZN(O19412));
  NANDX1 G21041 (.A1(W13630), .A2(W20669), .ZN(O19411));
  NANDX1 G21042 (.A1(W15729), .A2(W32129), .ZN(O19407));
  NANDX1 G21043 (.A1(W49433), .A2(W26414), .ZN(O19404));
  NANDX1 G21044 (.A1(W19681), .A2(W38798), .ZN(O19400));
  NANDX1 G21045 (.A1(W5344), .A2(W45288), .ZN(O19396));
  NANDX1 G21046 (.A1(W8051), .A2(W20988), .ZN(O19199));
  NANDX1 G21047 (.A1(W24910), .A2(W28129), .ZN(O19235));
  NANDX1 G21048 (.A1(W19593), .A2(W15119), .ZN(O19230));
  NANDX1 G21049 (.A1(W9149), .A2(W28164), .ZN(O19228));
  NANDX1 G21050 (.A1(W6816), .A2(W49037), .ZN(O19224));
  NANDX1 G21051 (.A1(W35617), .A2(W28999), .ZN(O19220));
  NANDX1 G21052 (.A1(W24554), .A2(W41446), .ZN(O19218));
  NANDX1 G21053 (.A1(I65), .A2(W33083), .ZN(O19213));
  NANDX1 G21054 (.A1(W7820), .A2(W16249), .ZN(O19210));
  NANDX1 G21055 (.A1(W2138), .A2(W10237), .ZN(O19207));
  NANDX1 G21056 (.A1(W25902), .A2(W39394), .ZN(O19206));
  NANDX1 G21057 (.A1(W28010), .A2(W22284), .ZN(O19204));
  NANDX1 G21058 (.A1(W49175), .A2(W5467), .ZN(O19200));
  NANDX1 G21059 (.A1(W311), .A2(W42245), .ZN(O19236));
  NANDX1 G21060 (.A1(W12814), .A2(W3647), .ZN(O19198));
  NANDX1 G21061 (.A1(W16352), .A2(W12554), .ZN(O19191));
  NANDX1 G21062 (.A1(W11071), .A2(W28631), .ZN(O19186));
  NANDX1 G21063 (.A1(W49133), .A2(W27252), .ZN(O19180));
  NANDX1 G21064 (.A1(W6956), .A2(W11776), .ZN(O19178));
  NANDX1 G21065 (.A1(W49448), .A2(W5075), .ZN(O19177));
  NANDX1 G21066 (.A1(W13488), .A2(W49018), .ZN(O19176));
  NANDX1 G21067 (.A1(W46681), .A2(W39036), .ZN(O19175));
  NANDX1 G21068 (.A1(W11205), .A2(W32939), .ZN(O19173));
  NANDX1 G21069 (.A1(W45314), .A2(W17429), .ZN(O19172));
  NANDX1 G21070 (.A1(W14828), .A2(W3531), .ZN(O19166));
  NANDX1 G21071 (.A1(W5063), .A2(W15028), .ZN(O19277));
  NANDX1 G21072 (.A1(W29940), .A2(W8104), .ZN(O19312));
  NANDX1 G21073 (.A1(I1651), .A2(W12168), .ZN(W50539));
  NANDX1 G21074 (.A1(W39476), .A2(W27681), .ZN(O19304));
  NANDX1 G21075 (.A1(W45025), .A2(W28174), .ZN(O19302));
  NANDX1 G21076 (.A1(W44083), .A2(W7536), .ZN(O19301));
  NANDX1 G21077 (.A1(W25233), .A2(W27788), .ZN(O19299));
  NANDX1 G21078 (.A1(W27395), .A2(W674), .ZN(O19295));
  NANDX1 G21079 (.A1(W41359), .A2(W32615), .ZN(O19288));
  NANDX1 G21080 (.A1(W18097), .A2(W24144), .ZN(O19287));
  NANDX1 G21081 (.A1(W43547), .A2(W36645), .ZN(O19286));
  NANDX1 G21082 (.A1(W5370), .A2(W29622), .ZN(O19280));
  NANDX1 G21083 (.A1(W48207), .A2(W23784), .ZN(O19479));
  NANDX1 G21084 (.A1(W40816), .A2(W22948), .ZN(O19275));
  NANDX1 G21085 (.A1(W46094), .A2(W32153), .ZN(O19272));
  NANDX1 G21086 (.A1(W35798), .A2(W46509), .ZN(O19268));
  NANDX1 G21087 (.A1(W4240), .A2(W4304), .ZN(O19257));
  NANDX1 G21088 (.A1(W34143), .A2(W391), .ZN(O19256));
  NANDX1 G21089 (.A1(W36187), .A2(W45409), .ZN(O19250));
  NANDX1 G21090 (.A1(W867), .A2(W8372), .ZN(O19249));
  NANDX1 G21091 (.A1(W31831), .A2(W17959), .ZN(O19244));
  NANDX1 G21092 (.A1(W7786), .A2(W747), .ZN(O19242));
  NANDX1 G21093 (.A1(W4086), .A2(W20561), .ZN(O19240));
  NANDX1 G21094 (.A1(W121), .A2(W22370), .ZN(O19237));
  NANDX1 G21095 (.A1(W6625), .A2(W13543), .ZN(O19633));
  NANDX1 G21096 (.A1(I1011), .A2(W18747), .ZN(O19672));
  NANDX1 G21097 (.A1(I541), .A2(W27817), .ZN(O19669));
  NANDX1 G21098 (.A1(W9698), .A2(W20321), .ZN(O19667));
  NANDX1 G21099 (.A1(W19638), .A2(W23318), .ZN(O19664));
  NANDX1 G21100 (.A1(W47414), .A2(W8622), .ZN(O19658));
  NANDX1 G21101 (.A1(W8006), .A2(W35435), .ZN(O19655));
  NANDX1 G21102 (.A1(W22260), .A2(W50563), .ZN(O19653));
  NANDX1 G21103 (.A1(W26059), .A2(W22717), .ZN(O19647));
  NANDX1 G21104 (.A1(W21897), .A2(W6190), .ZN(O19645));
  NANDX1 G21105 (.A1(W30697), .A2(W13681), .ZN(O19639));
  NANDX1 G21106 (.A1(W15941), .A2(W26647), .ZN(O19636));
  NANDX1 G21107 (.A1(W36704), .A2(W26203), .ZN(O19634));
  NANDX1 G21108 (.A1(W11777), .A2(W36558), .ZN(O19676));
  NANDX1 G21109 (.A1(W6135), .A2(W17336), .ZN(O19630));
  NANDX1 G21110 (.A1(W28873), .A2(W12280), .ZN(O19625));
  NANDX1 G21111 (.A1(W23080), .A2(W45951), .ZN(O19624));
  NANDX1 G21112 (.A1(W37599), .A2(W11506), .ZN(O19623));
  NANDX1 G21113 (.A1(W23533), .A2(W39208), .ZN(O19622));
  NANDX1 G21114 (.A1(W45008), .A2(W49715), .ZN(O19617));
  NANDX1 G21115 (.A1(W35745), .A2(W12745), .ZN(O19616));
  NANDX1 G21116 (.A1(W19411), .A2(W19352), .ZN(O19606));
  NANDX1 G21117 (.A1(W16977), .A2(W48523), .ZN(O19604));
  NANDX1 G21118 (.A1(W40720), .A2(W31676), .ZN(O19603));
  NANDX1 G21119 (.A1(W16689), .A2(W11094), .ZN(O19598));
  NANDX1 G21120 (.A1(W21461), .A2(W33422), .ZN(O19730));
  NANDX1 G21121 (.A1(W3948), .A2(W11293), .ZN(O19760));
  NANDX1 G21122 (.A1(W49055), .A2(W49527), .ZN(O19758));
  NANDX1 G21123 (.A1(W40185), .A2(W16423), .ZN(O19757));
  NANDX1 G21124 (.A1(W22537), .A2(W50909), .ZN(O19751));
  NANDX1 G21125 (.A1(W5417), .A2(W37968), .ZN(O19745));
  NANDX1 G21126 (.A1(W25870), .A2(W4221), .ZN(O19744));
  NANDX1 G21127 (.A1(W22538), .A2(I987), .ZN(O19743));
  NANDX1 G21128 (.A1(W26535), .A2(W20377), .ZN(O19741));
  NANDX1 G21129 (.A1(W12961), .A2(W25210), .ZN(O19740));
  NANDX1 G21130 (.A1(W627), .A2(W12687), .ZN(O19739));
  NANDX1 G21131 (.A1(W26498), .A2(W42109), .ZN(O19734));
  NANDX1 G21132 (.A1(W48283), .A2(W25354), .ZN(O19732));
  NANDX1 G21133 (.A1(W40889), .A2(W8793), .ZN(O19597));
  NANDX1 G21134 (.A1(W25667), .A2(W43389), .ZN(O19727));
  NANDX1 G21135 (.A1(W42738), .A2(W12170), .ZN(O19717));
  NANDX1 G21136 (.A1(W16354), .A2(W36509), .ZN(O19711));
  NANDX1 G21137 (.A1(W47539), .A2(W40349), .ZN(O19709));
  NANDX1 G21138 (.A1(W6216), .A2(W30861), .ZN(O19701));
  NANDX1 G21139 (.A1(W8863), .A2(W19154), .ZN(O19698));
  NANDX1 G21140 (.A1(W43431), .A2(W14677), .ZN(O19697));
  NANDX1 G21141 (.A1(W9422), .A2(W8277), .ZN(O19690));
  NANDX1 G21142 (.A1(W12079), .A2(W21154), .ZN(O19686));
  NANDX1 G21143 (.A1(W13758), .A2(W24951), .ZN(O19685));
  NANDX1 G21144 (.A1(W17117), .A2(W22112), .ZN(O19677));
  NANDX1 G21145 (.A1(W30124), .A2(W50116), .ZN(O19506));
  NANDX1 G21146 (.A1(W13870), .A2(W28247), .ZN(O19547));
  NANDX1 G21147 (.A1(W26924), .A2(W40788), .ZN(O19545));
  NANDX1 G21148 (.A1(W38141), .A2(W40304), .ZN(O19544));
  NANDX1 G21149 (.A1(W50698), .A2(W38605), .ZN(O19542));
  NANDX1 G21150 (.A1(W33617), .A2(W15506), .ZN(O19537));
  NANDX1 G21151 (.A1(W41298), .A2(W15971), .ZN(O19535));
  NANDX1 G21152 (.A1(W16474), .A2(W26493), .ZN(O19532));
  NANDX1 G21153 (.A1(W29146), .A2(W18055), .ZN(O19525));
  NANDX1 G21154 (.A1(W37445), .A2(W47613), .ZN(O19522));
  NANDX1 G21155 (.A1(W42302), .A2(W36199), .ZN(O19519));
  NANDX1 G21156 (.A1(W46836), .A2(W40936), .ZN(O19509));
  NANDX1 G21157 (.A1(W34726), .A2(W44863), .ZN(O19508));
  NANDX1 G21158 (.A1(W37251), .A2(W33791), .ZN(O19548));
  NANDX1 G21159 (.A1(W48160), .A2(W9963), .ZN(O19504));
  NANDX1 G21160 (.A1(W45086), .A2(W35158), .ZN(O19503));
  NANDX1 G21161 (.A1(W14716), .A2(W48147), .ZN(O19501));
  NANDX1 G21162 (.A1(W13023), .A2(I466), .ZN(O19497));
  NANDX1 G21163 (.A1(W18476), .A2(W34157), .ZN(O19495));
  NANDX1 G21164 (.A1(W34900), .A2(W9022), .ZN(O19494));
  NANDX1 G21165 (.A1(W2776), .A2(W47529), .ZN(O19492));
  NANDX1 G21166 (.A1(W46425), .A2(W19600), .ZN(O19489));
  NANDX1 G21167 (.A1(W44922), .A2(W7413), .ZN(O19487));
  NANDX1 G21168 (.A1(W35829), .A2(W8322), .ZN(O19486));
  NANDX1 G21169 (.A1(W27540), .A2(W7887), .ZN(O19481));
  NANDX1 G21170 (.A1(W23536), .A2(W2654), .ZN(O19580));
  NANDX1 G21171 (.A1(W24974), .A2(W23649), .ZN(O19596));
  NANDX1 G21172 (.A1(W36451), .A2(W11505), .ZN(O19595));
  NANDX1 G21173 (.A1(W37925), .A2(W1623), .ZN(O19593));
  NANDX1 G21174 (.A1(W45580), .A2(W4005), .ZN(O19591));
  NANDX1 G21175 (.A1(W48828), .A2(W14001), .ZN(O19590));
  NANDX1 G21176 (.A1(W21603), .A2(W19739), .ZN(O19588));
  NANDX1 G21177 (.A1(W3171), .A2(W20484), .ZN(O19587));
  NANDX1 G21178 (.A1(W14650), .A2(W48908), .ZN(O19586));
  NANDX1 G21179 (.A1(W21107), .A2(W1293), .ZN(O19585));
  NANDX1 G21180 (.A1(W17935), .A2(W20008), .ZN(O19582));
  NANDX1 G21181 (.A1(W16506), .A2(W4412), .ZN(O19581));
  NANDX1 G21182 (.A1(W29432), .A2(W16305), .ZN(O19163));
  NANDX1 G21183 (.A1(W35814), .A2(W11316), .ZN(O19577));
  NANDX1 G21184 (.A1(W8126), .A2(W8697), .ZN(O19573));
  NANDX1 G21185 (.A1(W1581), .A2(W14391), .ZN(O19570));
  NANDX1 G21186 (.A1(W40526), .A2(W19715), .ZN(O19569));
  NANDX1 G21187 (.A1(W43668), .A2(W25768), .ZN(O19566));
  NANDX1 G21188 (.A1(W189), .A2(W1707), .ZN(O19565));
  NANDX1 G21189 (.A1(W3648), .A2(W4070), .ZN(O19564));
  NANDX1 G21190 (.A1(W33759), .A2(W50445), .ZN(O19561));
  NANDX1 G21191 (.A1(W44763), .A2(W11753), .ZN(O19556));
  NANDX1 G21192 (.A1(W4359), .A2(W6507), .ZN(O19553));
  NANDX1 G21193 (.A1(W33137), .A2(W3917), .ZN(O19549));
  NANDX1 G21194 (.A1(W14441), .A2(W28872), .ZN(O18800));
  NANDX1 G21195 (.A1(W23504), .A2(W11403), .ZN(O18829));
  NANDX1 G21196 (.A1(I17), .A2(W14675), .ZN(O18824));
  NANDX1 G21197 (.A1(W42979), .A2(I990), .ZN(O18822));
  NANDX1 G21198 (.A1(W1401), .A2(W33018), .ZN(O18821));
  NANDX1 G21199 (.A1(W13923), .A2(I1357), .ZN(O18820));
  NANDX1 G21200 (.A1(W43657), .A2(W21525), .ZN(O18815));
  NANDX1 G21201 (.A1(W17504), .A2(W48872), .ZN(O18814));
  NANDX1 G21202 (.A1(W33848), .A2(W9751), .ZN(O18812));
  NANDX1 G21203 (.A1(W12313), .A2(W31461), .ZN(O18809));
  NANDX1 G21204 (.A1(W7008), .A2(W11407), .ZN(O18808));
  NANDX1 G21205 (.A1(W37413), .A2(W962), .ZN(O18807));
  NANDX1 G21206 (.A1(W16670), .A2(W46082), .ZN(O18802));
  NANDX1 G21207 (.A1(W22041), .A2(W750), .ZN(O18830));
  NANDX1 G21208 (.A1(W47822), .A2(I1514), .ZN(O18799));
  NANDX1 G21209 (.A1(W4311), .A2(W21014), .ZN(O18796));
  NANDX1 G21210 (.A1(W11866), .A2(I1568), .ZN(O18794));
  NANDX1 G21211 (.A1(W42890), .A2(W28104), .ZN(O18785));
  NANDX1 G21212 (.A1(W3467), .A2(W2229), .ZN(O18782));
  NANDX1 G21213 (.A1(W37248), .A2(I416), .ZN(O18781));
  NANDX1 G21214 (.A1(W47448), .A2(W29765), .ZN(O18780));
  NANDX1 G21215 (.A1(W4894), .A2(W32185), .ZN(O18778));
  NANDX1 G21216 (.A1(W1161), .A2(W44974), .ZN(O18777));
  NANDX1 G21217 (.A1(W9471), .A2(W13813), .ZN(O18776));
  NANDX1 G21218 (.A1(W36399), .A2(W47758), .ZN(O18775));
  NANDX1 G21219 (.A1(W6462), .A2(W14647), .ZN(O18853));
  NANDX1 G21220 (.A1(W5603), .A2(W45967), .ZN(O18892));
  NANDX1 G21221 (.A1(W7934), .A2(W40056), .ZN(O18890));
  NANDX1 G21222 (.A1(W40885), .A2(W37151), .ZN(O18887));
  NANDX1 G21223 (.A1(W37517), .A2(W46135), .ZN(O18885));
  NANDX1 G21224 (.A1(W3942), .A2(W22688), .ZN(O18881));
  NANDX1 G21225 (.A1(W39734), .A2(W40314), .ZN(O18878));
  NANDX1 G21226 (.A1(W15522), .A2(W1869), .ZN(O18873));
  NANDX1 G21227 (.A1(W29761), .A2(W643), .ZN(O18872));
  NANDX1 G21228 (.A1(W29201), .A2(W37650), .ZN(O18866));
  NANDX1 G21229 (.A1(W5925), .A2(W27470), .ZN(O18861));
  NANDX1 G21230 (.A1(W15193), .A2(W48818), .ZN(O18858));
  NANDX1 G21231 (.A1(W25654), .A2(W20023), .ZN(O18855));
  NANDX1 G21232 (.A1(W34219), .A2(W40625), .ZN(O18774));
  NANDX1 G21233 (.A1(W7679), .A2(W4156), .ZN(W50072));
  NANDX1 G21234 (.A1(W50059), .A2(I715), .ZN(O18850));
  NANDX1 G21235 (.A1(W43885), .A2(W41565), .ZN(O18848));
  NANDX1 G21236 (.A1(W16879), .A2(W49178), .ZN(O18846));
  NANDX1 G21237 (.A1(W49624), .A2(W47787), .ZN(O18845));
  NANDX1 G21238 (.A1(W30963), .A2(W27543), .ZN(O18842));
  NANDX1 G21239 (.A1(W96), .A2(W37625), .ZN(O18840));
  NANDX1 G21240 (.A1(W16435), .A2(W32407), .ZN(W50059));
  NANDX1 G21241 (.A1(W19742), .A2(W25837), .ZN(O18838));
  NANDX1 G21242 (.A1(W41053), .A2(W43926), .ZN(O18836));
  NANDX1 G21243 (.A1(W34956), .A2(W18976), .ZN(O18833));
  NANDX1 G21244 (.A1(W27034), .A2(W13595), .ZN(O18664));
  NANDX1 G21245 (.A1(W34977), .A2(W42049), .ZN(O18701));
  NANDX1 G21246 (.A1(W32945), .A2(W41288), .ZN(O18697));
  NANDX1 G21247 (.A1(W20999), .A2(W41258), .ZN(O18693));
  NANDX1 G21248 (.A1(W43414), .A2(W27884), .ZN(O18692));
  NANDX1 G21249 (.A1(W42030), .A2(W47274), .ZN(O18686));
  NANDX1 G21250 (.A1(W41955), .A2(W33394), .ZN(O18683));
  NANDX1 G21251 (.A1(W7875), .A2(W28990), .ZN(O18681));
  NANDX1 G21252 (.A1(W74), .A2(W36243), .ZN(W49893));
  NANDX1 G21253 (.A1(W21854), .A2(W22004), .ZN(O18677));
  NANDX1 G21254 (.A1(W18638), .A2(W49190), .ZN(O18673));
  NANDX1 G21255 (.A1(W12345), .A2(W13883), .ZN(O18672));
  NANDX1 G21256 (.A1(W7277), .A2(W34764), .ZN(O18666));
  NANDX1 G21257 (.A1(W8264), .A2(W3618), .ZN(O18704));
  NANDX1 G21258 (.A1(W17137), .A2(W5046), .ZN(O18658));
  NANDX1 G21259 (.A1(W15023), .A2(W29399), .ZN(O18649));
  NANDX1 G21260 (.A1(W39625), .A2(W15650), .ZN(O18647));
  NANDX1 G21261 (.A1(W42233), .A2(W22907), .ZN(O18644));
  NANDX1 G21262 (.A1(W14575), .A2(W17614), .ZN(O18640));
  NANDX1 G21263 (.A1(W29032), .A2(W24855), .ZN(O18637));
  NANDX1 G21264 (.A1(W2789), .A2(W38259), .ZN(O18636));
  NANDX1 G21265 (.A1(W48614), .A2(W36582), .ZN(O18634));
  NANDX1 G21266 (.A1(W36661), .A2(W47675), .ZN(O18630));
  NANDX1 G21267 (.A1(W40167), .A2(I266), .ZN(O18628));
  NANDX1 G21268 (.A1(W5667), .A2(W17711), .ZN(O18626));
  NANDX1 G21269 (.A1(W41997), .A2(W32887), .ZN(O18751));
  NANDX1 G21270 (.A1(W12400), .A2(W16901), .ZN(O18772));
  NANDX1 G21271 (.A1(W43669), .A2(W9168), .ZN(O18769));
  NANDX1 G21272 (.A1(W38321), .A2(W2916), .ZN(O18768));
  NANDX1 G21273 (.A1(W35850), .A2(W10810), .ZN(O18766));
  NANDX1 G21274 (.A1(W49570), .A2(W20597), .ZN(O18765));
  NANDX1 G21275 (.A1(W27821), .A2(W28182), .ZN(O18764));
  NANDX1 G21276 (.A1(W28203), .A2(W48563), .ZN(O18760));
  NANDX1 G21277 (.A1(W44904), .A2(W41058), .ZN(O18757));
  NANDX1 G21278 (.A1(W36758), .A2(W3313), .ZN(O18756));
  NANDX1 G21279 (.A1(I437), .A2(W10725), .ZN(O18755));
  NANDX1 G21280 (.A1(W22410), .A2(W46335), .ZN(O18752));
  NANDX1 G21281 (.A1(W10706), .A2(W32504), .ZN(W50116));
  NANDX1 G21282 (.A1(W9602), .A2(W9805), .ZN(O18748));
  NANDX1 G21283 (.A1(W42847), .A2(W6086), .ZN(O18747));
  NANDX1 G21284 (.A1(W30423), .A2(W31297), .ZN(O18743));
  NANDX1 G21285 (.A1(W35768), .A2(W38549), .ZN(O18741));
  NANDX1 G21286 (.A1(W15496), .A2(W2514), .ZN(O18740));
  NANDX1 G21287 (.A1(W6639), .A2(W9951), .ZN(O18734));
  NANDX1 G21288 (.A1(W36249), .A2(W38663), .ZN(O18729));
  NANDX1 G21289 (.A1(W45349), .A2(W46329), .ZN(O18717));
  NANDX1 G21290 (.A1(W22422), .A2(W10095), .ZN(O18714));
  NANDX1 G21291 (.A1(W4782), .A2(W40669), .ZN(O18707));
  NANDX1 G21292 (.A1(W37859), .A2(W26707), .ZN(O18705));
  NANDX1 G21293 (.A1(I146), .A2(W11242), .ZN(O19052));
  NANDX1 G21294 (.A1(W1366), .A2(W30413), .ZN(O19096));
  NANDX1 G21295 (.A1(W15055), .A2(W49668), .ZN(O19095));
  NANDX1 G21296 (.A1(W14128), .A2(W9776), .ZN(O19091));
  NANDX1 G21297 (.A1(W18149), .A2(W19449), .ZN(O19090));
  NANDX1 G21298 (.A1(W29852), .A2(W872), .ZN(O19079));
  NANDX1 G21299 (.A1(W35426), .A2(W16487), .ZN(O19078));
  NANDX1 G21300 (.A1(W46969), .A2(I649), .ZN(O19076));
  NANDX1 G21301 (.A1(W21728), .A2(W9104), .ZN(O19068));
  NANDX1 G21302 (.A1(W4724), .A2(W14946), .ZN(O19067));
  NANDX1 G21303 (.A1(W31085), .A2(W14442), .ZN(O19065));
  NANDX1 G21304 (.A1(W29247), .A2(W40478), .ZN(O19062));
  NANDX1 G21305 (.A1(W20016), .A2(W49276), .ZN(O19055));
  NANDX1 G21306 (.A1(W21960), .A2(W29833), .ZN(O19100));
  NANDX1 G21307 (.A1(W23098), .A2(W30980), .ZN(O19050));
  NANDX1 G21308 (.A1(W32527), .A2(W34354), .ZN(O19041));
  NANDX1 G21309 (.A1(W32288), .A2(W31984), .ZN(O19036));
  NANDX1 G21310 (.A1(W4931), .A2(W40952), .ZN(O19032));
  NANDX1 G21311 (.A1(W47560), .A2(W39120), .ZN(O19030));
  NANDX1 G21312 (.A1(W47010), .A2(W31261), .ZN(O19021));
  NANDX1 G21313 (.A1(W42299), .A2(W34392), .ZN(O19015));
  NANDX1 G21314 (.A1(W34583), .A2(I1839), .ZN(W50242));
  NANDX1 G21315 (.A1(W46834), .A2(W41410), .ZN(O19008));
  NANDX1 G21316 (.A1(W36805), .A2(W34186), .ZN(O19004));
  NANDX1 G21317 (.A1(W47768), .A2(W26905), .ZN(O19003));
  NANDX1 G21318 (.A1(W14165), .A2(W2468), .ZN(O19130));
  NANDX1 G21319 (.A1(W36805), .A2(W24818), .ZN(O19160));
  NANDX1 G21320 (.A1(W30475), .A2(W38623), .ZN(O19159));
  NANDX1 G21321 (.A1(W2888), .A2(W8112), .ZN(O19153));
  NANDX1 G21322 (.A1(W29257), .A2(W38632), .ZN(O19148));
  NANDX1 G21323 (.A1(W28638), .A2(W4082), .ZN(O19147));
  NANDX1 G21324 (.A1(W27161), .A2(W48717), .ZN(O19146));
  NANDX1 G21325 (.A1(W43555), .A2(W46555), .ZN(O19145));
  NANDX1 G21326 (.A1(W18798), .A2(W49987), .ZN(O19144));
  NANDX1 G21327 (.A1(W1033), .A2(W21664), .ZN(O19137));
  NANDX1 G21328 (.A1(W39564), .A2(W34410), .ZN(O19134));
  NANDX1 G21329 (.A1(W14982), .A2(W32685), .ZN(O19131));
  NANDX1 G21330 (.A1(W18856), .A2(W23349), .ZN(O18998));
  NANDX1 G21331 (.A1(W10715), .A2(W49894), .ZN(O19129));
  NANDX1 G21332 (.A1(W49220), .A2(W28369), .ZN(O19125));
  NANDX1 G21333 (.A1(W40687), .A2(W35705), .ZN(O19121));
  NANDX1 G21334 (.A1(W5748), .A2(W11347), .ZN(O19119));
  NANDX1 G21335 (.A1(W22433), .A2(W3280), .ZN(O19117));
  NANDX1 G21336 (.A1(W10691), .A2(W42144), .ZN(O19113));
  NANDX1 G21337 (.A1(W35264), .A2(W36255), .ZN(O19111));
  NANDX1 G21338 (.A1(W39021), .A2(W6182), .ZN(O19110));
  NANDX1 G21339 (.A1(I900), .A2(W30041), .ZN(O19107));
  NANDX1 G21340 (.A1(W38054), .A2(W47631), .ZN(O19103));
  NANDX1 G21341 (.A1(W63), .A2(W19722), .ZN(O19102));
  NANDX1 G21342 (.A1(W17571), .A2(W37761), .ZN(O18928));
  NANDX1 G21343 (.A1(W49678), .A2(W44714), .ZN(O18949));
  NANDX1 G21344 (.A1(I245), .A2(W1705), .ZN(O18948));
  NANDX1 G21345 (.A1(W36824), .A2(W16264), .ZN(O18947));
  NANDX1 G21346 (.A1(W39766), .A2(W29924), .ZN(O18946));
  NANDX1 G21347 (.A1(W8260), .A2(W34183), .ZN(O18941));
  NANDX1 G21348 (.A1(W35809), .A2(W3806), .ZN(O18940));
  NANDX1 G21349 (.A1(W2018), .A2(W33077), .ZN(O18939));
  NANDX1 G21350 (.A1(W29205), .A2(W40192), .ZN(O18937));
  NANDX1 G21351 (.A1(W21375), .A2(W36983), .ZN(O18935));
  NANDX1 G21352 (.A1(W5345), .A2(W46951), .ZN(O18934));
  NANDX1 G21353 (.A1(W1118), .A2(W22948), .ZN(O18932));
  NANDX1 G21354 (.A1(W23542), .A2(I614), .ZN(O18929));
  NANDX1 G21355 (.A1(W32320), .A2(W2347), .ZN(O18950));
  NANDX1 G21356 (.A1(W19888), .A2(W20143), .ZN(O18927));
  NANDX1 G21357 (.A1(W11294), .A2(W21708), .ZN(O18924));
  NANDX1 G21358 (.A1(W50121), .A2(W30433), .ZN(O18922));
  NANDX1 G21359 (.A1(W34589), .A2(W14182), .ZN(O18920));
  NANDX1 G21360 (.A1(W3047), .A2(W29391), .ZN(O18919));
  NANDX1 G21361 (.A1(W26470), .A2(W1337), .ZN(O18918));
  NANDX1 G21362 (.A1(W28063), .A2(W21752), .ZN(O18914));
  NANDX1 G21363 (.A1(W9403), .A2(W32582), .ZN(O18913));
  NANDX1 G21364 (.A1(W22443), .A2(W20313), .ZN(O18910));
  NANDX1 G21365 (.A1(W7312), .A2(W36157), .ZN(O18909));
  NANDX1 G21366 (.A1(W11603), .A2(W49209), .ZN(O18900));
  NANDX1 G21367 (.A1(W32662), .A2(W8838), .ZN(O18973));
  NANDX1 G21368 (.A1(W32895), .A2(W43637), .ZN(W50225));
  NANDX1 G21369 (.A1(W12586), .A2(W27703), .ZN(O18996));
  NANDX1 G21370 (.A1(W28260), .A2(W3542), .ZN(O18995));
  NANDX1 G21371 (.A1(W4696), .A2(W41612), .ZN(O18994));
  NANDX1 G21372 (.A1(W13337), .A2(W18013), .ZN(O18993));
  NANDX1 G21373 (.A1(W14930), .A2(W15062), .ZN(O18990));
  NANDX1 G21374 (.A1(W23338), .A2(W3015), .ZN(O18989));
  NANDX1 G21375 (.A1(W43153), .A2(W6959), .ZN(O18986));
  NANDX1 G21376 (.A1(W45269), .A2(W7966), .ZN(O18983));
  NANDX1 G21377 (.A1(W29932), .A2(W5841), .ZN(O18981));
  NANDX1 G21378 (.A1(W9225), .A2(W40679), .ZN(O18974));
  NANDX1 G21379 (.A1(W35270), .A2(W17189), .ZN(O17489));
  NANDX1 G21380 (.A1(W35101), .A2(W26168), .ZN(O18972));
  NANDX1 G21381 (.A1(W30455), .A2(W26315), .ZN(W50198));
  NANDX1 G21382 (.A1(W36171), .A2(W36849), .ZN(O18970));
  NANDX1 G21383 (.A1(W34867), .A2(W28655), .ZN(O18967));
  NANDX1 G21384 (.A1(W6522), .A2(W26537), .ZN(O18964));
  NANDX1 G21385 (.A1(W20383), .A2(W23524), .ZN(O18962));
  NANDX1 G21386 (.A1(W44665), .A2(W23455), .ZN(O18961));
  NANDX1 G21387 (.A1(W14391), .A2(W15533), .ZN(O18959));
  NANDX1 G21388 (.A1(W6539), .A2(W303), .ZN(O18957));
  NANDX1 G21389 (.A1(W17030), .A2(W36535), .ZN(O18954));
  NANDX1 G21390 (.A1(W45585), .A2(W34257), .ZN(O18951));
  NANDX1 G21391 (.A1(W4083), .A2(W22266), .ZN(O15959));
  NANDX1 G21392 (.A1(W5831), .A2(W16642), .ZN(O15995));
  NANDX1 G21393 (.A1(W4422), .A2(W5783), .ZN(W46966));
  NANDX1 G21394 (.A1(W46277), .A2(W41942), .ZN(O15987));
  NANDX1 G21395 (.A1(W24725), .A2(W14856), .ZN(O15983));
  NANDX1 G21396 (.A1(W7400), .A2(W45179), .ZN(O15981));
  NANDX1 G21397 (.A1(W38678), .A2(W37577), .ZN(O15980));
  NANDX1 G21398 (.A1(W45517), .A2(W23026), .ZN(O15975));
  NANDX1 G21399 (.A1(W575), .A2(W2393), .ZN(O15972));
  NANDX1 G21400 (.A1(W23932), .A2(W5844), .ZN(O15969));
  NANDX1 G21401 (.A1(W40559), .A2(W16091), .ZN(O15968));
  NANDX1 G21402 (.A1(W24374), .A2(W18630), .ZN(O15965));
  NANDX1 G21403 (.A1(W2280), .A2(W38051), .ZN(O15960));
  NANDX1 G21404 (.A1(W22741), .A2(W28092), .ZN(O15996));
  NANDX1 G21405 (.A1(W33910), .A2(W37483), .ZN(O15958));
  NANDX1 G21406 (.A1(W35804), .A2(W42629), .ZN(O15957));
  NANDX1 G21407 (.A1(W15542), .A2(W30691), .ZN(O15956));
  NANDX1 G21408 (.A1(W14867), .A2(W18379), .ZN(O15954));
  NANDX1 G21409 (.A1(W27019), .A2(W18356), .ZN(O15953));
  NANDX1 G21410 (.A1(W10727), .A2(W10629), .ZN(O15952));
  NANDX1 G21411 (.A1(W5067), .A2(W45328), .ZN(O15951));
  NANDX1 G21412 (.A1(W16626), .A2(W17881), .ZN(O15950));
  NANDX1 G21413 (.A1(W22089), .A2(W42361), .ZN(O15949));
  NANDX1 G21414 (.A1(W7652), .A2(W42439), .ZN(O15948));
  NANDX1 G21415 (.A1(W43542), .A2(W1039), .ZN(O15943));
  NANDX1 G21416 (.A1(W45907), .A2(W31891), .ZN(O16020));
  NANDX1 G21417 (.A1(W7443), .A2(W3202), .ZN(O16046));
  NANDX1 G21418 (.A1(W23760), .A2(I433), .ZN(O16043));
  NANDX1 G21419 (.A1(W34878), .A2(W16528), .ZN(O16041));
  NANDX1 G21420 (.A1(W32283), .A2(W14467), .ZN(O16039));
  NANDX1 G21421 (.A1(W18550), .A2(W10922), .ZN(O16036));
  NANDX1 G21422 (.A1(I914), .A2(W17503), .ZN(O16033));
  NANDX1 G21423 (.A1(W8539), .A2(W19776), .ZN(O16031));
  NANDX1 G21424 (.A1(W41839), .A2(W23201), .ZN(O16026));
  NANDX1 G21425 (.A1(W5449), .A2(W19417), .ZN(O16024));
  NANDX1 G21426 (.A1(W22203), .A2(W30096), .ZN(W47004));
  NANDX1 G21427 (.A1(W11341), .A2(W6389), .ZN(O16022));
  NANDX1 G21428 (.A1(W24059), .A2(W13371), .ZN(O16021));
  NANDX1 G21429 (.A1(W15417), .A2(W34598), .ZN(O15941));
  NANDX1 G21430 (.A1(W5024), .A2(W39055), .ZN(O16012));
  NANDX1 G21431 (.A1(W17320), .A2(W17198), .ZN(O16009));
  NANDX1 G21432 (.A1(W23293), .A2(W15143), .ZN(W46987));
  NANDX1 G21433 (.A1(W29829), .A2(W38271), .ZN(O16008));
  NANDX1 G21434 (.A1(W36504), .A2(W32907), .ZN(W46985));
  NANDX1 G21435 (.A1(W34838), .A2(W16440), .ZN(O16005));
  NANDX1 G21436 (.A1(W38377), .A2(W43518), .ZN(O16004));
  NANDX1 G21437 (.A1(W31038), .A2(W423), .ZN(O16003));
  NANDX1 G21438 (.A1(W21905), .A2(W37309), .ZN(O16002));
  NANDX1 G21439 (.A1(W39092), .A2(W25913), .ZN(O16000));
  NANDX1 G21440 (.A1(W26303), .A2(W14397), .ZN(O15999));
  NANDX1 G21441 (.A1(W15181), .A2(W37971), .ZN(O15862));
  NANDX1 G21442 (.A1(W40988), .A2(W5059), .ZN(O15888));
  NANDX1 G21443 (.A1(W32472), .A2(W13416), .ZN(O15886));
  NANDX1 G21444 (.A1(W23873), .A2(W22603), .ZN(O15883));
  NANDX1 G21445 (.A1(W11936), .A2(W23375), .ZN(O15882));
  NANDX1 G21446 (.A1(W5983), .A2(W2661), .ZN(O15878));
  NANDX1 G21447 (.A1(W37426), .A2(W44665), .ZN(O15876));
  NANDX1 G21448 (.A1(W9484), .A2(W21543), .ZN(O15875));
  NANDX1 G21449 (.A1(W43301), .A2(W22422), .ZN(W46826));
  NANDX1 G21450 (.A1(I1135), .A2(W44603), .ZN(O15870));
  NANDX1 G21451 (.A1(W1199), .A2(W17041), .ZN(O15864));
  NANDX1 G21452 (.A1(W19465), .A2(W38110), .ZN(W46812));
  NANDX1 G21453 (.A1(W20594), .A2(W15801), .ZN(W46811));
  NANDX1 G21454 (.A1(W35704), .A2(W43136), .ZN(O15889));
  NANDX1 G21455 (.A1(W21859), .A2(W1023), .ZN(O15858));
  NANDX1 G21456 (.A1(W20905), .A2(W13789), .ZN(O15854));
  NANDX1 G21457 (.A1(W34834), .A2(W38762), .ZN(O15852));
  NANDX1 G21458 (.A1(W14137), .A2(W15733), .ZN(O15851));
  NANDX1 G21459 (.A1(W6021), .A2(W25472), .ZN(O15848));
  NANDX1 G21460 (.A1(W18957), .A2(W24544), .ZN(W46793));
  NANDX1 G21461 (.A1(W6019), .A2(W40039), .ZN(O15837));
  NANDX1 G21462 (.A1(W13353), .A2(W45111), .ZN(O15833));
  NANDX1 G21463 (.A1(W18804), .A2(W8945), .ZN(O15831));
  NANDX1 G21464 (.A1(W21461), .A2(W38225), .ZN(O15829));
  NANDX1 G21465 (.A1(W13453), .A2(W21102), .ZN(O15828));
  NANDX1 G21466 (.A1(W45594), .A2(W11634), .ZN(O15922));
  NANDX1 G21467 (.A1(W20155), .A2(I1629), .ZN(O15939));
  NANDX1 G21468 (.A1(W14547), .A2(W19380), .ZN(O15938));
  NANDX1 G21469 (.A1(W6662), .A2(W43825), .ZN(O15937));
  NANDX1 G21470 (.A1(W42139), .A2(W23520), .ZN(O15936));
  NANDX1 G21471 (.A1(W30391), .A2(W34189), .ZN(O15933));
  NANDX1 G21472 (.A1(W5926), .A2(W874), .ZN(O15932));
  NANDX1 G21473 (.A1(W5772), .A2(W17854), .ZN(O15928));
  NANDX1 G21474 (.A1(W40311), .A2(W20957), .ZN(O15925));
  NANDX1 G21475 (.A1(W7950), .A2(W40326), .ZN(W46888));
  NANDX1 G21476 (.A1(W40377), .A2(W33262), .ZN(O15923));
  NANDX1 G21477 (.A1(W18268), .A2(W107), .ZN(W46886));
  NANDX1 G21478 (.A1(W46059), .A2(W8101), .ZN(O16049));
  NANDX1 G21479 (.A1(W32734), .A2(W11254), .ZN(O15916));
  NANDX1 G21480 (.A1(W31117), .A2(I1202), .ZN(O15911));
  NANDX1 G21481 (.A1(W21028), .A2(W39142), .ZN(O15910));
  NANDX1 G21482 (.A1(W34402), .A2(W30243), .ZN(O15906));
  NANDX1 G21483 (.A1(W37249), .A2(W4715), .ZN(O15901));
  NANDX1 G21484 (.A1(W36952), .A2(W11231), .ZN(O15900));
  NANDX1 G21485 (.A1(W40451), .A2(W14138), .ZN(O15896));
  NANDX1 G21486 (.A1(W17740), .A2(W44702), .ZN(O15893));
  NANDX1 G21487 (.A1(W21249), .A2(W30830), .ZN(O15891));
  NANDX1 G21488 (.A1(W21460), .A2(W30659), .ZN(W46848));
  NANDX1 G21489 (.A1(W13375), .A2(W8115), .ZN(O15890));
  NANDX1 G21490 (.A1(W8945), .A2(W25935), .ZN(O16235));
  NANDX1 G21491 (.A1(W34524), .A2(W44548), .ZN(O16267));
  NANDX1 G21492 (.A1(W28975), .A2(W30707), .ZN(W47274));
  NANDX1 G21493 (.A1(W26894), .A2(W10859), .ZN(O16263));
  NANDX1 G21494 (.A1(W38308), .A2(W29175), .ZN(O16259));
  NANDX1 G21495 (.A1(W38171), .A2(W37323), .ZN(O16256));
  NANDX1 G21496 (.A1(W28441), .A2(W14208), .ZN(O16254));
  NANDX1 G21497 (.A1(W1949), .A2(W7652), .ZN(W47260));
  NANDX1 G21498 (.A1(W3685), .A2(W37392), .ZN(O16248));
  NANDX1 G21499 (.A1(W11870), .A2(W3538), .ZN(O16247));
  NANDX1 G21500 (.A1(W5755), .A2(W23909), .ZN(O16246));
  NANDX1 G21501 (.A1(W9974), .A2(W27993), .ZN(O16245));
  NANDX1 G21502 (.A1(W34129), .A2(W7407), .ZN(O16237));
  NANDX1 G21503 (.A1(W10510), .A2(W46587), .ZN(O16268));
  NANDX1 G21504 (.A1(W18551), .A2(W45232), .ZN(O16230));
  NANDX1 G21505 (.A1(W1720), .A2(W45412), .ZN(O16228));
  NANDX1 G21506 (.A1(W6536), .A2(W44940), .ZN(O16227));
  NANDX1 G21507 (.A1(W10812), .A2(W2356), .ZN(O16226));
  NANDX1 G21508 (.A1(W43411), .A2(W19298), .ZN(O16222));
  NANDX1 G21509 (.A1(W35185), .A2(W14773), .ZN(W47226));
  NANDX1 G21510 (.A1(W23614), .A2(W42515), .ZN(O16221));
  NANDX1 G21511 (.A1(W14619), .A2(W931), .ZN(O16215));
  NANDX1 G21512 (.A1(W2999), .A2(W3123), .ZN(O16203));
  NANDX1 G21513 (.A1(W41079), .A2(W14751), .ZN(O16202));
  NANDX1 G21514 (.A1(I1478), .A2(W22443), .ZN(O16200));
  NANDX1 G21515 (.A1(I21), .A2(W14093), .ZN(O16301));
  NANDX1 G21516 (.A1(W44064), .A2(W27235), .ZN(O16350));
  NANDX1 G21517 (.A1(W45895), .A2(W15015), .ZN(W47369));
  NANDX1 G21518 (.A1(W38311), .A2(W36457), .ZN(O16343));
  NANDX1 G21519 (.A1(W3026), .A2(W26016), .ZN(O16339));
  NANDX1 G21520 (.A1(W27508), .A2(W6144), .ZN(O16337));
  NANDX1 G21521 (.A1(W37432), .A2(W1632), .ZN(O16334));
  NANDX1 G21522 (.A1(I1255), .A2(W19131), .ZN(O16328));
  NANDX1 G21523 (.A1(W4052), .A2(W26548), .ZN(O16317));
  NANDX1 G21524 (.A1(W1310), .A2(W9721), .ZN(O16316));
  NANDX1 G21525 (.A1(W15947), .A2(W7409), .ZN(O16315));
  NANDX1 G21526 (.A1(W10351), .A2(W30341), .ZN(O16311));
  NANDX1 G21527 (.A1(W7603), .A2(W29255), .ZN(O16303));
  NANDX1 G21528 (.A1(W21196), .A2(W28044), .ZN(O16193));
  NANDX1 G21529 (.A1(W18036), .A2(W26855), .ZN(O16295));
  NANDX1 G21530 (.A1(W23414), .A2(W8049), .ZN(O16292));
  NANDX1 G21531 (.A1(W18223), .A2(W14107), .ZN(O16289));
  NANDX1 G21532 (.A1(W45500), .A2(W23050), .ZN(O16288));
  NANDX1 G21533 (.A1(W45165), .A2(W44120), .ZN(O16284));
  NANDX1 G21534 (.A1(W615), .A2(W5689), .ZN(O16281));
  NANDX1 G21535 (.A1(W22704), .A2(W46793), .ZN(O16280));
  NANDX1 G21536 (.A1(W13267), .A2(W5962), .ZN(O16278));
  NANDX1 G21537 (.A1(W12388), .A2(W13428), .ZN(O16276));
  NANDX1 G21538 (.A1(W4968), .A2(I267), .ZN(O16270));
  NANDX1 G21539 (.A1(W18414), .A2(W17265), .ZN(O16269));
  NANDX1 G21540 (.A1(W20143), .A2(W44903), .ZN(O16079));
  NANDX1 G21541 (.A1(W23101), .A2(W44162), .ZN(O16115));
  NANDX1 G21542 (.A1(W31277), .A2(W1320), .ZN(O16113));
  NANDX1 G21543 (.A1(W17557), .A2(W9815), .ZN(O16111));
  NANDX1 G21544 (.A1(W15268), .A2(W29224), .ZN(O16105));
  NANDX1 G21545 (.A1(W2378), .A2(W40024), .ZN(O16102));
  NANDX1 G21546 (.A1(W25709), .A2(W21000), .ZN(O16100));
  NANDX1 G21547 (.A1(W5603), .A2(W40263), .ZN(O16099));
  NANDX1 G21548 (.A1(W22163), .A2(W39251), .ZN(O16098));
  NANDX1 G21549 (.A1(W11190), .A2(W9589), .ZN(O16097));
  NANDX1 G21550 (.A1(W23768), .A2(W2056), .ZN(O16096));
  NANDX1 G21551 (.A1(W37844), .A2(W15812), .ZN(O16094));
  NANDX1 G21552 (.A1(W34743), .A2(W30852), .ZN(O16088));
  NANDX1 G21553 (.A1(W29057), .A2(W41819), .ZN(O16119));
  NANDX1 G21554 (.A1(W27357), .A2(W43404), .ZN(O16078));
  NANDX1 G21555 (.A1(W30574), .A2(W35195), .ZN(O16076));
  NANDX1 G21556 (.A1(W18179), .A2(W11027), .ZN(O16073));
  NANDX1 G21557 (.A1(I252), .A2(W43216), .ZN(O16071));
  NANDX1 G21558 (.A1(W40542), .A2(W9390), .ZN(O16068));
  NANDX1 G21559 (.A1(W14723), .A2(W5392), .ZN(O16064));
  NANDX1 G21560 (.A1(W39241), .A2(W36121), .ZN(O16059));
  NANDX1 G21561 (.A1(W44689), .A2(W42180), .ZN(W47041));
  NANDX1 G21562 (.A1(W31968), .A2(W39779), .ZN(O16054));
  NANDX1 G21563 (.A1(W45867), .A2(W13523), .ZN(O16053));
  NANDX1 G21564 (.A1(W7068), .A2(W14129), .ZN(O16050));
  NANDX1 G21565 (.A1(W46353), .A2(W25205), .ZN(O16164));
  NANDX1 G21566 (.A1(W33315), .A2(W13971), .ZN(O16191));
  NANDX1 G21567 (.A1(W10904), .A2(W10749), .ZN(O16187));
  NANDX1 G21568 (.A1(W33289), .A2(W34939), .ZN(O16186));
  NANDX1 G21569 (.A1(W25266), .A2(W6343), .ZN(O16182));
  NANDX1 G21570 (.A1(W2281), .A2(W5237), .ZN(W47180));
  NANDX1 G21571 (.A1(W38629), .A2(W19431), .ZN(O16179));
  NANDX1 G21572 (.A1(W3570), .A2(W6358), .ZN(O16176));
  NANDX1 G21573 (.A1(W15288), .A2(W30145), .ZN(O16175));
  NANDX1 G21574 (.A1(W18005), .A2(W9491), .ZN(O16173));
  NANDX1 G21575 (.A1(W38806), .A2(W29464), .ZN(O16170));
  NANDX1 G21576 (.A1(W17385), .A2(W37324), .ZN(O16166));
  NANDX1 G21577 (.A1(W41356), .A2(W3101), .ZN(O15826));
  NANDX1 G21578 (.A1(W303), .A2(W12107), .ZN(W47162));
  NANDX1 G21579 (.A1(W10178), .A2(W27801), .ZN(O16156));
  NANDX1 G21580 (.A1(W33048), .A2(I1593), .ZN(O16155));
  NANDX1 G21581 (.A1(W3198), .A2(W41265), .ZN(O16154));
  NANDX1 G21582 (.A1(W29998), .A2(W46369), .ZN(O16153));
  NANDX1 G21583 (.A1(W30877), .A2(W35773), .ZN(O16151));
  NANDX1 G21584 (.A1(W7127), .A2(W12005), .ZN(O16137));
  NANDX1 G21585 (.A1(W44192), .A2(W33527), .ZN(O16135));
  NANDX1 G21586 (.A1(W32026), .A2(W11156), .ZN(O16133));
  NANDX1 G21587 (.A1(W6539), .A2(W21048), .ZN(O16130));
  NANDX1 G21588 (.A1(W85), .A2(W5329), .ZN(O16128));
  NANDX1 G21589 (.A1(W34648), .A2(W10369), .ZN(O15525));
  NANDX1 G21590 (.A1(W18465), .A2(W16856), .ZN(O15549));
  NANDX1 G21591 (.A1(W4050), .A2(W39000), .ZN(O15546));
  NANDX1 G21592 (.A1(W32774), .A2(W8816), .ZN(O15545));
  NANDX1 G21593 (.A1(W31477), .A2(W36295), .ZN(O15541));
  NANDX1 G21594 (.A1(W37861), .A2(W27812), .ZN(O15539));
  NANDX1 G21595 (.A1(W17831), .A2(W5970), .ZN(O15536));
  NANDX1 G21596 (.A1(W12970), .A2(W10139), .ZN(W46425));
  NANDX1 G21597 (.A1(W27493), .A2(W39341), .ZN(O15535));
  NANDX1 G21598 (.A1(W18153), .A2(W19215), .ZN(O15534));
  NANDX1 G21599 (.A1(W17328), .A2(W1993), .ZN(O15533));
  NANDX1 G21600 (.A1(W42380), .A2(W19873), .ZN(O15529));
  NANDX1 G21601 (.A1(W10616), .A2(W39945), .ZN(O15526));
  NANDX1 G21602 (.A1(W4758), .A2(W17188), .ZN(O15550));
  NANDX1 G21603 (.A1(W39561), .A2(W3928), .ZN(O15523));
  NANDX1 G21604 (.A1(W45571), .A2(W32153), .ZN(O15520));
  NANDX1 G21605 (.A1(W3614), .A2(W26270), .ZN(O15519));
  NANDX1 G21606 (.A1(W31835), .A2(W27930), .ZN(O15517));
  NANDX1 G21607 (.A1(W42206), .A2(W32179), .ZN(O15515));
  NANDX1 G21608 (.A1(W27574), .A2(W14910), .ZN(O15514));
  NANDX1 G21609 (.A1(I1078), .A2(W44384), .ZN(O15513));
  NANDX1 G21610 (.A1(W29693), .A2(W4820), .ZN(O15509));
  NANDX1 G21611 (.A1(W18676), .A2(W37022), .ZN(O15508));
  NANDX1 G21612 (.A1(W9656), .A2(W42719), .ZN(O15507));
  NANDX1 G21613 (.A1(W18227), .A2(W43526), .ZN(O15505));
  NANDX1 G21614 (.A1(W14953), .A2(W23049), .ZN(O15592));
  NANDX1 G21615 (.A1(W6452), .A2(W32580), .ZN(W46517));
  NANDX1 G21616 (.A1(W466), .A2(W7723), .ZN(O15614));
  NANDX1 G21617 (.A1(W14057), .A2(W5221), .ZN(O15613));
  NANDX1 G21618 (.A1(W23078), .A2(W76), .ZN(O15612));
  NANDX1 G21619 (.A1(W18700), .A2(W9607), .ZN(O15607));
  NANDX1 G21620 (.A1(W1870), .A2(W44816), .ZN(O15606));
  NANDX1 G21621 (.A1(W39260), .A2(W17158), .ZN(O15605));
  NANDX1 G21622 (.A1(W42609), .A2(W10939), .ZN(O15604));
  NANDX1 G21623 (.A1(W42421), .A2(W37304), .ZN(O15601));
  NANDX1 G21624 (.A1(W30099), .A2(I346), .ZN(O15600));
  NANDX1 G21625 (.A1(W41754), .A2(W19100), .ZN(O15598));
  NANDX1 G21626 (.A1(W21260), .A2(W31556), .ZN(O15596));
  NANDX1 G21627 (.A1(W28431), .A2(W88), .ZN(O15504));
  NANDX1 G21628 (.A1(I1374), .A2(W23100), .ZN(W46475));
  NANDX1 G21629 (.A1(W21572), .A2(W17161), .ZN(O15578));
  NANDX1 G21630 (.A1(W40271), .A2(W30099), .ZN(O15576));
  NANDX1 G21631 (.A1(W38999), .A2(W15186), .ZN(O15574));
  NANDX1 G21632 (.A1(W10068), .A2(W42862), .ZN(O15573));
  NANDX1 G21633 (.A1(W36720), .A2(W18631), .ZN(O15564));
  NANDX1 G21634 (.A1(W35755), .A2(W21957), .ZN(O15559));
  NANDX1 G21635 (.A1(W28453), .A2(W32129), .ZN(O15558));
  NANDX1 G21636 (.A1(W9795), .A2(W32268), .ZN(O15556));
  NANDX1 G21637 (.A1(W22558), .A2(W5361), .ZN(O15554));
  NANDX1 G21638 (.A1(W19717), .A2(W3237), .ZN(O15552));
  NANDX1 G21639 (.A1(W12266), .A2(W30669), .ZN(O15403));
  NANDX1 G21640 (.A1(W17471), .A2(W11824), .ZN(O15439));
  NANDX1 G21641 (.A1(W22512), .A2(W24261), .ZN(O15436));
  NANDX1 G21642 (.A1(W20830), .A2(W6834), .ZN(O15433));
  NANDX1 G21643 (.A1(W26505), .A2(W20815), .ZN(O15431));
  NANDX1 G21644 (.A1(W44735), .A2(W23094), .ZN(W46299));
  NANDX1 G21645 (.A1(W44760), .A2(W42254), .ZN(O15423));
  NANDX1 G21646 (.A1(W17997), .A2(W38156), .ZN(O15421));
  NANDX1 G21647 (.A1(W19474), .A2(W38907), .ZN(O15419));
  NANDX1 G21648 (.A1(W11568), .A2(W24782), .ZN(O15417));
  NANDX1 G21649 (.A1(W4254), .A2(W30084), .ZN(O15409));
  NANDX1 G21650 (.A1(W6290), .A2(W5039), .ZN(O15407));
  NANDX1 G21651 (.A1(W17350), .A2(W17554), .ZN(O15405));
  NANDX1 G21652 (.A1(W10815), .A2(W6156), .ZN(O15450));
  NANDX1 G21653 (.A1(W18917), .A2(W25806), .ZN(O15401));
  NANDX1 G21654 (.A1(W24564), .A2(W2845), .ZN(O15400));
  NANDX1 G21655 (.A1(W37106), .A2(W35283), .ZN(O15399));
  NANDX1 G21656 (.A1(W23486), .A2(W36131), .ZN(O15398));
  NANDX1 G21657 (.A1(W43137), .A2(W23502), .ZN(O15394));
  NANDX1 G21658 (.A1(W22718), .A2(W30905), .ZN(O15387));
  NANDX1 G21659 (.A1(W26097), .A2(W12617), .ZN(O15383));
  NANDX1 G21660 (.A1(W13179), .A2(W13277), .ZN(O15381));
  NANDX1 G21661 (.A1(W11663), .A2(I1914), .ZN(O15380));
  NANDX1 G21662 (.A1(W2335), .A2(W38015), .ZN(W46241));
  NANDX1 G21663 (.A1(W44469), .A2(W15443), .ZN(W46239));
  NANDX1 G21664 (.A1(W46345), .A2(W19790), .ZN(O15482));
  NANDX1 G21665 (.A1(W1522), .A2(W21171), .ZN(O15501));
  NANDX1 G21666 (.A1(W42089), .A2(W16278), .ZN(O15500));
  NANDX1 G21667 (.A1(W8889), .A2(W20659), .ZN(O15496));
  NANDX1 G21668 (.A1(W18382), .A2(W8767), .ZN(O15495));
  NANDX1 G21669 (.A1(W15142), .A2(W7205), .ZN(W46378));
  NANDX1 G21670 (.A1(W6477), .A2(W36862), .ZN(O15491));
  NANDX1 G21671 (.A1(W35036), .A2(W10777), .ZN(O15490));
  NANDX1 G21672 (.A1(W19739), .A2(W24681), .ZN(W46372));
  NANDX1 G21673 (.A1(W7643), .A2(W18498), .ZN(W46369));
  NANDX1 G21674 (.A1(W40764), .A2(W39196), .ZN(O15487));
  NANDX1 G21675 (.A1(W3210), .A2(W15605), .ZN(O15484));
  NANDX1 G21676 (.A1(W27983), .A2(W41976), .ZN(O15616));
  NANDX1 G21677 (.A1(W12325), .A2(W11301), .ZN(O15479));
  NANDX1 G21678 (.A1(W45606), .A2(W7054), .ZN(O15477));
  NANDX1 G21679 (.A1(W21754), .A2(W29404), .ZN(O15473));
  NANDX1 G21680 (.A1(W6620), .A2(W37954), .ZN(O15472));
  NANDX1 G21681 (.A1(W10952), .A2(W15107), .ZN(O15469));
  NANDX1 G21682 (.A1(W40768), .A2(W1644), .ZN(O15468));
  NANDX1 G21683 (.A1(W37043), .A2(W13340), .ZN(O15461));
  NANDX1 G21684 (.A1(W33154), .A2(W21365), .ZN(W46335));
  NANDX1 G21685 (.A1(W16078), .A2(W9241), .ZN(O15457));
  NANDX1 G21686 (.A1(W15258), .A2(I1021), .ZN(O15453));
  NANDX1 G21687 (.A1(W25051), .A2(W33839), .ZN(W46325));
  NANDX1 G21688 (.A1(W141), .A2(W25094), .ZN(O15754));
  NANDX1 G21689 (.A1(W10551), .A2(W45470), .ZN(O15783));
  NANDX1 G21690 (.A1(W33291), .A2(W11000), .ZN(O15781));
  NANDX1 G21691 (.A1(W7108), .A2(W1653), .ZN(W46714));
  NANDX1 G21692 (.A1(W7811), .A2(W20856), .ZN(O15778));
  NANDX1 G21693 (.A1(W9118), .A2(W42359), .ZN(W46707));
  NANDX1 G21694 (.A1(W37844), .A2(W1030), .ZN(O15772));
  NANDX1 G21695 (.A1(I117), .A2(W20482), .ZN(O15771));
  NANDX1 G21696 (.A1(W17956), .A2(W43932), .ZN(O15770));
  NANDX1 G21697 (.A1(W16428), .A2(W954), .ZN(O15766));
  NANDX1 G21698 (.A1(W18430), .A2(W35312), .ZN(O15764));
  NANDX1 G21699 (.A1(W26773), .A2(W29385), .ZN(O15758));
  NANDX1 G21700 (.A1(W26079), .A2(W39107), .ZN(O15755));
  NANDX1 G21701 (.A1(W44018), .A2(W7146), .ZN(O15784));
  NANDX1 G21702 (.A1(W37967), .A2(W9376), .ZN(O15753));
  NANDX1 G21703 (.A1(W17798), .A2(W30607), .ZN(O15751));
  NANDX1 G21704 (.A1(W31267), .A2(W38869), .ZN(O15748));
  NANDX1 G21705 (.A1(W40292), .A2(W42221), .ZN(O15745));
  NANDX1 G21706 (.A1(W38511), .A2(W17285), .ZN(O15739));
  NANDX1 G21707 (.A1(W24670), .A2(W6220), .ZN(O15735));
  NANDX1 G21708 (.A1(W18406), .A2(W17778), .ZN(O15731));
  NANDX1 G21709 (.A1(W9436), .A2(W26116), .ZN(O15728));
  NANDX1 G21710 (.A1(I1925), .A2(W25619), .ZN(O15727));
  NANDX1 G21711 (.A1(W4492), .A2(W10989), .ZN(O15726));
  NANDX1 G21712 (.A1(W30639), .A2(W40262), .ZN(O15723));
  NANDX1 G21713 (.A1(W18908), .A2(W43566), .ZN(O15797));
  NANDX1 G21714 (.A1(W39629), .A2(W40054), .ZN(O15825));
  NANDX1 G21715 (.A1(W33060), .A2(W5657), .ZN(O15823));
  NANDX1 G21716 (.A1(W15014), .A2(W24308), .ZN(W46764));
  NANDX1 G21717 (.A1(W20099), .A2(I1818), .ZN(O15819));
  NANDX1 G21718 (.A1(W41288), .A2(W28270), .ZN(W46753));
  NANDX1 G21719 (.A1(W20653), .A2(W46325), .ZN(O15812));
  NANDX1 G21720 (.A1(W32374), .A2(W35132), .ZN(O15810));
  NANDX1 G21721 (.A1(W46734), .A2(I1530), .ZN(O15809));
  NANDX1 G21722 (.A1(W45302), .A2(W12501), .ZN(W46748));
  NANDX1 G21723 (.A1(W10757), .A2(W2784), .ZN(O15806));
  NANDX1 G21724 (.A1(W45365), .A2(W45924), .ZN(O15801));
  NANDX1 G21725 (.A1(W11803), .A2(W25239), .ZN(O15722));
  NANDX1 G21726 (.A1(W41279), .A2(W44694), .ZN(W46734));
  NANDX1 G21727 (.A1(W24055), .A2(W3014), .ZN(W46732));
  NANDX1 G21728 (.A1(W41981), .A2(W4647), .ZN(O15795));
  NANDX1 G21729 (.A1(W11833), .A2(W46533), .ZN(W46729));
  NANDX1 G21730 (.A1(W10017), .A2(W1264), .ZN(O15794));
  NANDX1 G21731 (.A1(W22014), .A2(W2780), .ZN(O15793));
  NANDX1 G21732 (.A1(W2948), .A2(W5239), .ZN(O15792));
  NANDX1 G21733 (.A1(W45456), .A2(W18512), .ZN(O15791));
  NANDX1 G21734 (.A1(W29620), .A2(W25457), .ZN(O15790));
  NANDX1 G21735 (.A1(W40932), .A2(W26522), .ZN(O15787));
  NANDX1 G21736 (.A1(W6027), .A2(W40626), .ZN(O15786));
  NANDX1 G21737 (.A1(I877), .A2(W28752), .ZN(O15641));
  NANDX1 G21738 (.A1(W31394), .A2(W5400), .ZN(O15662));
  NANDX1 G21739 (.A1(W12889), .A2(I1232), .ZN(O15659));
  NANDX1 G21740 (.A1(W10436), .A2(W11625), .ZN(O15658));
  NANDX1 G21741 (.A1(W36605), .A2(W7211), .ZN(O15657));
  NANDX1 G21742 (.A1(W17462), .A2(W2328), .ZN(O15653));
  NANDX1 G21743 (.A1(W30188), .A2(W1302), .ZN(O15652));
  NANDX1 G21744 (.A1(W42745), .A2(W32768), .ZN(W46561));
  NANDX1 G21745 (.A1(W45463), .A2(W25568), .ZN(O15650));
  NANDX1 G21746 (.A1(W34428), .A2(W23375), .ZN(O15649));
  NANDX1 G21747 (.A1(W7086), .A2(W40190), .ZN(W46555));
  NANDX1 G21748 (.A1(W43100), .A2(W7384), .ZN(O15643));
  NANDX1 G21749 (.A1(W4828), .A2(W7010), .ZN(O15642));
  NANDX1 G21750 (.A1(W38031), .A2(W17892), .ZN(O15664));
  NANDX1 G21751 (.A1(W22366), .A2(W38809), .ZN(O15639));
  NANDX1 G21752 (.A1(W14352), .A2(W28426), .ZN(W46544));
  NANDX1 G21753 (.A1(W800), .A2(W38872), .ZN(O15638));
  NANDX1 G21754 (.A1(W5604), .A2(W36721), .ZN(O15633));
  NANDX1 G21755 (.A1(W40007), .A2(W38415), .ZN(O15630));
  NANDX1 G21756 (.A1(W43135), .A2(W26906), .ZN(O15629));
  NANDX1 G21757 (.A1(W1046), .A2(W33491), .ZN(W46531));
  NANDX1 G21758 (.A1(W41791), .A2(W22036), .ZN(O15627));
  NANDX1 G21759 (.A1(W28806), .A2(W23829), .ZN(O15625));
  NANDX1 G21760 (.A1(W33265), .A2(W21774), .ZN(O15620));
  NANDX1 G21761 (.A1(W35525), .A2(W28007), .ZN(O15618));
  NANDX1 G21762 (.A1(W39079), .A2(W10531), .ZN(W46621));
  NANDX1 G21763 (.A1(W13145), .A2(W1618), .ZN(W46641));
  NANDX1 G21764 (.A1(W26577), .A2(W7579), .ZN(O15717));
  NANDX1 G21765 (.A1(W4077), .A2(W17030), .ZN(W46638));
  NANDX1 G21766 (.A1(W8355), .A2(W18474), .ZN(O15714));
  NANDX1 G21767 (.A1(W10139), .A2(W3385), .ZN(W46635));
  NANDX1 G21768 (.A1(W22953), .A2(W19181), .ZN(O15712));
  NANDX1 G21769 (.A1(W2897), .A2(W32188), .ZN(O15710));
  NANDX1 G21770 (.A1(W26448), .A2(W7966), .ZN(O15705));
  NANDX1 G21771 (.A1(W5037), .A2(W36733), .ZN(W46624));
  NANDX1 G21772 (.A1(W34298), .A2(W40951), .ZN(O15703));
  NANDX1 G21773 (.A1(W5174), .A2(W12714), .ZN(O15702));
  NANDX1 G21774 (.A1(W27474), .A2(W46605), .ZN(O16351));
  NANDX1 G21775 (.A1(W27773), .A2(W32719), .ZN(O15692));
  NANDX1 G21776 (.A1(W690), .A2(W43276), .ZN(O15690));
  NANDX1 G21777 (.A1(W5126), .A2(W42296), .ZN(O15687));
  NANDX1 G21778 (.A1(I248), .A2(W42708), .ZN(O15685));
  NANDX1 G21779 (.A1(W4033), .A2(W18696), .ZN(O15679));
  NANDX1 G21780 (.A1(W10588), .A2(W3888), .ZN(O15676));
  NANDX1 G21781 (.A1(W29981), .A2(W43142), .ZN(W46589));
  NANDX1 G21782 (.A1(W5065), .A2(W43928), .ZN(O15674));
  NANDX1 G21783 (.A1(W39078), .A2(W41400), .ZN(O15672));
  NANDX1 G21784 (.A1(W34611), .A2(W29849), .ZN(O15669));
  NANDX1 G21785 (.A1(W23081), .A2(W9208), .ZN(O15667));
  NANDX1 G21786 (.A1(W1579), .A2(W10612), .ZN(O17076));
  NANDX1 G21787 (.A1(W41653), .A2(W36535), .ZN(O17114));
  NANDX1 G21788 (.A1(W43373), .A2(W21171), .ZN(O17111));
  NANDX1 G21789 (.A1(W13167), .A2(W38787), .ZN(O17107));
  NANDX1 G21790 (.A1(W19368), .A2(W28785), .ZN(O17103));
  NANDX1 G21791 (.A1(W22850), .A2(W16699), .ZN(O17102));
  NANDX1 G21792 (.A1(I1385), .A2(W2298), .ZN(O17099));
  NANDX1 G21793 (.A1(W7927), .A2(W19676), .ZN(O17094));
  NANDX1 G21794 (.A1(W15260), .A2(W13790), .ZN(O17093));
  NANDX1 G21795 (.A1(W5177), .A2(W5039), .ZN(O17089));
  NANDX1 G21796 (.A1(W31502), .A2(W6261), .ZN(W48183));
  NANDX1 G21797 (.A1(W8160), .A2(W22831), .ZN(O17086));
  NANDX1 G21798 (.A1(I332), .A2(W43051), .ZN(O17082));
  NANDX1 G21799 (.A1(W42648), .A2(W36499), .ZN(O17117));
  NANDX1 G21800 (.A1(W36557), .A2(W31596), .ZN(O17074));
  NANDX1 G21801 (.A1(W39788), .A2(W15602), .ZN(O17073));
  NANDX1 G21802 (.A1(W34217), .A2(W47066), .ZN(O17064));
  NANDX1 G21803 (.A1(W46561), .A2(W13973), .ZN(O17062));
  NANDX1 G21804 (.A1(W40396), .A2(W31177), .ZN(O17058));
  NANDX1 G21805 (.A1(W43223), .A2(W1516), .ZN(O17053));
  NANDX1 G21806 (.A1(W14537), .A2(W27555), .ZN(O17050));
  NANDX1 G21807 (.A1(W28758), .A2(W12063), .ZN(O17049));
  NANDX1 G21808 (.A1(W16083), .A2(W47369), .ZN(O17047));
  NANDX1 G21809 (.A1(I1826), .A2(W11388), .ZN(O17045));
  NANDX1 G21810 (.A1(W18538), .A2(W26111), .ZN(O17044));
  NANDX1 G21811 (.A1(W43423), .A2(W31741), .ZN(O17138));
  NANDX1 G21812 (.A1(W1364), .A2(W6618), .ZN(O17184));
  NANDX1 G21813 (.A1(W35059), .A2(W4070), .ZN(O17179));
  NANDX1 G21814 (.A1(W7755), .A2(W8446), .ZN(O17176));
  NANDX1 G21815 (.A1(W2303), .A2(W24965), .ZN(O17175));
  NANDX1 G21816 (.A1(W9887), .A2(I564), .ZN(O17174));
  NANDX1 G21817 (.A1(W45792), .A2(W44190), .ZN(O17165));
  NANDX1 G21818 (.A1(W35845), .A2(W7780), .ZN(O17164));
  NANDX1 G21819 (.A1(W7147), .A2(W25404), .ZN(O17163));
  NANDX1 G21820 (.A1(W29504), .A2(W30853), .ZN(O17162));
  NANDX1 G21821 (.A1(W15524), .A2(W27574), .ZN(O17154));
  NANDX1 G21822 (.A1(W28113), .A2(W8725), .ZN(O17143));
  NANDX1 G21823 (.A1(W30509), .A2(W15371), .ZN(O17141));
  NANDX1 G21824 (.A1(W15633), .A2(W15348), .ZN(O17040));
  NANDX1 G21825 (.A1(W33945), .A2(W43604), .ZN(W48234));
  NANDX1 G21826 (.A1(W30737), .A2(W19193), .ZN(O17132));
  NANDX1 G21827 (.A1(W14089), .A2(W25578), .ZN(W48226));
  NANDX1 G21828 (.A1(W10280), .A2(W19175), .ZN(O17129));
  NANDX1 G21829 (.A1(W31972), .A2(W22586), .ZN(O17128));
  NANDX1 G21830 (.A1(I791), .A2(W33698), .ZN(O17127));
  NANDX1 G21831 (.A1(W29961), .A2(W34591), .ZN(O17126));
  NANDX1 G21832 (.A1(W12132), .A2(W22134), .ZN(O17124));
  NANDX1 G21833 (.A1(W28171), .A2(W21216), .ZN(O17122));
  NANDX1 G21834 (.A1(W22469), .A2(W39714), .ZN(O17119));
  NANDX1 G21835 (.A1(W41021), .A2(W11689), .ZN(O17118));
  NANDX1 G21836 (.A1(I643), .A2(W40368), .ZN(W48022));
  NANDX1 G21837 (.A1(W46475), .A2(W32131), .ZN(O16973));
  NANDX1 G21838 (.A1(W36252), .A2(W18282), .ZN(O16966));
  NANDX1 G21839 (.A1(I1945), .A2(W8149), .ZN(O16965));
  NANDX1 G21840 (.A1(W40076), .A2(W2978), .ZN(O16958));
  NANDX1 G21841 (.A1(W31971), .A2(W20836), .ZN(O16957));
  NANDX1 G21842 (.A1(W29123), .A2(W4490), .ZN(O16956));
  NANDX1 G21843 (.A1(W9142), .A2(W19894), .ZN(O16951));
  NANDX1 G21844 (.A1(W24408), .A2(W4579), .ZN(O16949));
  NANDX1 G21845 (.A1(W8641), .A2(W14370), .ZN(O16948));
  NANDX1 G21846 (.A1(W11831), .A2(W3747), .ZN(O16946));
  NANDX1 G21847 (.A1(W11390), .A2(W39489), .ZN(O16944));
  NANDX1 G21848 (.A1(W38574), .A2(W16332), .ZN(O16942));
  NANDX1 G21849 (.A1(W47126), .A2(W1392), .ZN(O16977));
  NANDX1 G21850 (.A1(W5881), .A2(W15424), .ZN(O16940));
  NANDX1 G21851 (.A1(W14415), .A2(W404), .ZN(O16934));
  NANDX1 G21852 (.A1(W28342), .A2(W41880), .ZN(O16932));
  NANDX1 G21853 (.A1(W24583), .A2(W35837), .ZN(O16930));
  NANDX1 G21854 (.A1(W3336), .A2(W27038), .ZN(O16927));
  NANDX1 G21855 (.A1(W33524), .A2(W47145), .ZN(O16924));
  NANDX1 G21856 (.A1(W9970), .A2(W12812), .ZN(O16923));
  NANDX1 G21857 (.A1(W2381), .A2(W8056), .ZN(O16921));
  NANDX1 G21858 (.A1(W28008), .A2(W42946), .ZN(O16920));
  NANDX1 G21859 (.A1(W38591), .A2(W5794), .ZN(O16918));
  NANDX1 G21860 (.A1(W29608), .A2(W11674), .ZN(W47993));
  NANDX1 G21861 (.A1(W32554), .A2(W10098), .ZN(O17004));
  NANDX1 G21862 (.A1(W22800), .A2(W34713), .ZN(O17039));
  NANDX1 G21863 (.A1(W24924), .A2(W27657), .ZN(O17038));
  NANDX1 G21864 (.A1(W43236), .A2(W22233), .ZN(O17037));
  NANDX1 G21865 (.A1(W23961), .A2(W4870), .ZN(O17035));
  NANDX1 G21866 (.A1(W23056), .A2(W36125), .ZN(O17034));
  NANDX1 G21867 (.A1(W19866), .A2(W3426), .ZN(O17033));
  NANDX1 G21868 (.A1(W13401), .A2(W16520), .ZN(O17032));
  NANDX1 G21869 (.A1(W34178), .A2(W40670), .ZN(W48114));
  NANDX1 G21870 (.A1(W15797), .A2(W35571), .ZN(W48106));
  NANDX1 G21871 (.A1(W14017), .A2(W14091), .ZN(O17020));
  NANDX1 G21872 (.A1(W1922), .A2(W24928), .ZN(O17013));
  NANDX1 G21873 (.A1(W45255), .A2(W4570), .ZN(O17186));
  NANDX1 G21874 (.A1(I1324), .A2(W46714), .ZN(O17003));
  NANDX1 G21875 (.A1(W30030), .A2(W7194), .ZN(O17001));
  NANDX1 G21876 (.A1(W22960), .A2(W19591), .ZN(O17000));
  NANDX1 G21877 (.A1(W25031), .A2(W28059), .ZN(O16996));
  NANDX1 G21878 (.A1(W35050), .A2(W2642), .ZN(O16995));
  NANDX1 G21879 (.A1(I1248), .A2(W28280), .ZN(O16994));
  NANDX1 G21880 (.A1(W384), .A2(W6786), .ZN(W48073));
  NANDX1 G21881 (.A1(W37041), .A2(W8312), .ZN(O16989));
  NANDX1 G21882 (.A1(W37401), .A2(W24314), .ZN(O16985));
  NANDX1 G21883 (.A1(W7961), .A2(W6499), .ZN(O16982));
  NANDX1 G21884 (.A1(W34743), .A2(W26476), .ZN(O16980));
  NANDX1 G21885 (.A1(W12839), .A2(W37049), .ZN(O17371));
  NANDX1 G21886 (.A1(W43477), .A2(W44135), .ZN(O17397));
  NANDX1 G21887 (.A1(W3112), .A2(W22219), .ZN(O17395));
  NANDX1 G21888 (.A1(I212), .A2(W9067), .ZN(O17387));
  NANDX1 G21889 (.A1(W36615), .A2(W19027), .ZN(O17386));
  NANDX1 G21890 (.A1(W9421), .A2(W2548), .ZN(O17385));
  NANDX1 G21891 (.A1(W4653), .A2(W14758), .ZN(O17383));
  NANDX1 G21892 (.A1(W1503), .A2(W17723), .ZN(O17382));
  NANDX1 G21893 (.A1(W17291), .A2(W18952), .ZN(O17381));
  NANDX1 G21894 (.A1(W346), .A2(W29070), .ZN(O17379));
  NANDX1 G21895 (.A1(W2495), .A2(I353), .ZN(O17377));
  NANDX1 G21896 (.A1(W14291), .A2(W10939), .ZN(O17376));
  NANDX1 G21897 (.A1(W27732), .A2(W42092), .ZN(O17374));
  NANDX1 G21898 (.A1(W30591), .A2(W31133), .ZN(O17399));
  NANDX1 G21899 (.A1(W43176), .A2(W16798), .ZN(O17369));
  NANDX1 G21900 (.A1(W39992), .A2(W7265), .ZN(O17363));
  NANDX1 G21901 (.A1(W17487), .A2(W5529), .ZN(O17360));
  NANDX1 G21902 (.A1(W6936), .A2(W191), .ZN(O17356));
  NANDX1 G21903 (.A1(W28778), .A2(W22395), .ZN(O17354));
  NANDX1 G21904 (.A1(W25430), .A2(I22), .ZN(O17352));
  NANDX1 G21905 (.A1(W11830), .A2(W2443), .ZN(O17349));
  NANDX1 G21906 (.A1(W20006), .A2(W27376), .ZN(O17346));
  NANDX1 G21907 (.A1(W15406), .A2(W40976), .ZN(O17343));
  NANDX1 G21908 (.A1(W27799), .A2(W28765), .ZN(O17342));
  NANDX1 G21909 (.A1(W14956), .A2(W47216), .ZN(O17340));
  NANDX1 G21910 (.A1(W25584), .A2(W48389), .ZN(O17437));
  NANDX1 G21911 (.A1(W15198), .A2(W43402), .ZN(O17482));
  NANDX1 G21912 (.A1(W7463), .A2(W5585), .ZN(O17479));
  NANDX1 G21913 (.A1(W15265), .A2(W16083), .ZN(O17476));
  NANDX1 G21914 (.A1(W29156), .A2(W32443), .ZN(O17475));
  NANDX1 G21915 (.A1(I715), .A2(W9803), .ZN(O17470));
  NANDX1 G21916 (.A1(W45832), .A2(W35774), .ZN(O17469));
  NANDX1 G21917 (.A1(W20730), .A2(W32464), .ZN(O17465));
  NANDX1 G21918 (.A1(W37362), .A2(W35100), .ZN(O17453));
  NANDX1 G21919 (.A1(W38157), .A2(W22463), .ZN(O17451));
  NANDX1 G21920 (.A1(W6374), .A2(W19078), .ZN(O17449));
  NANDX1 G21921 (.A1(W6024), .A2(W5219), .ZN(W48577));
  NANDX1 G21922 (.A1(W9133), .A2(W46635), .ZN(O17439));
  NANDX1 G21923 (.A1(W11185), .A2(W1296), .ZN(O17336));
  NANDX1 G21924 (.A1(W46595), .A2(W7354), .ZN(O17436));
  NANDX1 G21925 (.A1(W3542), .A2(W45299), .ZN(O17434));
  NANDX1 G21926 (.A1(W36580), .A2(W36205), .ZN(O17432));
  NANDX1 G21927 (.A1(W1621), .A2(W14453), .ZN(O17424));
  NANDX1 G21928 (.A1(W5103), .A2(W3096), .ZN(W48540));
  NANDX1 G21929 (.A1(W46589), .A2(W43), .ZN(W48537));
  NANDX1 G21930 (.A1(W8329), .A2(W7491), .ZN(O17419));
  NANDX1 G21931 (.A1(I168), .A2(W35509), .ZN(O17412));
  NANDX1 G21932 (.A1(W7755), .A2(W7592), .ZN(O17407));
  NANDX1 G21933 (.A1(W22553), .A2(W45925), .ZN(O17405));
  NANDX1 G21934 (.A1(W14555), .A2(W29202), .ZN(O17403));
  NANDX1 G21935 (.A1(W45929), .A2(W29296), .ZN(O17231));
  NANDX1 G21936 (.A1(W41825), .A2(W20228), .ZN(O17267));
  NANDX1 G21937 (.A1(W21639), .A2(W22478), .ZN(O17264));
  NANDX1 G21938 (.A1(W11075), .A2(W14010), .ZN(O17262));
  NANDX1 G21939 (.A1(W39088), .A2(W26567), .ZN(O17261));
  NANDX1 G21940 (.A1(W40484), .A2(W3187), .ZN(O17258));
  NANDX1 G21941 (.A1(W1479), .A2(W27915), .ZN(O17257));
  NANDX1 G21942 (.A1(W15450), .A2(W21249), .ZN(O17253));
  NANDX1 G21943 (.A1(W25638), .A2(W34383), .ZN(O17250));
  NANDX1 G21944 (.A1(W38186), .A2(W14652), .ZN(O17245));
  NANDX1 G21945 (.A1(W12404), .A2(W22641), .ZN(O17241));
  NANDX1 G21946 (.A1(W28254), .A2(W35355), .ZN(O17239));
  NANDX1 G21947 (.A1(W14957), .A2(W35045), .ZN(O17232));
  NANDX1 G21948 (.A1(W37439), .A2(W41252), .ZN(O17268));
  NANDX1 G21949 (.A1(W13411), .A2(W11793), .ZN(O17229));
  NANDX1 G21950 (.A1(W47632), .A2(W21014), .ZN(O17227));
  NANDX1 G21951 (.A1(W31985), .A2(W45267), .ZN(O17222));
  NANDX1 G21952 (.A1(W29122), .A2(W23796), .ZN(W48322));
  NANDX1 G21953 (.A1(W41031), .A2(W22186), .ZN(O17217));
  NANDX1 G21954 (.A1(W15437), .A2(W47299), .ZN(O17214));
  NANDX1 G21955 (.A1(I5), .A2(W21923), .ZN(O17209));
  NANDX1 G21956 (.A1(I1917), .A2(W20025), .ZN(O17203));
  NANDX1 G21957 (.A1(W3811), .A2(W44646), .ZN(O17198));
  NANDX1 G21958 (.A1(W2643), .A2(W45726), .ZN(O17197));
  NANDX1 G21959 (.A1(W24240), .A2(W3674), .ZN(O17189));
  NANDX1 G21960 (.A1(W32725), .A2(W26595), .ZN(O17301));
  NANDX1 G21961 (.A1(W42862), .A2(W43957), .ZN(O17334));
  NANDX1 G21962 (.A1(W29225), .A2(W31663), .ZN(O17329));
  NANDX1 G21963 (.A1(W4848), .A2(W8360), .ZN(O17327));
  NANDX1 G21964 (.A1(W22765), .A2(W34822), .ZN(O17322));
  NANDX1 G21965 (.A1(W31906), .A2(W44903), .ZN(O17317));
  NANDX1 G21966 (.A1(W18206), .A2(W15402), .ZN(O17316));
  NANDX1 G21967 (.A1(W47763), .A2(W41248), .ZN(O17314));
  NANDX1 G21968 (.A1(W8430), .A2(W20525), .ZN(O17313));
  NANDX1 G21969 (.A1(W3006), .A2(W39264), .ZN(O17311));
  NANDX1 G21970 (.A1(W15588), .A2(W7826), .ZN(O17310));
  NANDX1 G21971 (.A1(W1270), .A2(W28023), .ZN(O17309));
  NANDX1 G21972 (.A1(W41647), .A2(I693), .ZN(O16913));
  NANDX1 G21973 (.A1(W18865), .A2(W27566), .ZN(O17298));
  NANDX1 G21974 (.A1(W10129), .A2(W32671), .ZN(O17296));
  NANDX1 G21975 (.A1(W7933), .A2(W22608), .ZN(O17288));
  NANDX1 G21976 (.A1(I458), .A2(W8667), .ZN(W48396));
  NANDX1 G21977 (.A1(W34729), .A2(I1092), .ZN(W48395));
  NANDX1 G21978 (.A1(W37465), .A2(W27008), .ZN(O17286));
  NANDX1 G21979 (.A1(W37615), .A2(W36679), .ZN(O17284));
  NANDX1 G21980 (.A1(W12187), .A2(W26001), .ZN(O17277));
  NANDX1 G21981 (.A1(W6604), .A2(W44687), .ZN(O17276));
  NANDX1 G21982 (.A1(W15795), .A2(W26721), .ZN(O17275));
  NANDX1 G21983 (.A1(W41791), .A2(W44619), .ZN(O17273));
  NANDX1 G21984 (.A1(W40396), .A2(W19474), .ZN(O16521));
  NANDX1 G21985 (.A1(W5529), .A2(W20543), .ZN(O16556));
  NANDX1 G21986 (.A1(W43417), .A2(W4494), .ZN(O16553));
  NANDX1 G21987 (.A1(W3293), .A2(W2051), .ZN(O16551));
  NANDX1 G21988 (.A1(W638), .A2(W24507), .ZN(O16547));
  NANDX1 G21989 (.A1(W3105), .A2(W25718), .ZN(O16542));
  NANDX1 G21990 (.A1(W30435), .A2(W10835), .ZN(O16541));
  NANDX1 G21991 (.A1(W38862), .A2(W9396), .ZN(O16539));
  NANDX1 G21992 (.A1(W22823), .A2(W11942), .ZN(W47584));
  NANDX1 G21993 (.A1(W32912), .A2(W17298), .ZN(O16528));
  NANDX1 G21994 (.A1(W28885), .A2(W25022), .ZN(O16526));
  NANDX1 G21995 (.A1(W38475), .A2(W11053), .ZN(O16525));
  NANDX1 G21996 (.A1(W10505), .A2(W8290), .ZN(O16522));
  NANDX1 G21997 (.A1(W44531), .A2(W6922), .ZN(O16564));
  NANDX1 G21998 (.A1(W3484), .A2(W43395), .ZN(W47565));
  NANDX1 G21999 (.A1(W1242), .A2(I661), .ZN(O16514));
  NANDX1 G22000 (.A1(W45469), .A2(W11223), .ZN(O16512));
  NANDX1 G22001 (.A1(W17101), .A2(W2187), .ZN(O16508));
  NANDX1 G22002 (.A1(W4557), .A2(W23876), .ZN(O16507));
  NANDX1 G22003 (.A1(W47388), .A2(W45832), .ZN(O16506));
  NANDX1 G22004 (.A1(W34526), .A2(I349), .ZN(O16504));
  NANDX1 G22005 (.A1(W12164), .A2(W1532), .ZN(W47539));
  NANDX1 G22006 (.A1(W17192), .A2(W2174), .ZN(O16493));
  NANDX1 G22007 (.A1(W22950), .A2(W8791), .ZN(W47531));
  NANDX1 G22008 (.A1(W13501), .A2(W13895), .ZN(O16488));
  NANDX1 G22009 (.A1(W6023), .A2(W40386), .ZN(O16589));
  NANDX1 G22010 (.A1(W47214), .A2(W3195), .ZN(O16618));
  NANDX1 G22011 (.A1(W11182), .A2(I444), .ZN(O16617));
  NANDX1 G22012 (.A1(W25607), .A2(W7093), .ZN(O16614));
  NANDX1 G22013 (.A1(W28578), .A2(W27130), .ZN(O16612));
  NANDX1 G22014 (.A1(W43386), .A2(W7176), .ZN(W47665));
  NANDX1 G22015 (.A1(W47227), .A2(W33396), .ZN(O16608));
  NANDX1 G22016 (.A1(W12123), .A2(W8771), .ZN(O16607));
  NANDX1 G22017 (.A1(W18622), .A2(W21780), .ZN(O16606));
  NANDX1 G22018 (.A1(W911), .A2(W29855), .ZN(O16605));
  NANDX1 G22019 (.A1(W2587), .A2(W8328), .ZN(O16602));
  NANDX1 G22020 (.A1(W45771), .A2(W24773), .ZN(O16601));
  NANDX1 G22021 (.A1(W32519), .A2(W27702), .ZN(W47649));
  NANDX1 G22022 (.A1(W22130), .A2(W4628), .ZN(O16487));
  NANDX1 G22023 (.A1(W40844), .A2(W26105), .ZN(O16588));
  NANDX1 G22024 (.A1(W18508), .A2(W46573), .ZN(O16585));
  NANDX1 G22025 (.A1(W3105), .A2(W25814), .ZN(O16581));
  NANDX1 G22026 (.A1(W42614), .A2(W7115), .ZN(O16580));
  NANDX1 G22027 (.A1(I227), .A2(W14532), .ZN(O16577));
  NANDX1 G22028 (.A1(W10908), .A2(W19038), .ZN(W47626));
  NANDX1 G22029 (.A1(W4016), .A2(W31629), .ZN(O16576));
  NANDX1 G22030 (.A1(W7774), .A2(W45125), .ZN(O16571));
  NANDX1 G22031 (.A1(W38348), .A2(W29940), .ZN(O16570));
  NANDX1 G22032 (.A1(W27763), .A2(W4162), .ZN(O16565));
  NANDX1 G22033 (.A1(W40524), .A2(W36610), .ZN(W47611));
  NANDX1 G22034 (.A1(W19214), .A2(W1483), .ZN(W47414));
  NANDX1 G22035 (.A1(W6065), .A2(W32780), .ZN(O16416));
  NANDX1 G22036 (.A1(W3638), .A2(W15409), .ZN(O16414));
  NANDX1 G22037 (.A1(W36143), .A2(W12870), .ZN(O16412));
  NANDX1 G22038 (.A1(W5853), .A2(W18905), .ZN(O16411));
  NANDX1 G22039 (.A1(W45758), .A2(W15902), .ZN(O16407));
  NANDX1 G22040 (.A1(W16390), .A2(W12161), .ZN(O16399));
  NANDX1 G22041 (.A1(W38123), .A2(W33216), .ZN(O16398));
  NANDX1 G22042 (.A1(W25447), .A2(W4368), .ZN(O16395));
  NANDX1 G22043 (.A1(W40372), .A2(W24473), .ZN(O16393));
  NANDX1 G22044 (.A1(W26453), .A2(W23905), .ZN(O16389));
  NANDX1 G22045 (.A1(W19864), .A2(W14923), .ZN(O16388));
  NANDX1 G22046 (.A1(I938), .A2(W22405), .ZN(O16387));
  NANDX1 G22047 (.A1(W420), .A2(W43644), .ZN(O16419));
  NANDX1 G22048 (.A1(W8774), .A2(W31703), .ZN(O16383));
  NANDX1 G22049 (.A1(W12394), .A2(W17801), .ZN(O16381));
  NANDX1 G22050 (.A1(W2234), .A2(W2542), .ZN(W47404));
  NANDX1 G22051 (.A1(W19848), .A2(W25485), .ZN(O16373));
  NANDX1 G22052 (.A1(W27346), .A2(W24696), .ZN(O16372));
  NANDX1 G22053 (.A1(W3313), .A2(W20427), .ZN(O16368));
  NANDX1 G22054 (.A1(W45336), .A2(W46005), .ZN(O16366));
  NANDX1 G22055 (.A1(W3456), .A2(W3698), .ZN(O16358));
  NANDX1 G22056 (.A1(W11359), .A2(W42693), .ZN(O16354));
  NANDX1 G22057 (.A1(W14856), .A2(W39263), .ZN(W47375));
  NANDX1 G22058 (.A1(W22526), .A2(W26056), .ZN(O16352));
  NANDX1 G22059 (.A1(W33052), .A2(W25362), .ZN(O16445));
  NANDX1 G22060 (.A1(W15400), .A2(W22614), .ZN(W47514));
  NANDX1 G22061 (.A1(W5214), .A2(W14100), .ZN(W47510));
  NANDX1 G22062 (.A1(W10775), .A2(W35846), .ZN(O16474));
  NANDX1 G22063 (.A1(W2353), .A2(W37021), .ZN(O16470));
  NANDX1 G22064 (.A1(W16349), .A2(W43815), .ZN(O16469));
  NANDX1 G22065 (.A1(W44895), .A2(W6445), .ZN(O16468));
  NANDX1 G22066 (.A1(W42993), .A2(W20621), .ZN(O16464));
  NANDX1 G22067 (.A1(W22573), .A2(W21652), .ZN(O16454));
  NANDX1 G22068 (.A1(W41009), .A2(W38181), .ZN(O16453));
  NANDX1 G22069 (.A1(W18301), .A2(W2958), .ZN(O16450));
  NANDX1 G22070 (.A1(W33093), .A2(W7086), .ZN(O16447));
  NANDX1 G22071 (.A1(W35037), .A2(W6479), .ZN(O16623));
  NANDX1 G22072 (.A1(W8766), .A2(W27670), .ZN(O16443));
  NANDX1 G22073 (.A1(W41829), .A2(W20320), .ZN(O16442));
  NANDX1 G22074 (.A1(W18992), .A2(W16796), .ZN(O16440));
  NANDX1 G22075 (.A1(W7814), .A2(W6986), .ZN(O16439));
  NANDX1 G22076 (.A1(W22732), .A2(W34812), .ZN(O16438));
  NANDX1 G22077 (.A1(W28935), .A2(W17039), .ZN(O16432));
  NANDX1 G22078 (.A1(W29225), .A2(W41974), .ZN(O16429));
  NANDX1 G22079 (.A1(W22446), .A2(W9992), .ZN(W47458));
  NANDX1 G22080 (.A1(W11973), .A2(W21087), .ZN(O16425));
  NANDX1 G22081 (.A1(W3077), .A2(W22269), .ZN(O16423));
  NANDX1 G22082 (.A1(W38031), .A2(W8302), .ZN(O16422));
  NANDX1 G22083 (.A1(W14630), .A2(W20756), .ZN(O16809));
  NANDX1 G22084 (.A1(W26451), .A2(W28261), .ZN(W47919));
  NANDX1 G22085 (.A1(W44478), .A2(W5255), .ZN(O16843));
  NANDX1 G22086 (.A1(W22362), .A2(W37332), .ZN(O16838));
  NANDX1 G22087 (.A1(W30593), .A2(W33888), .ZN(O16833));
  NANDX1 G22088 (.A1(W8307), .A2(W12019), .ZN(O16832));
  NANDX1 G22089 (.A1(W16322), .A2(W18671), .ZN(O16830));
  NANDX1 G22090 (.A1(W38873), .A2(W2750), .ZN(O16827));
  NANDX1 G22091 (.A1(W6304), .A2(W5514), .ZN(O16825));
  NANDX1 G22092 (.A1(W30392), .A2(W18470), .ZN(W47897));
  NANDX1 G22093 (.A1(W23550), .A2(W14257), .ZN(O16820));
  NANDX1 G22094 (.A1(W31184), .A2(W36586), .ZN(O16813));
  NANDX1 G22095 (.A1(W45853), .A2(W35692), .ZN(O16811));
  NANDX1 G22096 (.A1(W36501), .A2(W27165), .ZN(O16848));
  NANDX1 G22097 (.A1(W30768), .A2(W47557), .ZN(O16808));
  NANDX1 G22098 (.A1(W2529), .A2(W39432), .ZN(O16807));
  NANDX1 G22099 (.A1(W33085), .A2(W18101), .ZN(O16803));
  NANDX1 G22100 (.A1(W32608), .A2(W39505), .ZN(O16801));
  NANDX1 G22101 (.A1(W45254), .A2(W8889), .ZN(O16800));
  NANDX1 G22102 (.A1(W39280), .A2(W13654), .ZN(O16798));
  NANDX1 G22103 (.A1(W24163), .A2(W29664), .ZN(W47860));
  NANDX1 G22104 (.A1(W21093), .A2(W31182), .ZN(O16790));
  NANDX1 G22105 (.A1(W28398), .A2(W9082), .ZN(O16789));
  NANDX1 G22106 (.A1(W44096), .A2(W33760), .ZN(O16788));
  NANDX1 G22107 (.A1(W45443), .A2(W15667), .ZN(W47854));
  NANDX1 G22108 (.A1(W43682), .A2(W7094), .ZN(O16886));
  NANDX1 G22109 (.A1(I1284), .A2(W2040), .ZN(O16911));
  NANDX1 G22110 (.A1(W23769), .A2(W15819), .ZN(O16909));
  NANDX1 G22111 (.A1(W2110), .A2(W28172), .ZN(O16908));
  NANDX1 G22112 (.A1(W1226), .A2(I562), .ZN(O16906));
  NANDX1 G22113 (.A1(W21468), .A2(W38890), .ZN(O16900));
  NANDX1 G22114 (.A1(W25687), .A2(W20429), .ZN(O16898));
  NANDX1 G22115 (.A1(W18805), .A2(W14484), .ZN(O16897));
  NANDX1 G22116 (.A1(W43103), .A2(W7236), .ZN(O16895));
  NANDX1 G22117 (.A1(W31855), .A2(W26722), .ZN(O16894));
  NANDX1 G22118 (.A1(W26815), .A2(W2885), .ZN(O16890));
  NANDX1 G22119 (.A1(W22833), .A2(W5261), .ZN(O16889));
  NANDX1 G22120 (.A1(W18017), .A2(W22853), .ZN(O16774));
  NANDX1 G22121 (.A1(W39674), .A2(W42147), .ZN(O16882));
  NANDX1 G22122 (.A1(W32169), .A2(W16031), .ZN(O16881));
  NANDX1 G22123 (.A1(W4943), .A2(I856), .ZN(O16873));
  NANDX1 G22124 (.A1(W9589), .A2(W16861), .ZN(O16870));
  NANDX1 G22125 (.A1(W46841), .A2(W1015), .ZN(O16865));
  NANDX1 G22126 (.A1(W5876), .A2(W22729), .ZN(O16863));
  NANDX1 G22127 (.A1(W11536), .A2(W43652), .ZN(O16861));
  NANDX1 G22128 (.A1(W14483), .A2(W33724), .ZN(W47933));
  NANDX1 G22129 (.A1(W11519), .A2(W38897), .ZN(O16857));
  NANDX1 G22130 (.A1(W28829), .A2(W1267), .ZN(O16856));
  NANDX1 G22131 (.A1(W21489), .A2(W46709), .ZN(O16853));
  NANDX1 G22132 (.A1(W45988), .A2(W18760), .ZN(O16652));
  NANDX1 G22133 (.A1(W29822), .A2(W42723), .ZN(O16687));
  NANDX1 G22134 (.A1(W4510), .A2(W19531), .ZN(O16684));
  NANDX1 G22135 (.A1(W34600), .A2(W13901), .ZN(O16683));
  NANDX1 G22136 (.A1(W39052), .A2(W7565), .ZN(O16677));
  NANDX1 G22137 (.A1(W34120), .A2(W39258), .ZN(O16676));
  NANDX1 G22138 (.A1(W3047), .A2(W45468), .ZN(O16673));
  NANDX1 G22139 (.A1(W11477), .A2(W17456), .ZN(O16670));
  NANDX1 G22140 (.A1(W9387), .A2(W31562), .ZN(O16669));
  NANDX1 G22141 (.A1(I676), .A2(W11416), .ZN(O16664));
  NANDX1 G22142 (.A1(W36278), .A2(W1098), .ZN(O16658));
  NANDX1 G22143 (.A1(W1990), .A2(W5952), .ZN(O16657));
  NANDX1 G22144 (.A1(W33766), .A2(W45234), .ZN(O16655));
  NANDX1 G22145 (.A1(W39127), .A2(W38036), .ZN(O16690));
  NANDX1 G22146 (.A1(W41539), .A2(I1038), .ZN(O16647));
  NANDX1 G22147 (.A1(W21201), .A2(W14634), .ZN(O16644));
  NANDX1 G22148 (.A1(W40569), .A2(W8796), .ZN(O16642));
  NANDX1 G22149 (.A1(W33992), .A2(W20451), .ZN(O16641));
  NANDX1 G22150 (.A1(W33547), .A2(W44748), .ZN(O16638));
  NANDX1 G22151 (.A1(W42733), .A2(W42595), .ZN(O16635));
  NANDX1 G22152 (.A1(W14660), .A2(W26039), .ZN(O16634));
  NANDX1 G22153 (.A1(W25045), .A2(W15399), .ZN(W47689));
  NANDX1 G22154 (.A1(W12359), .A2(W4900), .ZN(O16631));
  NANDX1 G22155 (.A1(W26518), .A2(W42527), .ZN(O16629));
  NANDX1 G22156 (.A1(W11739), .A2(W20911), .ZN(O16628));
  NANDX1 G22157 (.A1(W27943), .A2(W23307), .ZN(O16739));
  NANDX1 G22158 (.A1(W3225), .A2(W3211), .ZN(O16770));
  NANDX1 G22159 (.A1(W34372), .A2(W40646), .ZN(O16769));
  NANDX1 G22160 (.A1(W17503), .A2(W36595), .ZN(O16763));
  NANDX1 G22161 (.A1(W585), .A2(W30464), .ZN(W47824));
  NANDX1 G22162 (.A1(W36302), .A2(I271), .ZN(O16759));
  NANDX1 G22163 (.A1(W38887), .A2(W38572), .ZN(O16757));
  NANDX1 G22164 (.A1(W4003), .A2(W16248), .ZN(O16756));
  NANDX1 G22165 (.A1(W29050), .A2(W14509), .ZN(O16753));
  NANDX1 G22166 (.A1(W40322), .A2(W33386), .ZN(O16747));
  NANDX1 G22167 (.A1(W12802), .A2(W14346), .ZN(O16744));
  NANDX1 G22168 (.A1(W27796), .A2(W40450), .ZN(O16742));
  NANDX1 G22169 (.A1(W5816), .A2(W14860), .ZN(O11670));
  NANDX1 G22170 (.A1(W25688), .A2(W5875), .ZN(O16735));
  NANDX1 G22171 (.A1(W38353), .A2(W18391), .ZN(O16732));
  NANDX1 G22172 (.A1(W4726), .A2(W40867), .ZN(O16729));
  NANDX1 G22173 (.A1(W32189), .A2(W11362), .ZN(O16722));
  NANDX1 G22174 (.A1(W33281), .A2(W20364), .ZN(O16721));
  NANDX1 G22175 (.A1(W17652), .A2(W12930), .ZN(O16720));
  NANDX1 G22176 (.A1(W3887), .A2(W35422), .ZN(O16717));
  NANDX1 G22177 (.A1(W32936), .A2(W7879), .ZN(O16714));
  NANDX1 G22178 (.A1(W14832), .A2(W45715), .ZN(W47768));
  NANDX1 G22179 (.A1(W2695), .A2(W26244), .ZN(O16698));
  NANDX1 G22180 (.A1(W41751), .A2(W33033), .ZN(O16695));
  NANDX1 G22181 (.A1(W17568), .A2(W25837), .ZN(W34941));
  NANDX1 G22182 (.A1(W3851), .A2(W20466), .ZN(W34963));
  NANDX1 G22183 (.A1(I928), .A2(W28405), .ZN(O7538));
  NANDX1 G22184 (.A1(W34647), .A2(W31742), .ZN(W34957));
  NANDX1 G22185 (.A1(W6490), .A2(W15628), .ZN(W34956));
  NANDX1 G22186 (.A1(W19835), .A2(W14908), .ZN(O7535));
  NANDX1 G22187 (.A1(W23990), .A2(W12218), .ZN(O7534));
  NANDX1 G22188 (.A1(W26284), .A2(W26694), .ZN(W34952));
  NANDX1 G22189 (.A1(W26510), .A2(W31078), .ZN(O7532));
  NANDX1 G22190 (.A1(W7029), .A2(W19051), .ZN(W34948));
  NANDX1 G22191 (.A1(W34646), .A2(W17461), .ZN(W34947));
  NANDX1 G22192 (.A1(W17890), .A2(W25675), .ZN(O7531));
  NANDX1 G22193 (.A1(W8723), .A2(I609), .ZN(O7529));
  NANDX1 G22194 (.A1(W14523), .A2(W8730), .ZN(O7539));
  NANDX1 G22195 (.A1(W3605), .A2(W68), .ZN(W34939));
  NANDX1 G22196 (.A1(W18997), .A2(W20751), .ZN(W34937));
  NANDX1 G22197 (.A1(W34419), .A2(W15899), .ZN(O7526));
  NANDX1 G22198 (.A1(W16869), .A2(W22388), .ZN(O7525));
  NANDX1 G22199 (.A1(W20905), .A2(W26960), .ZN(W34932));
  NANDX1 G22200 (.A1(W26991), .A2(W21230), .ZN(O7523));
  NANDX1 G22201 (.A1(W407), .A2(I448), .ZN(O7520));
  NANDX1 G22202 (.A1(W27057), .A2(I1088), .ZN(O7517));
  NANDX1 G22203 (.A1(W34801), .A2(W8619), .ZN(W34921));
  NANDX1 G22204 (.A1(W11734), .A2(W25040), .ZN(O7512));
  NANDX1 G22205 (.A1(W10812), .A2(W34362), .ZN(O7511));
  NANDX1 G22206 (.A1(W17217), .A2(W11798), .ZN(O7575));
  NANDX1 G22207 (.A1(W30876), .A2(W33745), .ZN(W35042));
  NANDX1 G22208 (.A1(W5582), .A2(W8983), .ZN(W35041));
  NANDX1 G22209 (.A1(W23412), .A2(W28541), .ZN(O7587));
  NANDX1 G22210 (.A1(W15563), .A2(W8563), .ZN(W35035));
  NANDX1 G22211 (.A1(W12724), .A2(W22496), .ZN(O7586));
  NANDX1 G22212 (.A1(W25793), .A2(W791), .ZN(W35033));
  NANDX1 G22213 (.A1(W27129), .A2(W24114), .ZN(O7584));
  NANDX1 G22214 (.A1(W7151), .A2(I286), .ZN(O7581));
  NANDX1 G22215 (.A1(W10960), .A2(W29334), .ZN(O7580));
  NANDX1 G22216 (.A1(W4928), .A2(W14149), .ZN(O7579));
  NANDX1 G22217 (.A1(W23079), .A2(W15235), .ZN(W35019));
  NANDX1 G22218 (.A1(W22584), .A2(W22530), .ZN(W35016));
  NANDX1 G22219 (.A1(W2407), .A2(W24762), .ZN(O7507));
  NANDX1 G22220 (.A1(W25067), .A2(W34078), .ZN(O7574));
  NANDX1 G22221 (.A1(W21493), .A2(W19857), .ZN(O7573));
  NANDX1 G22222 (.A1(W12911), .A2(W29284), .ZN(O7568));
  NANDX1 G22223 (.A1(W11730), .A2(W4000), .ZN(O7566));
  NANDX1 G22224 (.A1(W34683), .A2(W32363), .ZN(O7565));
  NANDX1 G22225 (.A1(W20577), .A2(W11160), .ZN(W34999));
  NANDX1 G22226 (.A1(W21914), .A2(W33788), .ZN(O7559));
  NANDX1 G22227 (.A1(W31742), .A2(W194), .ZN(O7554));
  NANDX1 G22228 (.A1(W20858), .A2(W15037), .ZN(O7551));
  NANDX1 G22229 (.A1(W2016), .A2(W15762), .ZN(O7544));
  NANDX1 G22230 (.A1(W32882), .A2(W8390), .ZN(W34968));
  NANDX1 G22231 (.A1(W30516), .A2(W28628), .ZN(O7446));
  NANDX1 G22232 (.A1(W29691), .A2(W13283), .ZN(O7458));
  NANDX1 G22233 (.A1(W1795), .A2(W13024), .ZN(W34810));
  NANDX1 G22234 (.A1(W26442), .A2(W20440), .ZN(W34807));
  NANDX1 G22235 (.A1(W22845), .A2(W10762), .ZN(O7457));
  NANDX1 G22236 (.A1(W7172), .A2(W12569), .ZN(O7455));
  NANDX1 G22237 (.A1(W31592), .A2(W11166), .ZN(W34801));
  NANDX1 G22238 (.A1(W32733), .A2(W11495), .ZN(W34794));
  NANDX1 G22239 (.A1(W29922), .A2(W28869), .ZN(O7451));
  NANDX1 G22240 (.A1(W18649), .A2(W3933), .ZN(O7450));
  NANDX1 G22241 (.A1(W18973), .A2(W31580), .ZN(W34789));
  NANDX1 G22242 (.A1(W6665), .A2(W28798), .ZN(O7449));
  NANDX1 G22243 (.A1(W9254), .A2(W31313), .ZN(W34784));
  NANDX1 G22244 (.A1(W4882), .A2(W30913), .ZN(O7464));
  NANDX1 G22245 (.A1(W33715), .A2(W29659), .ZN(O7444));
  NANDX1 G22246 (.A1(W24444), .A2(W30322), .ZN(O7440));
  NANDX1 G22247 (.A1(W18691), .A2(W24078), .ZN(O7438));
  NANDX1 G22248 (.A1(W17818), .A2(W7638), .ZN(W34768));
  NANDX1 G22249 (.A1(W16341), .A2(W21841), .ZN(W34767));
  NANDX1 G22250 (.A1(I1422), .A2(W32368), .ZN(O7435));
  NANDX1 G22251 (.A1(W8684), .A2(W756), .ZN(O7434));
  NANDX1 G22252 (.A1(W7292), .A2(W17695), .ZN(O7433));
  NANDX1 G22253 (.A1(I1427), .A2(W22829), .ZN(W34752));
  NANDX1 G22254 (.A1(W11509), .A2(W34339), .ZN(W34743));
  NANDX1 G22255 (.A1(W29298), .A2(W8706), .ZN(O7424));
  NANDX1 G22256 (.A1(W9255), .A2(W11292), .ZN(O7486));
  NANDX1 G22257 (.A1(W19413), .A2(W12056), .ZN(O7506));
  NANDX1 G22258 (.A1(W26014), .A2(W29796), .ZN(O7504));
  NANDX1 G22259 (.A1(W14722), .A2(W7635), .ZN(O7498));
  NANDX1 G22260 (.A1(W10561), .A2(W16239), .ZN(W34892));
  NANDX1 G22261 (.A1(W30040), .A2(W15439), .ZN(W34890));
  NANDX1 G22262 (.A1(W11182), .A2(W2418), .ZN(W34885));
  NANDX1 G22263 (.A1(W24885), .A2(W20979), .ZN(W34883));
  NANDX1 G22264 (.A1(W4695), .A2(W18897), .ZN(W34878));
  NANDX1 G22265 (.A1(I1060), .A2(W2255), .ZN(O7490));
  NANDX1 G22266 (.A1(W25926), .A2(W20709), .ZN(O7488));
  NANDX1 G22267 (.A1(W11430), .A2(W30652), .ZN(W34865));
  NANDX1 G22268 (.A1(W22355), .A2(W12485), .ZN(O7589));
  NANDX1 G22269 (.A1(W13628), .A2(I1831), .ZN(O7485));
  NANDX1 G22270 (.A1(W22034), .A2(W4731), .ZN(O7484));
  NANDX1 G22271 (.A1(W18039), .A2(W16047), .ZN(W34850));
  NANDX1 G22272 (.A1(W22342), .A2(W17172), .ZN(W34848));
  NANDX1 G22273 (.A1(W19908), .A2(W8877), .ZN(W34844));
  NANDX1 G22274 (.A1(W34640), .A2(W20423), .ZN(W34841));
  NANDX1 G22275 (.A1(W1603), .A2(W24987), .ZN(O7472));
  NANDX1 G22276 (.A1(W4548), .A2(W1944), .ZN(W34834));
  NANDX1 G22277 (.A1(W7187), .A2(W13365), .ZN(W34828));
  NANDX1 G22278 (.A1(I43), .A2(W11652), .ZN(O7469));
  NANDX1 G22279 (.A1(W1699), .A2(W609), .ZN(W34822));
  NANDX1 G22280 (.A1(W27769), .A2(W27505), .ZN(W35204));
  NANDX1 G22281 (.A1(W21452), .A2(W34992), .ZN(W35247));
  NANDX1 G22282 (.A1(W17699), .A2(W22912), .ZN(O7692));
  NANDX1 G22283 (.A1(W7902), .A2(W11332), .ZN(W35243));
  NANDX1 G22284 (.A1(W34109), .A2(W33216), .ZN(W35234));
  NANDX1 G22285 (.A1(W5006), .A2(W20887), .ZN(W35228));
  NANDX1 G22286 (.A1(W5996), .A2(W12956), .ZN(O7685));
  NANDX1 G22287 (.A1(W2267), .A2(W1340), .ZN(W35225));
  NANDX1 G22288 (.A1(W22225), .A2(W2311), .ZN(W35224));
  NANDX1 G22289 (.A1(W17834), .A2(W81), .ZN(W35215));
  NANDX1 G22290 (.A1(W6349), .A2(W20543), .ZN(O7679));
  NANDX1 G22291 (.A1(W9472), .A2(W7170), .ZN(O7678));
  NANDX1 G22292 (.A1(W31078), .A2(W399), .ZN(O7677));
  NANDX1 G22293 (.A1(W31288), .A2(W12277), .ZN(O7697));
  NANDX1 G22294 (.A1(W19490), .A2(W9870), .ZN(O7674));
  NANDX1 G22295 (.A1(W34852), .A2(W281), .ZN(W35199));
  NANDX1 G22296 (.A1(W31068), .A2(W14513), .ZN(W35198));
  NANDX1 G22297 (.A1(W9205), .A2(I290), .ZN(W35194));
  NANDX1 G22298 (.A1(W27785), .A2(W16577), .ZN(O7671));
  NANDX1 G22299 (.A1(W17249), .A2(W3019), .ZN(O7668));
  NANDX1 G22300 (.A1(I635), .A2(W16149), .ZN(O7667));
  NANDX1 G22301 (.A1(I977), .A2(W28060), .ZN(W35185));
  NANDX1 G22302 (.A1(I1556), .A2(W1186), .ZN(O7666));
  NANDX1 G22303 (.A1(W21001), .A2(W3809), .ZN(O7662));
  NANDX1 G22304 (.A1(W13401), .A2(W7735), .ZN(W35177));
  NANDX1 G22305 (.A1(W590), .A2(W21689), .ZN(O7711));
  NANDX1 G22306 (.A1(W10948), .A2(W1608), .ZN(O7742));
  NANDX1 G22307 (.A1(W11622), .A2(W33483), .ZN(O7740));
  NANDX1 G22308 (.A1(W30065), .A2(W2889), .ZN(W35312));
  NANDX1 G22309 (.A1(W27771), .A2(W6363), .ZN(O7728));
  NANDX1 G22310 (.A1(W7192), .A2(W10402), .ZN(O7723));
  NANDX1 G22311 (.A1(W16360), .A2(W15720), .ZN(O7722));
  NANDX1 G22312 (.A1(W15557), .A2(W29804), .ZN(O7718));
  NANDX1 G22313 (.A1(W27239), .A2(I1103), .ZN(O7717));
  NANDX1 G22314 (.A1(W18668), .A2(W33061), .ZN(W35282));
  NANDX1 G22315 (.A1(W24231), .A2(W33078), .ZN(W35281));
  NANDX1 G22316 (.A1(W5421), .A2(W34638), .ZN(O7713));
  NANDX1 G22317 (.A1(W27668), .A2(W7369), .ZN(O7712));
  NANDX1 G22318 (.A1(W17504), .A2(W18909), .ZN(W35174));
  NANDX1 G22319 (.A1(W8783), .A2(W17193), .ZN(W35276));
  NANDX1 G22320 (.A1(W29384), .A2(W9925), .ZN(O7708));
  NANDX1 G22321 (.A1(W8803), .A2(W4903), .ZN(O7707));
  NANDX1 G22322 (.A1(W17137), .A2(W24397), .ZN(O7706));
  NANDX1 G22323 (.A1(W12922), .A2(W28018), .ZN(O7705));
  NANDX1 G22324 (.A1(W20098), .A2(W175), .ZN(O7704));
  NANDX1 G22325 (.A1(W27508), .A2(W3112), .ZN(W35265));
  NANDX1 G22326 (.A1(W8177), .A2(I534), .ZN(O7702));
  NANDX1 G22327 (.A1(W10433), .A2(W23170), .ZN(W35260));
  NANDX1 G22328 (.A1(W20040), .A2(W35248), .ZN(O7699));
  NANDX1 G22329 (.A1(W32042), .A2(W22872), .ZN(W35255));
  NANDX1 G22330 (.A1(W3437), .A2(W23557), .ZN(W35077));
  NANDX1 G22331 (.A1(W7567), .A2(W24098), .ZN(O7627));
  NANDX1 G22332 (.A1(W17666), .A2(W13899), .ZN(W35105));
  NANDX1 G22333 (.A1(W12217), .A2(W27210), .ZN(O7626));
  NANDX1 G22334 (.A1(W37), .A2(W28463), .ZN(W35101));
  NANDX1 G22335 (.A1(W34578), .A2(W5795), .ZN(W35100));
  NANDX1 G22336 (.A1(W20023), .A2(W23694), .ZN(O7623));
  NANDX1 G22337 (.A1(W17128), .A2(W33856), .ZN(W35088));
  NANDX1 G22338 (.A1(I1188), .A2(W11882), .ZN(W35087));
  NANDX1 G22339 (.A1(W24099), .A2(W4316), .ZN(O7617));
  NANDX1 G22340 (.A1(W35065), .A2(W13721), .ZN(O7616));
  NANDX1 G22341 (.A1(W13971), .A2(W15354), .ZN(W35084));
  NANDX1 G22342 (.A1(W20027), .A2(W21923), .ZN(O7613));
  NANDX1 G22343 (.A1(W18256), .A2(W7801), .ZN(W35114));
  NANDX1 G22344 (.A1(W32528), .A2(W15453), .ZN(W35074));
  NANDX1 G22345 (.A1(W15708), .A2(W28536), .ZN(O7603));
  NANDX1 G22346 (.A1(W25669), .A2(W21265), .ZN(W35063));
  NANDX1 G22347 (.A1(W17394), .A2(W20562), .ZN(O7602));
  NANDX1 G22348 (.A1(W13914), .A2(W27437), .ZN(O7600));
  NANDX1 G22349 (.A1(W28874), .A2(W1838), .ZN(W35059));
  NANDX1 G22350 (.A1(W8689), .A2(W5644), .ZN(O7599));
  NANDX1 G22351 (.A1(W27505), .A2(W33890), .ZN(W35054));
  NANDX1 G22352 (.A1(W11085), .A2(W5438), .ZN(O7593));
  NANDX1 G22353 (.A1(W9429), .A2(W24356), .ZN(O7592));
  NANDX1 G22354 (.A1(W13841), .A2(I1575), .ZN(O7590));
  NANDX1 G22355 (.A1(W28428), .A2(W13730), .ZN(W35144));
  NANDX1 G22356 (.A1(W10881), .A2(W8853), .ZN(W35172));
  NANDX1 G22357 (.A1(W10974), .A2(W8536), .ZN(O7660));
  NANDX1 G22358 (.A1(W22211), .A2(W5002), .ZN(O7658));
  NANDX1 G22359 (.A1(W2104), .A2(W2408), .ZN(W35166));
  NANDX1 G22360 (.A1(W29657), .A2(W6640), .ZN(O7656));
  NANDX1 G22361 (.A1(W17220), .A2(W25712), .ZN(W35160));
  NANDX1 G22362 (.A1(W9990), .A2(W35042), .ZN(W35158));
  NANDX1 G22363 (.A1(W25804), .A2(W3097), .ZN(W35155));
  NANDX1 G22364 (.A1(W4613), .A2(W3254), .ZN(O7647));
  NANDX1 G22365 (.A1(W18573), .A2(W15009), .ZN(O7646));
  NANDX1 G22366 (.A1(W423), .A2(W26092), .ZN(W35146));
  NANDX1 G22367 (.A1(W17574), .A2(W29769), .ZN(O7418));
  NANDX1 G22368 (.A1(W33168), .A2(W31855), .ZN(W35139));
  NANDX1 G22369 (.A1(I520), .A2(W20614), .ZN(W35138));
  NANDX1 G22370 (.A1(W9697), .A2(W25611), .ZN(W35134));
  NANDX1 G22371 (.A1(W29154), .A2(W23679), .ZN(W35133));
  NANDX1 G22372 (.A1(W5790), .A2(W30684), .ZN(W35130));
  NANDX1 G22373 (.A1(W4036), .A2(W35012), .ZN(W35129));
  NANDX1 G22374 (.A1(W4309), .A2(W34153), .ZN(O7642));
  NANDX1 G22375 (.A1(W27310), .A2(W24487), .ZN(O7640));
  NANDX1 G22376 (.A1(W26998), .A2(W9448), .ZN(O7639));
  NANDX1 G22377 (.A1(W12885), .A2(W9177), .ZN(O7638));
  NANDX1 G22378 (.A1(W7641), .A2(W20155), .ZN(O7634));
  NANDX1 G22379 (.A1(W14041), .A2(W26060), .ZN(W34366));
  NANDX1 G22380 (.A1(W31335), .A2(W13065), .ZN(W34392));
  NANDX1 G22381 (.A1(W31637), .A2(W29402), .ZN(O7227));
  NANDX1 G22382 (.A1(W6753), .A2(W18810), .ZN(W34387));
  NANDX1 G22383 (.A1(W9525), .A2(W14897), .ZN(W34384));
  NANDX1 G22384 (.A1(W3966), .A2(W11329), .ZN(O7220));
  NANDX1 G22385 (.A1(W20318), .A2(W24759), .ZN(W34379));
  NANDX1 G22386 (.A1(W5417), .A2(W22523), .ZN(W34376));
  NANDX1 G22387 (.A1(W24933), .A2(W3539), .ZN(O7219));
  NANDX1 G22388 (.A1(W20820), .A2(W28029), .ZN(O7218));
  NANDX1 G22389 (.A1(W6725), .A2(W18002), .ZN(W34372));
  NANDX1 G22390 (.A1(W18922), .A2(W29688), .ZN(O7217));
  NANDX1 G22391 (.A1(W7142), .A2(W25298), .ZN(O7215));
  NANDX1 G22392 (.A1(W4567), .A2(W23919), .ZN(O7229));
  NANDX1 G22393 (.A1(W8334), .A2(W29138), .ZN(W34362));
  NANDX1 G22394 (.A1(W25854), .A2(W18382), .ZN(O7211));
  NANDX1 G22395 (.A1(W24257), .A2(W5187), .ZN(O7210));
  NANDX1 G22396 (.A1(I214), .A2(W15940), .ZN(W34356));
  NANDX1 G22397 (.A1(W9441), .A2(W21071), .ZN(W34355));
  NANDX1 G22398 (.A1(W18911), .A2(W5447), .ZN(O7207));
  NANDX1 G22399 (.A1(W33075), .A2(W33488), .ZN(O7204));
  NANDX1 G22400 (.A1(W13969), .A2(W11410), .ZN(W34343));
  NANDX1 G22401 (.A1(W28761), .A2(W30291), .ZN(O7202));
  NANDX1 G22402 (.A1(W23084), .A2(W22909), .ZN(W34339));
  NANDX1 G22403 (.A1(W11623), .A2(W18439), .ZN(O7198));
  NANDX1 G22404 (.A1(W26230), .A2(W31353), .ZN(O7241));
  NANDX1 G22405 (.A1(W26548), .A2(W9053), .ZN(W34450));
  NANDX1 G22406 (.A1(W21900), .A2(W33657), .ZN(W34447));
  NANDX1 G22407 (.A1(W20662), .A2(W8277), .ZN(O7261));
  NANDX1 G22408 (.A1(W7500), .A2(W17345), .ZN(O7260));
  NANDX1 G22409 (.A1(W3269), .A2(W27421), .ZN(O7259));
  NANDX1 G22410 (.A1(W8810), .A2(W18822), .ZN(O7257));
  NANDX1 G22411 (.A1(W27701), .A2(W15706), .ZN(O7254));
  NANDX1 G22412 (.A1(W22860), .A2(W20410), .ZN(O7253));
  NANDX1 G22413 (.A1(W31479), .A2(W8736), .ZN(O7248));
  NANDX1 G22414 (.A1(W6832), .A2(W6648), .ZN(O7245));
  NANDX1 G22415 (.A1(W32468), .A2(W27831), .ZN(O7244));
  NANDX1 G22416 (.A1(W5350), .A2(W5525), .ZN(W34417));
  NANDX1 G22417 (.A1(W23998), .A2(W26569), .ZN(W34330));
  NANDX1 G22418 (.A1(W17546), .A2(W12544), .ZN(W34412));
  NANDX1 G22419 (.A1(W18878), .A2(W13969), .ZN(O7240));
  NANDX1 G22420 (.A1(W8897), .A2(I1725), .ZN(W34410));
  NANDX1 G22421 (.A1(W6573), .A2(W31241), .ZN(W34408));
  NANDX1 G22422 (.A1(W26573), .A2(W25696), .ZN(O7237));
  NANDX1 G22423 (.A1(W5698), .A2(W29402), .ZN(W34404));
  NANDX1 G22424 (.A1(W13158), .A2(W7610), .ZN(O7235));
  NANDX1 G22425 (.A1(W19036), .A2(W419), .ZN(O7234));
  NANDX1 G22426 (.A1(W27814), .A2(W22027), .ZN(W34400));
  NANDX1 G22427 (.A1(W5953), .A2(W5886), .ZN(O7233));
  NANDX1 G22428 (.A1(W24847), .A2(W12850), .ZN(W34395));
  NANDX1 G22429 (.A1(W31401), .A2(W33327), .ZN(O7139));
  NANDX1 G22430 (.A1(W14684), .A2(I1092), .ZN(W34261));
  NANDX1 G22431 (.A1(W2943), .A2(W558), .ZN(W34260));
  NANDX1 G22432 (.A1(W34100), .A2(W20462), .ZN(W34257));
  NANDX1 G22433 (.A1(W8150), .A2(W18532), .ZN(W34255));
  NANDX1 G22434 (.A1(W6299), .A2(W26233), .ZN(W34254));
  NANDX1 G22435 (.A1(W895), .A2(W5102), .ZN(O7154));
  NANDX1 G22436 (.A1(W7926), .A2(W27738), .ZN(O7153));
  NANDX1 G22437 (.A1(W26638), .A2(W9217), .ZN(W34248));
  NANDX1 G22438 (.A1(W7385), .A2(W154), .ZN(O7150));
  NANDX1 G22439 (.A1(W4828), .A2(I1290), .ZN(O7149));
  NANDX1 G22440 (.A1(W20501), .A2(I604), .ZN(W34238));
  NANDX1 G22441 (.A1(W21430), .A2(W3187), .ZN(O7141));
  NANDX1 G22442 (.A1(W14836), .A2(W17578), .ZN(W34264));
  NANDX1 G22443 (.A1(W13797), .A2(W19312), .ZN(W34230));
  NANDX1 G22444 (.A1(W11884), .A2(W4611), .ZN(O7136));
  NANDX1 G22445 (.A1(W11781), .A2(W3857), .ZN(O7135));
  NANDX1 G22446 (.A1(W16413), .A2(W26838), .ZN(O7133));
  NANDX1 G22447 (.A1(W2303), .A2(W10669), .ZN(O7132));
  NANDX1 G22448 (.A1(W12023), .A2(W29981), .ZN(O7131));
  NANDX1 G22449 (.A1(W34091), .A2(W6289), .ZN(W34219));
  NANDX1 G22450 (.A1(W34041), .A2(W20860), .ZN(O7128));
  NANDX1 G22451 (.A1(W19140), .A2(W1712), .ZN(W34211));
  NANDX1 G22452 (.A1(W26454), .A2(W17010), .ZN(W34207));
  NANDX1 G22453 (.A1(W28133), .A2(W14526), .ZN(W34205));
  NANDX1 G22454 (.A1(W24571), .A2(W33494), .ZN(W34302));
  NANDX1 G22455 (.A1(W34177), .A2(W27892), .ZN(W34326));
  NANDX1 G22456 (.A1(W17068), .A2(W1052), .ZN(W34322));
  NANDX1 G22457 (.A1(W1092), .A2(W21278), .ZN(W34320));
  NANDX1 G22458 (.A1(W32972), .A2(W15161), .ZN(O7193));
  NANDX1 G22459 (.A1(W21656), .A2(W22535), .ZN(O7192));
  NANDX1 G22460 (.A1(W7585), .A2(W18103), .ZN(W34317));
  NANDX1 G22461 (.A1(W4264), .A2(W20439), .ZN(W34309));
  NANDX1 G22462 (.A1(W1588), .A2(W25579), .ZN(O7186));
  NANDX1 G22463 (.A1(W17324), .A2(W5268), .ZN(O7185));
  NANDX1 G22464 (.A1(W26282), .A2(W16220), .ZN(O7184));
  NANDX1 G22465 (.A1(W15205), .A2(W9227), .ZN(W34303));
  NANDX1 G22466 (.A1(W17833), .A2(W31115), .ZN(O7263));
  NANDX1 G22467 (.A1(W29957), .A2(W31265), .ZN(O7183));
  NANDX1 G22468 (.A1(W16524), .A2(W6798), .ZN(O7181));
  NANDX1 G22469 (.A1(W2636), .A2(I1425), .ZN(O7179));
  NANDX1 G22470 (.A1(W27800), .A2(W19115), .ZN(O7173));
  NANDX1 G22471 (.A1(W32492), .A2(W1288), .ZN(O7172));
  NANDX1 G22472 (.A1(W24316), .A2(W5059), .ZN(W34288));
  NANDX1 G22473 (.A1(W26138), .A2(W28632), .ZN(O7161));
  NANDX1 G22474 (.A1(W26374), .A2(W22619), .ZN(O7160));
  NANDX1 G22475 (.A1(W24465), .A2(I1646), .ZN(W34273));
  NANDX1 G22476 (.A1(W9492), .A2(W3735), .ZN(O7158));
  NANDX1 G22477 (.A1(W10204), .A2(W1924), .ZN(O7157));
  NANDX1 G22478 (.A1(W17822), .A2(W16244), .ZN(W34622));
  NANDX1 G22479 (.A1(W14211), .A2(W18231), .ZN(W34646));
  NANDX1 G22480 (.A1(W5819), .A2(I887), .ZN(O7371));
  NANDX1 G22481 (.A1(W30770), .A2(W12414), .ZN(W34642));
  NANDX1 G22482 (.A1(W24788), .A2(W2238), .ZN(W34640));
  NANDX1 G22483 (.A1(W29245), .A2(W16992), .ZN(O7369));
  NANDX1 G22484 (.A1(W8775), .A2(W29302), .ZN(O7366));
  NANDX1 G22485 (.A1(W25838), .A2(W25923), .ZN(W34632));
  NANDX1 G22486 (.A1(W28327), .A2(W4699), .ZN(O7364));
  NANDX1 G22487 (.A1(W28702), .A2(W32103), .ZN(O7363));
  NANDX1 G22488 (.A1(W16997), .A2(W32970), .ZN(O7362));
  NANDX1 G22489 (.A1(W3208), .A2(W18819), .ZN(W34626));
  NANDX1 G22490 (.A1(W16869), .A2(W8026), .ZN(W34625));
  NANDX1 G22491 (.A1(W31441), .A2(W18702), .ZN(W34647));
  NANDX1 G22492 (.A1(W886), .A2(W32565), .ZN(O7360));
  NANDX1 G22493 (.A1(W32065), .A2(W31994), .ZN(O7359));
  NANDX1 G22494 (.A1(W27026), .A2(W29087), .ZN(O7357));
  NANDX1 G22495 (.A1(W574), .A2(W31482), .ZN(O7356));
  NANDX1 G22496 (.A1(W30590), .A2(W3156), .ZN(W34612));
  NANDX1 G22497 (.A1(W18208), .A2(W15458), .ZN(O7346));
  NANDX1 G22498 (.A1(W1545), .A2(W8890), .ZN(W34596));
  NANDX1 G22499 (.A1(W23389), .A2(W19381), .ZN(O7345));
  NANDX1 G22500 (.A1(W2370), .A2(W12190), .ZN(W34594));
  NANDX1 G22501 (.A1(W1878), .A2(W14265), .ZN(W34593));
  NANDX1 G22502 (.A1(W33362), .A2(W6340), .ZN(O7344));
  NANDX1 G22503 (.A1(W23685), .A2(I386), .ZN(W34674));
  NANDX1 G22504 (.A1(W20151), .A2(W25553), .ZN(O7416));
  NANDX1 G22505 (.A1(W20794), .A2(W33263), .ZN(O7408));
  NANDX1 G22506 (.A1(W9661), .A2(W32685), .ZN(O7407));
  NANDX1 G22507 (.A1(W3603), .A2(W20908), .ZN(O7404));
  NANDX1 G22508 (.A1(W25008), .A2(W15221), .ZN(O7403));
  NANDX1 G22509 (.A1(W28551), .A2(W30232), .ZN(W34702));
  NANDX1 G22510 (.A1(W17238), .A2(W33099), .ZN(O7399));
  NANDX1 G22511 (.A1(W21988), .A2(W34543), .ZN(W34696));
  NANDX1 G22512 (.A1(W6118), .A2(W8819), .ZN(W34694));
  NANDX1 G22513 (.A1(W14507), .A2(W500), .ZN(W34692));
  NANDX1 G22514 (.A1(W4377), .A2(W5588), .ZN(W34688));
  NANDX1 G22515 (.A1(W3932), .A2(W32593), .ZN(O7390));
  NANDX1 G22516 (.A1(W19207), .A2(I1994), .ZN(O7343));
  NANDX1 G22517 (.A1(W6880), .A2(W8219), .ZN(O7388));
  NANDX1 G22518 (.A1(W32411), .A2(W17893), .ZN(W34672));
  NANDX1 G22519 (.A1(I1218), .A2(W12836), .ZN(W34667));
  NANDX1 G22520 (.A1(I745), .A2(W7500), .ZN(O7382));
  NANDX1 G22521 (.A1(W32462), .A2(W806), .ZN(O7380));
  NANDX1 G22522 (.A1(W10493), .A2(W13399), .ZN(O7378));
  NANDX1 G22523 (.A1(W14409), .A2(W2202), .ZN(W34657));
  NANDX1 G22524 (.A1(W25493), .A2(W30878), .ZN(W34653));
  NANDX1 G22525 (.A1(W90), .A2(W6393), .ZN(O7373));
  NANDX1 G22526 (.A1(W19065), .A2(W14944), .ZN(W34650));
  NANDX1 G22527 (.A1(W30255), .A2(W29090), .ZN(W34649));
  NANDX1 G22528 (.A1(W7155), .A2(W85), .ZN(O7282));
  NANDX1 G22529 (.A1(W32961), .A2(W3026), .ZN(O7302));
  NANDX1 G22530 (.A1(W14147), .A2(W7495), .ZN(O7298));
  NANDX1 G22531 (.A1(W6569), .A2(W23827), .ZN(W34501));
  NANDX1 G22532 (.A1(W20919), .A2(I423), .ZN(O7290));
  NANDX1 G22533 (.A1(W25878), .A2(W13822), .ZN(W34493));
  NANDX1 G22534 (.A1(W11713), .A2(W2766), .ZN(O7288));
  NANDX1 G22535 (.A1(W26864), .A2(W23924), .ZN(O7286));
  NANDX1 G22536 (.A1(W25316), .A2(W2126), .ZN(O7285));
  NANDX1 G22537 (.A1(W1840), .A2(W28821), .ZN(W34484));
  NANDX1 G22538 (.A1(W14927), .A2(W4600), .ZN(W34482));
  NANDX1 G22539 (.A1(W22836), .A2(W31855), .ZN(W34481));
  NANDX1 G22540 (.A1(W19793), .A2(W427), .ZN(W34479));
  NANDX1 G22541 (.A1(W26222), .A2(W1642), .ZN(O7304));
  NANDX1 G22542 (.A1(W20546), .A2(W7753), .ZN(O7280));
  NANDX1 G22543 (.A1(W21888), .A2(W17312), .ZN(O7278));
  NANDX1 G22544 (.A1(W31310), .A2(W13155), .ZN(O7277));
  NANDX1 G22545 (.A1(W28361), .A2(W25790), .ZN(W34471));
  NANDX1 G22546 (.A1(W13985), .A2(W23810), .ZN(O7274));
  NANDX1 G22547 (.A1(W15749), .A2(W32625), .ZN(W34466));
  NANDX1 G22548 (.A1(W4092), .A2(W2799), .ZN(O7272));
  NANDX1 G22549 (.A1(W22530), .A2(W5060), .ZN(O7270));
  NANDX1 G22550 (.A1(W31614), .A2(W11558), .ZN(O7268));
  NANDX1 G22551 (.A1(W7536), .A2(W6188), .ZN(W34457));
  NANDX1 G22552 (.A1(W13018), .A2(W4157), .ZN(O7266));
  NANDX1 G22553 (.A1(W793), .A2(W25891), .ZN(W34553));
  NANDX1 G22554 (.A1(W23940), .A2(W21951), .ZN(O7339));
  NANDX1 G22555 (.A1(W22828), .A2(W25243), .ZN(W34583));
  NANDX1 G22556 (.A1(W10584), .A2(W11853), .ZN(O7338));
  NANDX1 G22557 (.A1(W7300), .A2(W15980), .ZN(W34578));
  NANDX1 G22558 (.A1(W30355), .A2(W15394), .ZN(O7332));
  NANDX1 G22559 (.A1(W26284), .A2(W4093), .ZN(W34569));
  NANDX1 G22560 (.A1(W34528), .A2(W13189), .ZN(W34567));
  NANDX1 G22561 (.A1(W32374), .A2(W16088), .ZN(W34564));
  NANDX1 G22562 (.A1(W21012), .A2(W22284), .ZN(W34562));
  NANDX1 G22563 (.A1(W31779), .A2(W12488), .ZN(W34560));
  NANDX1 G22564 (.A1(W4525), .A2(W14317), .ZN(W34557));
  NANDX1 G22565 (.A1(W9263), .A2(I833), .ZN(W35330));
  NANDX1 G22566 (.A1(W8225), .A2(W31611), .ZN(O7324));
  NANDX1 G22567 (.A1(W13892), .A2(W3383), .ZN(W34549));
  NANDX1 G22568 (.A1(W32289), .A2(W30412), .ZN(O7322));
  NANDX1 G22569 (.A1(W6672), .A2(W29179), .ZN(W34543));
  NANDX1 G22570 (.A1(W22625), .A2(W26487), .ZN(W34540));
  NANDX1 G22571 (.A1(W20898), .A2(W18143), .ZN(O7314));
  NANDX1 G22572 (.A1(W15735), .A2(W6029), .ZN(W34534));
  NANDX1 G22573 (.A1(W20217), .A2(W3806), .ZN(O7312));
  NANDX1 G22574 (.A1(W1736), .A2(W16979), .ZN(W34526));
  NANDX1 G22575 (.A1(W1543), .A2(W7874), .ZN(W34524));
  NANDX1 G22576 (.A1(W30733), .A2(W21925), .ZN(O7305));
  NANDX1 G22577 (.A1(W14407), .A2(W13195), .ZN(O8179));
  NANDX1 G22578 (.A1(W7272), .A2(W7754), .ZN(O8194));
  NANDX1 G22579 (.A1(W16583), .A2(W3352), .ZN(O8192));
  NANDX1 G22580 (.A1(W28944), .A2(W26941), .ZN(O8189));
  NANDX1 G22581 (.A1(W7480), .A2(W19614), .ZN(O8188));
  NANDX1 G22582 (.A1(W34653), .A2(W22845), .ZN(W36079));
  NANDX1 G22583 (.A1(W30215), .A2(W22308), .ZN(O8187));
  NANDX1 G22584 (.A1(W17176), .A2(W5826), .ZN(W36073));
  NANDX1 G22585 (.A1(W14747), .A2(W4815), .ZN(W36070));
  NANDX1 G22586 (.A1(I1194), .A2(W6501), .ZN(O8182));
  NANDX1 G22587 (.A1(W32232), .A2(W10962), .ZN(W36067));
  NANDX1 G22588 (.A1(W32651), .A2(W23266), .ZN(W36065));
  NANDX1 G22589 (.A1(W5665), .A2(W27171), .ZN(O8180));
  NANDX1 G22590 (.A1(W12363), .A2(W28706), .ZN(W36092));
  NANDX1 G22591 (.A1(W31378), .A2(W11469), .ZN(W36061));
  NANDX1 G22592 (.A1(W1513), .A2(W22879), .ZN(O8176));
  NANDX1 G22593 (.A1(W33095), .A2(W29621), .ZN(O8170));
  NANDX1 G22594 (.A1(W2200), .A2(W30699), .ZN(O8169));
  NANDX1 G22595 (.A1(W29340), .A2(W7481), .ZN(O8168));
  NANDX1 G22596 (.A1(W21264), .A2(W12122), .ZN(O8167));
  NANDX1 G22597 (.A1(W9648), .A2(W22883), .ZN(W36047));
  NANDX1 G22598 (.A1(W20017), .A2(W8062), .ZN(O8166));
  NANDX1 G22599 (.A1(W370), .A2(I1585), .ZN(O8165));
  NANDX1 G22600 (.A1(W9154), .A2(W10160), .ZN(O8164));
  NANDX1 G22601 (.A1(W8747), .A2(W32809), .ZN(O8163));
  NANDX1 G22602 (.A1(W14096), .A2(W22437), .ZN(O8215));
  NANDX1 G22603 (.A1(W26173), .A2(W25277), .ZN(O8236));
  NANDX1 G22604 (.A1(W26490), .A2(W17850), .ZN(W36164));
  NANDX1 G22605 (.A1(W8686), .A2(W32636), .ZN(W36161));
  NANDX1 G22606 (.A1(W15507), .A2(W20512), .ZN(O8234));
  NANDX1 G22607 (.A1(W15074), .A2(W36111), .ZN(W36157));
  NANDX1 G22608 (.A1(W20590), .A2(W26614), .ZN(O8230));
  NANDX1 G22609 (.A1(W26834), .A2(W15782), .ZN(W36149));
  NANDX1 G22610 (.A1(W9947), .A2(W27102), .ZN(O8226));
  NANDX1 G22611 (.A1(W5280), .A2(W15631), .ZN(W36143));
  NANDX1 G22612 (.A1(I1626), .A2(W26083), .ZN(W36139));
  NANDX1 G22613 (.A1(W19986), .A2(W28972), .ZN(W36133));
  NANDX1 G22614 (.A1(W30844), .A2(W21613), .ZN(O8220));
  NANDX1 G22615 (.A1(I1040), .A2(W18481), .ZN(W36042));
  NANDX1 G22616 (.A1(W13576), .A2(W31827), .ZN(W36121));
  NANDX1 G22617 (.A1(W28438), .A2(W21834), .ZN(O8214));
  NANDX1 G22618 (.A1(W2934), .A2(W3333), .ZN(O8212));
  NANDX1 G22619 (.A1(W21991), .A2(W28367), .ZN(O8208));
  NANDX1 G22620 (.A1(W25575), .A2(W13171), .ZN(O8206));
  NANDX1 G22621 (.A1(W32878), .A2(W27434), .ZN(O8205));
  NANDX1 G22622 (.A1(W15614), .A2(W17017), .ZN(W36106));
  NANDX1 G22623 (.A1(W15594), .A2(W5021), .ZN(O8203));
  NANDX1 G22624 (.A1(W8518), .A2(W21835), .ZN(W36104));
  NANDX1 G22625 (.A1(W1638), .A2(W31368), .ZN(O8201));
  NANDX1 G22626 (.A1(W964), .A2(W33158), .ZN(O8199));
  NANDX1 G22627 (.A1(W31580), .A2(I1619), .ZN(W35929));
  NANDX1 G22628 (.A1(W9306), .A2(W18162), .ZN(O8112));
  NANDX1 G22629 (.A1(W5782), .A2(I521), .ZN(W35958));
  NANDX1 G22630 (.A1(W31388), .A2(W29316), .ZN(W35956));
  NANDX1 G22631 (.A1(W2788), .A2(W17532), .ZN(O8107));
  NANDX1 G22632 (.A1(W3195), .A2(W22109), .ZN(O8106));
  NANDX1 G22633 (.A1(W22508), .A2(W1031), .ZN(W35950));
  NANDX1 G22634 (.A1(W3212), .A2(W31354), .ZN(W35946));
  NANDX1 G22635 (.A1(W25862), .A2(W9516), .ZN(O8103));
  NANDX1 G22636 (.A1(W8726), .A2(W13756), .ZN(O8101));
  NANDX1 G22637 (.A1(W4789), .A2(W22696), .ZN(O8100));
  NANDX1 G22638 (.A1(W11226), .A2(W7737), .ZN(O8098));
  NANDX1 G22639 (.A1(W32074), .A2(W28762), .ZN(O8093));
  NANDX1 G22640 (.A1(W31100), .A2(W25987), .ZN(W35963));
  NANDX1 G22641 (.A1(W25110), .A2(W7659), .ZN(W35925));
  NANDX1 G22642 (.A1(W18898), .A2(W6543), .ZN(O8089));
  NANDX1 G22643 (.A1(W7978), .A2(W33644), .ZN(W35923));
  NANDX1 G22644 (.A1(W25925), .A2(W1874), .ZN(W35921));
  NANDX1 G22645 (.A1(W10172), .A2(W20784), .ZN(O8087));
  NANDX1 G22646 (.A1(W35672), .A2(W18473), .ZN(W35912));
  NANDX1 G22647 (.A1(W20635), .A2(W22026), .ZN(O8080));
  NANDX1 G22648 (.A1(W28399), .A2(W31160), .ZN(O8079));
  NANDX1 G22649 (.A1(W26572), .A2(W142), .ZN(O8078));
  NANDX1 G22650 (.A1(W14324), .A2(W29700), .ZN(O8076));
  NANDX1 G22651 (.A1(W32648), .A2(W16826), .ZN(W35903));
  NANDX1 G22652 (.A1(W7197), .A2(W21616), .ZN(W36004));
  NANDX1 G22653 (.A1(W22869), .A2(W24282), .ZN(W36040));
  NANDX1 G22654 (.A1(W421), .A2(W16461), .ZN(W36037));
  NANDX1 G22655 (.A1(W10424), .A2(W17308), .ZN(O8159));
  NANDX1 G22656 (.A1(W30135), .A2(W35556), .ZN(W36031));
  NANDX1 G22657 (.A1(W32568), .A2(W20112), .ZN(O8151));
  NANDX1 G22658 (.A1(W12886), .A2(W9327), .ZN(O8150));
  NANDX1 G22659 (.A1(W1837), .A2(W12263), .ZN(W36023));
  NANDX1 G22660 (.A1(W25961), .A2(W6471), .ZN(O8148));
  NANDX1 G22661 (.A1(W7079), .A2(W28231), .ZN(W36017));
  NANDX1 G22662 (.A1(W21588), .A2(W34084), .ZN(W36016));
  NANDX1 G22663 (.A1(W22035), .A2(W26998), .ZN(O8144));
  NANDX1 G22664 (.A1(W29644), .A2(W21178), .ZN(O8237));
  NANDX1 G22665 (.A1(W31784), .A2(W11219), .ZN(W36002));
  NANDX1 G22666 (.A1(W31754), .A2(W34917), .ZN(O8134));
  NANDX1 G22667 (.A1(W12309), .A2(W14614), .ZN(O8132));
  NANDX1 G22668 (.A1(W25728), .A2(W10160), .ZN(W35993));
  NANDX1 G22669 (.A1(W34145), .A2(W4882), .ZN(O8129));
  NANDX1 G22670 (.A1(W24296), .A2(W5554), .ZN(O8127));
  NANDX1 G22671 (.A1(W9093), .A2(W31170), .ZN(W35976));
  NANDX1 G22672 (.A1(W34667), .A2(W31241), .ZN(O8120));
  NANDX1 G22673 (.A1(W20366), .A2(W18473), .ZN(W35972));
  NANDX1 G22674 (.A1(W35215), .A2(W25042), .ZN(O8117));
  NANDX1 G22675 (.A1(W35776), .A2(W12731), .ZN(W35968));
  NANDX1 G22676 (.A1(W30488), .A2(W26247), .ZN(O8358));
  NANDX1 G22677 (.A1(W34305), .A2(W286), .ZN(W36403));
  NANDX1 G22678 (.A1(W22923), .A2(W20790), .ZN(W36399));
  NANDX1 G22679 (.A1(W3799), .A2(W25310), .ZN(O8374));
  NANDX1 G22680 (.A1(W13), .A2(W25205), .ZN(W36396));
  NANDX1 G22681 (.A1(W15351), .A2(W17597), .ZN(O8372));
  NANDX1 G22682 (.A1(W28646), .A2(W8616), .ZN(O8370));
  NANDX1 G22683 (.A1(W10200), .A2(W12216), .ZN(O8369));
  NANDX1 G22684 (.A1(W30893), .A2(W14082), .ZN(O8366));
  NANDX1 G22685 (.A1(W1353), .A2(W25786), .ZN(O8365));
  NANDX1 G22686 (.A1(W24085), .A2(W33457), .ZN(O8364));
  NANDX1 G22687 (.A1(W8106), .A2(W27179), .ZN(O8361));
  NANDX1 G22688 (.A1(W4453), .A2(W22346), .ZN(O8360));
  NANDX1 G22689 (.A1(W3660), .A2(W20955), .ZN(W36405));
  NANDX1 G22690 (.A1(W15666), .A2(W32467), .ZN(O8353));
  NANDX1 G22691 (.A1(W31494), .A2(W19116), .ZN(O8350));
  NANDX1 G22692 (.A1(W3206), .A2(W14045), .ZN(O8348));
  NANDX1 G22693 (.A1(W2350), .A2(W15711), .ZN(O8346));
  NANDX1 G22694 (.A1(W33406), .A2(W6411), .ZN(O8345));
  NANDX1 G22695 (.A1(W34679), .A2(W1671), .ZN(O8344));
  NANDX1 G22696 (.A1(W24393), .A2(W6134), .ZN(O8342));
  NANDX1 G22697 (.A1(W26871), .A2(W21022), .ZN(O8339));
  NANDX1 G22698 (.A1(W26515), .A2(W20863), .ZN(O8338));
  NANDX1 G22699 (.A1(W30615), .A2(W10806), .ZN(W36342));
  NANDX1 G22700 (.A1(W31836), .A2(W8502), .ZN(W36329));
  NANDX1 G22701 (.A1(W5994), .A2(W10028), .ZN(O8399));
  NANDX1 G22702 (.A1(W322), .A2(W21927), .ZN(O8426));
  NANDX1 G22703 (.A1(W32906), .A2(W4690), .ZN(O8425));
  NANDX1 G22704 (.A1(W8233), .A2(I215), .ZN(W36480));
  NANDX1 G22705 (.A1(W27074), .A2(W29849), .ZN(O8419));
  NANDX1 G22706 (.A1(W31783), .A2(W35326), .ZN(W36474));
  NANDX1 G22707 (.A1(W33656), .A2(W23839), .ZN(O8416));
  NANDX1 G22708 (.A1(W7932), .A2(W25040), .ZN(W36470));
  NANDX1 G22709 (.A1(W22107), .A2(W11541), .ZN(W36463));
  NANDX1 G22710 (.A1(I1141), .A2(W19836), .ZN(W36460));
  NANDX1 G22711 (.A1(W7665), .A2(W895), .ZN(O8408));
  NANDX1 G22712 (.A1(W13212), .A2(W30669), .ZN(W36456));
  NANDX1 G22713 (.A1(W8743), .A2(W5816), .ZN(W36453));
  NANDX1 G22714 (.A1(W34743), .A2(W5004), .ZN(W36327));
  NANDX1 G22715 (.A1(W30263), .A2(W2777), .ZN(O8395));
  NANDX1 G22716 (.A1(W4261), .A2(W10391), .ZN(O8394));
  NANDX1 G22717 (.A1(W3604), .A2(W14400), .ZN(W36433));
  NANDX1 G22718 (.A1(W5040), .A2(W6049), .ZN(O8393));
  NANDX1 G22719 (.A1(W28776), .A2(W8601), .ZN(O8387));
  NANDX1 G22720 (.A1(W1968), .A2(W18953), .ZN(W36418));
  NANDX1 G22721 (.A1(W23546), .A2(W16067), .ZN(W36413));
  NANDX1 G22722 (.A1(I1510), .A2(W1420), .ZN(W36411));
  NANDX1 G22723 (.A1(W18946), .A2(W5774), .ZN(O8380));
  NANDX1 G22724 (.A1(W13726), .A2(W23468), .ZN(O8379));
  NANDX1 G22725 (.A1(W24049), .A2(W1816), .ZN(O8378));
  NANDX1 G22726 (.A1(W29534), .A2(W17756), .ZN(O8254));
  NANDX1 G22727 (.A1(W17028), .A2(I1917), .ZN(W36252));
  NANDX1 G22728 (.A1(W19233), .A2(W8379), .ZN(W36248));
  NANDX1 G22729 (.A1(W13637), .A2(W16884), .ZN(W36247));
  NANDX1 G22730 (.A1(W11635), .A2(W20528), .ZN(W36240));
  NANDX1 G22731 (.A1(W22697), .A2(W2514), .ZN(O8276));
  NANDX1 G22732 (.A1(W17230), .A2(W13594), .ZN(W36235));
  NANDX1 G22733 (.A1(W29777), .A2(W11899), .ZN(O8272));
  NANDX1 G22734 (.A1(W4446), .A2(W34770), .ZN(W36226));
  NANDX1 G22735 (.A1(W29267), .A2(W3510), .ZN(O8260));
  NANDX1 G22736 (.A1(I1894), .A2(W12047), .ZN(W36211));
  NANDX1 G22737 (.A1(W2196), .A2(W12467), .ZN(W36210));
  NANDX1 G22738 (.A1(W33486), .A2(W8809), .ZN(W36201));
  NANDX1 G22739 (.A1(W24015), .A2(W29356), .ZN(W36255));
  NANDX1 G22740 (.A1(I564), .A2(W24289), .ZN(W36196));
  NANDX1 G22741 (.A1(W10374), .A2(W5779), .ZN(W36194));
  NANDX1 G22742 (.A1(W8218), .A2(W26287), .ZN(O8252));
  NANDX1 G22743 (.A1(W34620), .A2(W3360), .ZN(O8251));
  NANDX1 G22744 (.A1(W9590), .A2(I1634), .ZN(W36187));
  NANDX1 G22745 (.A1(W26732), .A2(W35074), .ZN(W36186));
  NANDX1 G22746 (.A1(W5938), .A2(W18629), .ZN(O8246));
  NANDX1 G22747 (.A1(W5384), .A2(W5796), .ZN(O8245));
  NANDX1 G22748 (.A1(W18151), .A2(W28950), .ZN(W36180));
  NANDX1 G22749 (.A1(W21713), .A2(W15974), .ZN(O8240));
  NANDX1 G22750 (.A1(W546), .A2(W28967), .ZN(O8239));
  NANDX1 G22751 (.A1(W18834), .A2(W3377), .ZN(W36294));
  NANDX1 G22752 (.A1(W12143), .A2(W10112), .ZN(O8327));
  NANDX1 G22753 (.A1(W9900), .A2(I826), .ZN(O8325));
  NANDX1 G22754 (.A1(W5765), .A2(W26485), .ZN(W36309));
  NANDX1 G22755 (.A1(W18483), .A2(W19964), .ZN(O8317));
  NANDX1 G22756 (.A1(W9015), .A2(W19157), .ZN(O8314));
  NANDX1 G22757 (.A1(W9462), .A2(I1026), .ZN(W36302));
  NANDX1 G22758 (.A1(W29988), .A2(W34752), .ZN(O8313));
  NANDX1 G22759 (.A1(W30598), .A2(W2019), .ZN(O8312));
  NANDX1 G22760 (.A1(W25987), .A2(W4293), .ZN(W36299));
  NANDX1 G22761 (.A1(W23061), .A2(W488), .ZN(O8311));
  NANDX1 G22762 (.A1(W5365), .A2(I1717), .ZN(O8310));
  NANDX1 G22763 (.A1(W33169), .A2(W5827), .ZN(O8074));
  NANDX1 G22764 (.A1(W9257), .A2(W21844), .ZN(O8306));
  NANDX1 G22765 (.A1(W11197), .A2(W30908), .ZN(O8302));
  NANDX1 G22766 (.A1(W17863), .A2(W29331), .ZN(O8301));
  NANDX1 G22767 (.A1(W29684), .A2(I337), .ZN(O8300));
  NANDX1 G22768 (.A1(W2772), .A2(W15325), .ZN(O8299));
  NANDX1 G22769 (.A1(W17745), .A2(W6151), .ZN(O8293));
  NANDX1 G22770 (.A1(W155), .A2(W8162), .ZN(O8292));
  NANDX1 G22771 (.A1(W9653), .A2(W30012), .ZN(W36267));
  NANDX1 G22772 (.A1(W20155), .A2(I1442), .ZN(W36264));
  NANDX1 G22773 (.A1(W8250), .A2(W19677), .ZN(O8288));
  NANDX1 G22774 (.A1(W13586), .A2(W4963), .ZN(O8284));
  NANDX1 G22775 (.A1(W26549), .A2(W5426), .ZN(W35534));
  NANDX1 G22776 (.A1(W22577), .A2(W1442), .ZN(W35565));
  NANDX1 G22777 (.A1(W1045), .A2(W19690), .ZN(W35564));
  NANDX1 G22778 (.A1(W871), .A2(W22931), .ZN(W35563));
  NANDX1 G22779 (.A1(W29603), .A2(W30559), .ZN(O7884));
  NANDX1 G22780 (.A1(W26282), .A2(W13579), .ZN(O7883));
  NANDX1 G22781 (.A1(W4459), .A2(I684), .ZN(O7878));
  NANDX1 G22782 (.A1(W7577), .A2(W20909), .ZN(O7876));
  NANDX1 G22783 (.A1(I1775), .A2(W12490), .ZN(O7875));
  NANDX1 G22784 (.A1(W557), .A2(W13113), .ZN(O7874));
  NANDX1 G22785 (.A1(W20848), .A2(W1079), .ZN(O7870));
  NANDX1 G22786 (.A1(W21584), .A2(W11839), .ZN(O7868));
  NANDX1 G22787 (.A1(W12905), .A2(W19260), .ZN(W35539));
  NANDX1 G22788 (.A1(W27978), .A2(W28611), .ZN(W35566));
  NANDX1 G22789 (.A1(W20884), .A2(W10331), .ZN(O7861));
  NANDX1 G22790 (.A1(I471), .A2(W9446), .ZN(W35529));
  NANDX1 G22791 (.A1(W6463), .A2(W21846), .ZN(O7856));
  NANDX1 G22792 (.A1(W5247), .A2(W12196), .ZN(O7855));
  NANDX1 G22793 (.A1(W15152), .A2(W23411), .ZN(O7853));
  NANDX1 G22794 (.A1(W13446), .A2(W8032), .ZN(O7851));
  NANDX1 G22795 (.A1(W26013), .A2(W517), .ZN(W35509));
  NANDX1 G22796 (.A1(W10541), .A2(W16800), .ZN(W35508));
  NANDX1 G22797 (.A1(W26256), .A2(W26829), .ZN(O7849));
  NANDX1 G22798 (.A1(W15536), .A2(W30847), .ZN(O7848));
  NANDX1 G22799 (.A1(W28505), .A2(W26103), .ZN(O7845));
  NANDX1 G22800 (.A1(W15128), .A2(W13886), .ZN(W35596));
  NANDX1 G22801 (.A1(W7354), .A2(W28013), .ZN(W35638));
  NANDX1 G22802 (.A1(W31353), .A2(I1393), .ZN(O7931));
  NANDX1 G22803 (.A1(W21919), .A2(W23939), .ZN(W35631));
  NANDX1 G22804 (.A1(W33743), .A2(W6519), .ZN(W35629));
  NANDX1 G22805 (.A1(W35431), .A2(W28368), .ZN(O7927));
  NANDX1 G22806 (.A1(W31847), .A2(W3873), .ZN(W35627));
  NANDX1 G22807 (.A1(W6964), .A2(W16337), .ZN(W35624));
  NANDX1 G22808 (.A1(W4896), .A2(W34217), .ZN(O7924));
  NANDX1 G22809 (.A1(W2673), .A2(W3240), .ZN(O7921));
  NANDX1 G22810 (.A1(W10529), .A2(W28523), .ZN(O7917));
  NANDX1 G22811 (.A1(W27792), .A2(W19783), .ZN(W35601));
  NANDX1 G22812 (.A1(W1199), .A2(W35409), .ZN(W35597));
  NANDX1 G22813 (.A1(W6052), .A2(W1621), .ZN(O7840));
  NANDX1 G22814 (.A1(W16075), .A2(W1575), .ZN(O7906));
  NANDX1 G22815 (.A1(W26174), .A2(W15359), .ZN(O7900));
  NANDX1 G22816 (.A1(W5588), .A2(W15755), .ZN(W35585));
  NANDX1 G22817 (.A1(W18750), .A2(W5529), .ZN(O7897));
  NANDX1 G22818 (.A1(W11597), .A2(I1674), .ZN(O7895));
  NANDX1 G22819 (.A1(W16123), .A2(W9956), .ZN(W35580));
  NANDX1 G22820 (.A1(W28444), .A2(W26550), .ZN(O7894));
  NANDX1 G22821 (.A1(W14189), .A2(W2606), .ZN(O7893));
  NANDX1 G22822 (.A1(W13855), .A2(W14499), .ZN(O7891));
  NANDX1 G22823 (.A1(W32581), .A2(I771), .ZN(O7890));
  NANDX1 G22824 (.A1(W31801), .A2(W17047), .ZN(O7885));
  NANDX1 G22825 (.A1(W18196), .A2(W2500), .ZN(W35359));
  NANDX1 G22826 (.A1(W34765), .A2(W13412), .ZN(O7782));
  NANDX1 G22827 (.A1(W29489), .A2(W35190), .ZN(O7781));
  NANDX1 G22828 (.A1(W5135), .A2(W20827), .ZN(O7776));
  NANDX1 G22829 (.A1(W15842), .A2(W11369), .ZN(W35391));
  NANDX1 G22830 (.A1(W25324), .A2(W7323), .ZN(O7774));
  NANDX1 G22831 (.A1(I1068), .A2(W12854), .ZN(W35388));
  NANDX1 G22832 (.A1(W14228), .A2(W4752), .ZN(W35386));
  NANDX1 G22833 (.A1(W25127), .A2(W13513), .ZN(W35373));
  NANDX1 G22834 (.A1(W24199), .A2(W18388), .ZN(O7766));
  NANDX1 G22835 (.A1(W29724), .A2(W18374), .ZN(O7763));
  NANDX1 G22836 (.A1(W12685), .A2(W30238), .ZN(W35362));
  NANDX1 G22837 (.A1(W19375), .A2(W6097), .ZN(O7760));
  NANDX1 G22838 (.A1(W8532), .A2(W4079), .ZN(O7790));
  NANDX1 G22839 (.A1(W26229), .A2(W21526), .ZN(O7759));
  NANDX1 G22840 (.A1(W19377), .A2(W33695), .ZN(W35354));
  NANDX1 G22841 (.A1(W17575), .A2(W22750), .ZN(W35348));
  NANDX1 G22842 (.A1(W17565), .A2(W20305), .ZN(O7753));
  NANDX1 G22843 (.A1(W30547), .A2(W11291), .ZN(O7752));
  NANDX1 G22844 (.A1(W21296), .A2(I108), .ZN(O7751));
  NANDX1 G22845 (.A1(W25347), .A2(W1276), .ZN(O7749));
  NANDX1 G22846 (.A1(W22807), .A2(W4952), .ZN(O7748));
  NANDX1 G22847 (.A1(W16771), .A2(W21764), .ZN(O7747));
  NANDX1 G22848 (.A1(W11532), .A2(W3808), .ZN(O7745));
  NANDX1 G22849 (.A1(W15113), .A2(W13619), .ZN(W35335));
  NANDX1 G22850 (.A1(W11504), .A2(W13541), .ZN(W35453));
  NANDX1 G22851 (.A1(W5341), .A2(W30933), .ZN(O7839));
  NANDX1 G22852 (.A1(W20854), .A2(W454), .ZN(O7833));
  NANDX1 G22853 (.A1(W954), .A2(W11888), .ZN(O7831));
  NANDX1 G22854 (.A1(W24323), .A2(W24760), .ZN(O7824));
  NANDX1 G22855 (.A1(W18522), .A2(W21352), .ZN(W35469));
  NANDX1 G22856 (.A1(W11177), .A2(W5752), .ZN(W35468));
  NANDX1 G22857 (.A1(W16337), .A2(W4064), .ZN(O7820));
  NANDX1 G22858 (.A1(W32815), .A2(W32690), .ZN(W35466));
  NANDX1 G22859 (.A1(W18020), .A2(W2855), .ZN(W35465));
  NANDX1 G22860 (.A1(W23552), .A2(W7356), .ZN(O7817));
  NANDX1 G22861 (.A1(W23290), .A2(W35395), .ZN(O7814));
  NANDX1 G22862 (.A1(W30804), .A2(W9488), .ZN(O7934));
  NANDX1 G22863 (.A1(W8109), .A2(W29202), .ZN(W35449));
  NANDX1 G22864 (.A1(W18062), .A2(W17771), .ZN(O7811));
  NANDX1 G22865 (.A1(W32975), .A2(W9661), .ZN(O7809));
  NANDX1 G22866 (.A1(W3291), .A2(W4115), .ZN(W35443));
  NANDX1 G22867 (.A1(W2314), .A2(W35144), .ZN(O7807));
  NANDX1 G22868 (.A1(W28444), .A2(W17832), .ZN(O7802));
  NANDX1 G22869 (.A1(W12829), .A2(W25010), .ZN(W35432));
  NANDX1 G22870 (.A1(W30572), .A2(W2841), .ZN(O7800));
  NANDX1 G22871 (.A1(W31932), .A2(W20876), .ZN(O7798));
  NANDX1 G22872 (.A1(W26324), .A2(W32437), .ZN(O7795));
  NANDX1 G22873 (.A1(W637), .A2(W33275), .ZN(O7794));
  NANDX1 G22874 (.A1(W4143), .A2(W12133), .ZN(W35803));
  NANDX1 G22875 (.A1(W27044), .A2(W34115), .ZN(O8031));
  NANDX1 G22876 (.A1(W20617), .A2(W10126), .ZN(W35824));
  NANDX1 G22877 (.A1(W21290), .A2(W7956), .ZN(W35823));
  NANDX1 G22878 (.A1(W19490), .A2(W24146), .ZN(W35822));
  NANDX1 G22879 (.A1(W12832), .A2(W557), .ZN(O8030));
  NANDX1 G22880 (.A1(W14872), .A2(W28501), .ZN(O8028));
  NANDX1 G22881 (.A1(W11112), .A2(W4659), .ZN(W35815));
  NANDX1 G22882 (.A1(W5826), .A2(W16249), .ZN(W35814));
  NANDX1 G22883 (.A1(W12656), .A2(W6033), .ZN(O8025));
  NANDX1 G22884 (.A1(W29523), .A2(W31630), .ZN(O8023));
  NANDX1 G22885 (.A1(W13597), .A2(W26170), .ZN(W35809));
  NANDX1 G22886 (.A1(W33086), .A2(W8610), .ZN(O8022));
  NANDX1 G22887 (.A1(W34191), .A2(W8391), .ZN(W35826));
  NANDX1 G22888 (.A1(W9202), .A2(W3918), .ZN(W35802));
  NANDX1 G22889 (.A1(W344), .A2(W540), .ZN(O8021));
  NANDX1 G22890 (.A1(W7217), .A2(W29550), .ZN(W35797));
  NANDX1 G22891 (.A1(W12074), .A2(W35547), .ZN(O8020));
  NANDX1 G22892 (.A1(W20254), .A2(W13826), .ZN(O8017));
  NANDX1 G22893 (.A1(W3136), .A2(I1100), .ZN(O8014));
  NANDX1 G22894 (.A1(W34037), .A2(I531), .ZN(O8012));
  NANDX1 G22895 (.A1(W16655), .A2(I1262), .ZN(O8010));
  NANDX1 G22896 (.A1(W28620), .A2(W17617), .ZN(W35781));
  NANDX1 G22897 (.A1(W15408), .A2(W8916), .ZN(W35771));
  NANDX1 G22898 (.A1(W28331), .A2(W34387), .ZN(O8004));
  NANDX1 G22899 (.A1(W32511), .A2(W7565), .ZN(O8050));
  NANDX1 G22900 (.A1(W4944), .A2(W10903), .ZN(O8068));
  NANDX1 G22901 (.A1(W7432), .A2(W12892), .ZN(W35893));
  NANDX1 G22902 (.A1(W25479), .A2(W26569), .ZN(O8064));
  NANDX1 G22903 (.A1(W26659), .A2(W12030), .ZN(O8059));
  NANDX1 G22904 (.A1(W10937), .A2(W12207), .ZN(O8058));
  NANDX1 G22905 (.A1(W32866), .A2(W30569), .ZN(W35875));
  NANDX1 G22906 (.A1(W29158), .A2(W16405), .ZN(W35869));
  NANDX1 G22907 (.A1(W3439), .A2(W7665), .ZN(O8054));
  NANDX1 G22908 (.A1(I320), .A2(W17280), .ZN(W35867));
  NANDX1 G22909 (.A1(W30374), .A2(W34649), .ZN(O8053));
  NANDX1 G22910 (.A1(W21903), .A2(W10196), .ZN(O8052));
  NANDX1 G22911 (.A1(W9031), .A2(W24523), .ZN(W35769));
  NANDX1 G22912 (.A1(W5271), .A2(W34105), .ZN(W35862));
  NANDX1 G22913 (.A1(W6264), .A2(W28777), .ZN(O8047));
  NANDX1 G22914 (.A1(W20953), .A2(W24383), .ZN(W35853));
  NANDX1 G22915 (.A1(W33841), .A2(W30170), .ZN(W35848));
  NANDX1 G22916 (.A1(W13978), .A2(W3453), .ZN(W35844));
  NANDX1 G22917 (.A1(W33469), .A2(W1748), .ZN(O8041));
  NANDX1 G22918 (.A1(W2788), .A2(W20274), .ZN(O8040));
  NANDX1 G22919 (.A1(W2069), .A2(W32463), .ZN(W35840));
  NANDX1 G22920 (.A1(W12808), .A2(W20770), .ZN(W35839));
  NANDX1 G22921 (.A1(W5056), .A2(W23021), .ZN(O8037));
  NANDX1 G22922 (.A1(W19489), .A2(W17768), .ZN(W35827));
  NANDX1 G22923 (.A1(W3530), .A2(W14852), .ZN(O7955));
  NANDX1 G22924 (.A1(W18462), .A2(W2189), .ZN(W35703));
  NANDX1 G22925 (.A1(W35634), .A2(W27017), .ZN(W35701));
  NANDX1 G22926 (.A1(W6498), .A2(W34376), .ZN(O7966));
  NANDX1 G22927 (.A1(W25582), .A2(W11361), .ZN(O7965));
  NANDX1 G22928 (.A1(W15887), .A2(W17523), .ZN(O7964));
  NANDX1 G22929 (.A1(W29279), .A2(W33754), .ZN(W35694));
  NANDX1 G22930 (.A1(W19183), .A2(W18140), .ZN(W35692));
  NANDX1 G22931 (.A1(W30289), .A2(W27473), .ZN(W35690));
  NANDX1 G22932 (.A1(W2975), .A2(W14015), .ZN(O7963));
  NANDX1 G22933 (.A1(W3111), .A2(W30960), .ZN(W35686));
  NANDX1 G22934 (.A1(W25368), .A2(W32316), .ZN(W35683));
  NANDX1 G22935 (.A1(W2916), .A2(W28525), .ZN(O7960));
  NANDX1 G22936 (.A1(W15393), .A2(W13701), .ZN(W35706));
  NANDX1 G22937 (.A1(W29498), .A2(W7309), .ZN(O7954));
  NANDX1 G22938 (.A1(W7930), .A2(W6942), .ZN(O7953));
  NANDX1 G22939 (.A1(W35565), .A2(W20540), .ZN(W35672));
  NANDX1 G22940 (.A1(W7884), .A2(W977), .ZN(W35670));
  NANDX1 G22941 (.A1(W31680), .A2(W15098), .ZN(O7950));
  NANDX1 G22942 (.A1(I1986), .A2(W11209), .ZN(W35664));
  NANDX1 G22943 (.A1(W20375), .A2(W12308), .ZN(W35655));
  NANDX1 G22944 (.A1(W7769), .A2(W14881), .ZN(O7944));
  NANDX1 G22945 (.A1(W33619), .A2(W3634), .ZN(O7938));
  NANDX1 G22946 (.A1(W10329), .A2(W23824), .ZN(W35646));
  NANDX1 G22947 (.A1(W25448), .A2(W11037), .ZN(W35645));
  NANDX1 G22948 (.A1(W10), .A2(W29721), .ZN(O7993));
  NANDX1 G22949 (.A1(W34809), .A2(W17140), .ZN(W35763));
  NANDX1 G22950 (.A1(W19533), .A2(W19606), .ZN(W35761));
  NANDX1 G22951 (.A1(W33583), .A2(W28294), .ZN(O8001));
  NANDX1 G22952 (.A1(W5487), .A2(W5357), .ZN(W35759));
  NANDX1 G22953 (.A1(W27757), .A2(W27943), .ZN(O8000));
  NANDX1 G22954 (.A1(W545), .A2(W18215), .ZN(O7999));
  NANDX1 G22955 (.A1(W4100), .A2(W3389), .ZN(W35755));
  NANDX1 G22956 (.A1(W2018), .A2(W24831), .ZN(W35754));
  NANDX1 G22957 (.A1(W27723), .A2(W21462), .ZN(W35751));
  NANDX1 G22958 (.A1(W26625), .A2(W813), .ZN(W35747));
  NANDX1 G22959 (.A1(W26209), .A2(W32467), .ZN(W35745));
  NANDX1 G22960 (.A1(W27594), .A2(W4255), .ZN(O7118));
  NANDX1 G22961 (.A1(W16983), .A2(W9832), .ZN(O7992));
  NANDX1 G22962 (.A1(W20310), .A2(W21772), .ZN(O7985));
  NANDX1 G22963 (.A1(W28125), .A2(W6873), .ZN(W35733));
  NANDX1 G22964 (.A1(W31874), .A2(W1582), .ZN(O7983));
  NANDX1 G22965 (.A1(W27101), .A2(W33284), .ZN(W35729));
  NANDX1 G22966 (.A1(W26742), .A2(W17353), .ZN(O7982));
  NANDX1 G22967 (.A1(W18866), .A2(W28291), .ZN(O7980));
  NANDX1 G22968 (.A1(W5092), .A2(W194), .ZN(W35719));
  NANDX1 G22969 (.A1(W31567), .A2(W9233), .ZN(O7974));
  NANDX1 G22970 (.A1(W11397), .A2(W10366), .ZN(O7973));
  NANDX1 G22971 (.A1(W7342), .A2(W2699), .ZN(W35710));
  NANDX1 G22972 (.A1(W18086), .A2(W5222), .ZN(W32637));
  NANDX1 G22973 (.A1(W19988), .A2(W31948), .ZN(W32667));
  NANDX1 G22974 (.A1(W3929), .A2(W24717), .ZN(W32665));
  NANDX1 G22975 (.A1(W9008), .A2(W19282), .ZN(O6335));
  NANDX1 G22976 (.A1(W1690), .A2(I68), .ZN(W32660));
  NANDX1 G22977 (.A1(W18499), .A2(I227), .ZN(W32656));
  NANDX1 G22978 (.A1(W12040), .A2(W28568), .ZN(W32653));
  NANDX1 G22979 (.A1(W16579), .A2(W1781), .ZN(O6331));
  NANDX1 G22980 (.A1(W22215), .A2(W12920), .ZN(W32648));
  NANDX1 G22981 (.A1(W22076), .A2(W2336), .ZN(O6330));
  NANDX1 G22982 (.A1(I1353), .A2(W21027), .ZN(O6329));
  NANDX1 G22983 (.A1(W17695), .A2(W28499), .ZN(W32641));
  NANDX1 G22984 (.A1(W19899), .A2(W5757), .ZN(W32640));
  NANDX1 G22985 (.A1(W21012), .A2(W3499), .ZN(W32669));
  NANDX1 G22986 (.A1(W8207), .A2(W21732), .ZN(W32635));
  NANDX1 G22987 (.A1(W22256), .A2(I1687), .ZN(W32633));
  NANDX1 G22988 (.A1(W20376), .A2(W17229), .ZN(O6321));
  NANDX1 G22989 (.A1(W32493), .A2(W20963), .ZN(O6320));
  NANDX1 G22990 (.A1(W28255), .A2(W1861), .ZN(O6318));
  NANDX1 G22991 (.A1(W25628), .A2(W7566), .ZN(W32621));
  NANDX1 G22992 (.A1(W29450), .A2(W31740), .ZN(W32618));
  NANDX1 G22993 (.A1(W15008), .A2(W32600), .ZN(W32617));
  NANDX1 G22994 (.A1(W23651), .A2(W24165), .ZN(W32616));
  NANDX1 G22995 (.A1(W7252), .A2(W25831), .ZN(O6314));
  NANDX1 G22996 (.A1(W646), .A2(W26625), .ZN(O6312));
  NANDX1 G22997 (.A1(W17280), .A2(W21259), .ZN(W32719));
  NANDX1 G22998 (.A1(W12312), .A2(W25558), .ZN(W32769));
  NANDX1 G22999 (.A1(W2738), .A2(I1985), .ZN(W32768));
  NANDX1 G23000 (.A1(W6032), .A2(W9042), .ZN(O6388));
  NANDX1 G23001 (.A1(W12308), .A2(W22866), .ZN(O6386));
  NANDX1 G23002 (.A1(W1224), .A2(W6058), .ZN(W32753));
  NANDX1 G23003 (.A1(W27390), .A2(W13695), .ZN(O6373));
  NANDX1 G23004 (.A1(W5256), .A2(W18938), .ZN(W32731));
  NANDX1 G23005 (.A1(W20434), .A2(I1478), .ZN(O6370));
  NANDX1 G23006 (.A1(W10108), .A2(W15636), .ZN(O6369));
  NANDX1 G23007 (.A1(W21101), .A2(W19424), .ZN(W32725));
  NANDX1 G23008 (.A1(W24989), .A2(W12993), .ZN(W32722));
  NANDX1 G23009 (.A1(W26178), .A2(W21919), .ZN(W32720));
  NANDX1 G23010 (.A1(W15814), .A2(W2371), .ZN(O6311));
  NANDX1 G23011 (.A1(W10260), .A2(W27945), .ZN(O6365));
  NANDX1 G23012 (.A1(W28209), .A2(W23082), .ZN(O6364));
  NANDX1 G23013 (.A1(W3384), .A2(W9019), .ZN(O6363));
  NANDX1 G23014 (.A1(W14351), .A2(W27895), .ZN(W32708));
  NANDX1 G23015 (.A1(W24202), .A2(W20185), .ZN(O6357));
  NANDX1 G23016 (.A1(W1161), .A2(W2430), .ZN(O6354));
  NANDX1 G23017 (.A1(W15621), .A2(W9530), .ZN(W32695));
  NANDX1 G23018 (.A1(W27723), .A2(W22748), .ZN(W32694));
  NANDX1 G23019 (.A1(W19477), .A2(W28666), .ZN(W32689));
  NANDX1 G23020 (.A1(W27820), .A2(W31163), .ZN(W32688));
  NANDX1 G23021 (.A1(W15436), .A2(W12374), .ZN(O6343));
  NANDX1 G23022 (.A1(W4393), .A2(W8127), .ZN(O6254));
  NANDX1 G23023 (.A1(W7165), .A2(W6227), .ZN(W32530));
  NANDX1 G23024 (.A1(W13526), .A2(W4797), .ZN(O6270));
  NANDX1 G23025 (.A1(W19265), .A2(W29544), .ZN(O6267));
  NANDX1 G23026 (.A1(W18979), .A2(W14325), .ZN(O6265));
  NANDX1 G23027 (.A1(W9755), .A2(W5831), .ZN(O6264));
  NANDX1 G23028 (.A1(W10679), .A2(W22217), .ZN(O6262));
  NANDX1 G23029 (.A1(I188), .A2(W6491), .ZN(W32512));
  NANDX1 G23030 (.A1(W6594), .A2(W1005), .ZN(O6261));
  NANDX1 G23031 (.A1(W31382), .A2(W26261), .ZN(O6259));
  NANDX1 G23032 (.A1(W31584), .A2(W5130), .ZN(O6258));
  NANDX1 G23033 (.A1(W12054), .A2(I1772), .ZN(O6257));
  NANDX1 G23034 (.A1(W21), .A2(W10603), .ZN(W32495));
  NANDX1 G23035 (.A1(W15), .A2(W19568), .ZN(W32532));
  NANDX1 G23036 (.A1(W23193), .A2(W25410), .ZN(O6253));
  NANDX1 G23037 (.A1(W24815), .A2(W20889), .ZN(O6250));
  NANDX1 G23038 (.A1(W22451), .A2(W4379), .ZN(W32480));
  NANDX1 G23039 (.A1(I1526), .A2(W768), .ZN(W32479));
  NANDX1 G23040 (.A1(W24842), .A2(W7155), .ZN(O6249));
  NANDX1 G23041 (.A1(W18662), .A2(W21287), .ZN(W32473));
  NANDX1 G23042 (.A1(W10084), .A2(W28339), .ZN(W32463));
  NANDX1 G23043 (.A1(W26384), .A2(W25082), .ZN(W32461));
  NANDX1 G23044 (.A1(W5957), .A2(W2681), .ZN(W32458));
  NANDX1 G23045 (.A1(W26101), .A2(W15969), .ZN(O6243));
  NANDX1 G23046 (.A1(W15445), .A2(W8939), .ZN(W32455));
  NANDX1 G23047 (.A1(W30853), .A2(W8403), .ZN(O6292));
  NANDX1 G23048 (.A1(W7590), .A2(W32578), .ZN(W32604));
  NANDX1 G23049 (.A1(W9314), .A2(W24168), .ZN(W32599));
  NANDX1 G23050 (.A1(W18607), .A2(W5224), .ZN(W32595));
  NANDX1 G23051 (.A1(W17253), .A2(W9253), .ZN(W32585));
  NANDX1 G23052 (.A1(W4452), .A2(W11356), .ZN(W32575));
  NANDX1 G23053 (.A1(W5382), .A2(W4152), .ZN(O6296));
  NANDX1 G23054 (.A1(W1553), .A2(W27725), .ZN(W32570));
  NANDX1 G23055 (.A1(W4270), .A2(W9737), .ZN(W32568));
  NANDX1 G23056 (.A1(W5489), .A2(W592), .ZN(O6293));
  NANDX1 G23057 (.A1(I1847), .A2(W1886), .ZN(W32566));
  NANDX1 G23058 (.A1(W5547), .A2(W22192), .ZN(W32565));
  NANDX1 G23059 (.A1(W4690), .A2(W541), .ZN(W32772));
  NANDX1 G23060 (.A1(W9425), .A2(W13490), .ZN(O6288));
  NANDX1 G23061 (.A1(W19048), .A2(W18289), .ZN(O6286));
  NANDX1 G23062 (.A1(W9874), .A2(W118), .ZN(O6284));
  NANDX1 G23063 (.A1(W22789), .A2(W11250), .ZN(O6283));
  NANDX1 G23064 (.A1(W20840), .A2(W17850), .ZN(O6278));
  NANDX1 G23065 (.A1(W28315), .A2(W10250), .ZN(O6277));
  NANDX1 G23066 (.A1(W23292), .A2(W31674), .ZN(O6276));
  NANDX1 G23067 (.A1(W13605), .A2(W24969), .ZN(O6275));
  NANDX1 G23068 (.A1(W7338), .A2(W12322), .ZN(O6273));
  NANDX1 G23069 (.A1(W10840), .A2(W20396), .ZN(O6272));
  NANDX1 G23070 (.A1(W19034), .A2(I812), .ZN(W32533));
  NANDX1 G23071 (.A1(W28467), .A2(I260), .ZN(O6464));
  NANDX1 G23072 (.A1(W7688), .A2(W16227), .ZN(W32976));
  NANDX1 G23073 (.A1(W10735), .A2(W8248), .ZN(O6482));
  NANDX1 G23074 (.A1(W28298), .A2(W13879), .ZN(W32972));
  NANDX1 G23075 (.A1(W31291), .A2(W30701), .ZN(O6480));
  NANDX1 G23076 (.A1(W8984), .A2(W7052), .ZN(W32970));
  NANDX1 G23077 (.A1(W26898), .A2(W28827), .ZN(W32961));
  NANDX1 G23078 (.A1(W262), .A2(W353), .ZN(O6474));
  NANDX1 G23079 (.A1(W29241), .A2(W16818), .ZN(W32949));
  NANDX1 G23080 (.A1(W18083), .A2(W30477), .ZN(W32947));
  NANDX1 G23081 (.A1(W12096), .A2(W32238), .ZN(O6467));
  NANDX1 G23082 (.A1(W22850), .A2(W24994), .ZN(W32943));
  NANDX1 G23083 (.A1(W15961), .A2(W22682), .ZN(W32942));
  NANDX1 G23084 (.A1(W15583), .A2(W29952), .ZN(O6483));
  NANDX1 G23085 (.A1(W18789), .A2(W25204), .ZN(O6463));
  NANDX1 G23086 (.A1(W6252), .A2(W29194), .ZN(W32933));
  NANDX1 G23087 (.A1(W22938), .A2(W6879), .ZN(O6461));
  NANDX1 G23088 (.A1(W13414), .A2(W8907), .ZN(W32923));
  NANDX1 G23089 (.A1(W17024), .A2(W22165), .ZN(W32909));
  NANDX1 G23090 (.A1(W25455), .A2(W17476), .ZN(W32907));
  NANDX1 G23091 (.A1(W8719), .A2(W1356), .ZN(O6452));
  NANDX1 G23092 (.A1(W12042), .A2(W24032), .ZN(W32904));
  NANDX1 G23093 (.A1(W3428), .A2(W32458), .ZN(W32903));
  NANDX1 G23094 (.A1(W20631), .A2(W1245), .ZN(W32902));
  NANDX1 G23095 (.A1(W24306), .A2(W9144), .ZN(W32899));
  NANDX1 G23096 (.A1(W604), .A2(W4758), .ZN(O6501));
  NANDX1 G23097 (.A1(W7903), .A2(W7477), .ZN(O6518));
  NANDX1 G23098 (.A1(I1166), .A2(W25462), .ZN(O6515));
  NANDX1 G23099 (.A1(W27539), .A2(W6678), .ZN(W33038));
  NANDX1 G23100 (.A1(W24292), .A2(W4688), .ZN(O6514));
  NANDX1 G23101 (.A1(W30249), .A2(W18342), .ZN(W33036));
  NANDX1 G23102 (.A1(W8478), .A2(W4343), .ZN(W33030));
  NANDX1 G23103 (.A1(W19951), .A2(W12630), .ZN(O6511));
  NANDX1 G23104 (.A1(W19869), .A2(W5511), .ZN(O6509));
  NANDX1 G23105 (.A1(W19131), .A2(W16461), .ZN(O6507));
  NANDX1 G23106 (.A1(W27038), .A2(W31439), .ZN(W33018));
  NANDX1 G23107 (.A1(W15589), .A2(W2744), .ZN(W33016));
  NANDX1 G23108 (.A1(W8631), .A2(W22358), .ZN(O6504));
  NANDX1 G23109 (.A1(W9215), .A2(W21572), .ZN(O6451));
  NANDX1 G23110 (.A1(W31728), .A2(W13236), .ZN(W33005));
  NANDX1 G23111 (.A1(W32715), .A2(W26267), .ZN(O6500));
  NANDX1 G23112 (.A1(W28973), .A2(I684), .ZN(O6499));
  NANDX1 G23113 (.A1(W4700), .A2(W27947), .ZN(W32997));
  NANDX1 G23114 (.A1(W20395), .A2(I1195), .ZN(O6494));
  NANDX1 G23115 (.A1(W2802), .A2(W8750), .ZN(W32992));
  NANDX1 G23116 (.A1(W8298), .A2(W4081), .ZN(O6492));
  NANDX1 G23117 (.A1(W17086), .A2(W20606), .ZN(O6489));
  NANDX1 G23118 (.A1(W4783), .A2(W32115), .ZN(O6487));
  NANDX1 G23119 (.A1(W15863), .A2(W21898), .ZN(O6486));
  NANDX1 G23120 (.A1(W17810), .A2(W25540), .ZN(O6484));
  NANDX1 G23121 (.A1(W20861), .A2(W16302), .ZN(O6402));
  NANDX1 G23122 (.A1(W6693), .A2(W15616), .ZN(O6425));
  NANDX1 G23123 (.A1(W23363), .A2(W29082), .ZN(W32837));
  NANDX1 G23124 (.A1(I1882), .A2(W23006), .ZN(O6419));
  NANDX1 G23125 (.A1(W6442), .A2(W9350), .ZN(O6418));
  NANDX1 G23126 (.A1(W9157), .A2(W20333), .ZN(W32824));
  NANDX1 G23127 (.A1(W16988), .A2(W19997), .ZN(W32819));
  NANDX1 G23128 (.A1(W25371), .A2(W12220), .ZN(W32815));
  NANDX1 G23129 (.A1(W1757), .A2(W11696), .ZN(O6408));
  NANDX1 G23130 (.A1(W14981), .A2(W15170), .ZN(O6407));
  NANDX1 G23131 (.A1(W1006), .A2(W11446), .ZN(W32810));
  NANDX1 G23132 (.A1(W21108), .A2(W10590), .ZN(W32808));
  NANDX1 G23133 (.A1(W10584), .A2(W24415), .ZN(W32806));
  NANDX1 G23134 (.A1(W8628), .A2(W6220), .ZN(W32842));
  NANDX1 G23135 (.A1(W25687), .A2(W24024), .ZN(O6400));
  NANDX1 G23136 (.A1(W7147), .A2(W19001), .ZN(W32794));
  NANDX1 G23137 (.A1(W20818), .A2(W24772), .ZN(W32789));
  NANDX1 G23138 (.A1(W1318), .A2(W17157), .ZN(W32784));
  NANDX1 G23139 (.A1(W22206), .A2(W24906), .ZN(W32783));
  NANDX1 G23140 (.A1(W12073), .A2(W9727), .ZN(W32781));
  NANDX1 G23141 (.A1(W27070), .A2(W32570), .ZN(W32780));
  NANDX1 G23142 (.A1(W6984), .A2(W2994), .ZN(W32779));
  NANDX1 G23143 (.A1(W1580), .A2(W1520), .ZN(O6391));
  NANDX1 G23144 (.A1(W22822), .A2(W7502), .ZN(W32774));
  NANDX1 G23145 (.A1(I1385), .A2(W20466), .ZN(O6390));
  NANDX1 G23146 (.A1(W32227), .A2(W8535), .ZN(O6440));
  NANDX1 G23147 (.A1(W5853), .A2(W29024), .ZN(W32897));
  NANDX1 G23148 (.A1(W4059), .A2(W811), .ZN(O6449));
  NANDX1 G23149 (.A1(W10343), .A2(W8111), .ZN(O6447));
  NANDX1 G23150 (.A1(W9817), .A2(W2849), .ZN(W32889));
  NANDX1 G23151 (.A1(W4927), .A2(W4335), .ZN(W32888));
  NANDX1 G23152 (.A1(W21782), .A2(W19148), .ZN(O6446));
  NANDX1 G23153 (.A1(W27615), .A2(W16823), .ZN(W32885));
  NANDX1 G23154 (.A1(W14256), .A2(W31576), .ZN(W32883));
  NANDX1 G23155 (.A1(W8040), .A2(W9509), .ZN(W32878));
  NANDX1 G23156 (.A1(W9846), .A2(W15624), .ZN(O6443));
  NANDX1 G23157 (.A1(W14034), .A2(W23972), .ZN(W32875));
  NANDX1 G23158 (.A1(W14584), .A2(W27916), .ZN(W32453));
  NANDX1 G23159 (.A1(W15592), .A2(W3476), .ZN(O6439));
  NANDX1 G23160 (.A1(W19460), .A2(W3656), .ZN(O6438));
  NANDX1 G23161 (.A1(I834), .A2(W21061), .ZN(O6437));
  NANDX1 G23162 (.A1(W23937), .A2(W30004), .ZN(W32864));
  NANDX1 G23163 (.A1(W17020), .A2(W24699), .ZN(W32863));
  NANDX1 G23164 (.A1(W2549), .A2(W28270), .ZN(W32862));
  NANDX1 G23165 (.A1(W30196), .A2(W22990), .ZN(W32861));
  NANDX1 G23166 (.A1(W2826), .A2(W8970), .ZN(W32859));
  NANDX1 G23167 (.A1(W6340), .A2(W9844), .ZN(W32854));
  NANDX1 G23168 (.A1(W3450), .A2(W27719), .ZN(O6430));
  NANDX1 G23169 (.A1(W11491), .A2(W17143), .ZN(O6428));
  NANDX1 G23170 (.A1(W25428), .A2(W14719), .ZN(O6077));
  NANDX1 G23171 (.A1(W1008), .A2(W7399), .ZN(O6090));
  NANDX1 G23172 (.A1(W15075), .A2(W27717), .ZN(W32097));
  NANDX1 G23173 (.A1(W18203), .A2(W5898), .ZN(O6089));
  NANDX1 G23174 (.A1(W5228), .A2(W21085), .ZN(O6087));
  NANDX1 G23175 (.A1(W20041), .A2(W22532), .ZN(W32087));
  NANDX1 G23176 (.A1(W24110), .A2(W29966), .ZN(O6085));
  NANDX1 G23177 (.A1(W19552), .A2(W26002), .ZN(O6084));
  NANDX1 G23178 (.A1(W21268), .A2(W16617), .ZN(O6083));
  NANDX1 G23179 (.A1(W24780), .A2(W3082), .ZN(W32077));
  NANDX1 G23180 (.A1(W28389), .A2(W27556), .ZN(W32075));
  NANDX1 G23181 (.A1(W4006), .A2(W14627), .ZN(W32071));
  NANDX1 G23182 (.A1(W26903), .A2(W17703), .ZN(W32069));
  NANDX1 G23183 (.A1(W17194), .A2(W11316), .ZN(W32101));
  NANDX1 G23184 (.A1(W8884), .A2(W20919), .ZN(W32066));
  NANDX1 G23185 (.A1(W6482), .A2(W4147), .ZN(O6072));
  NANDX1 G23186 (.A1(W4190), .A2(W22941), .ZN(W32053));
  NANDX1 G23187 (.A1(W10345), .A2(W12450), .ZN(W32052));
  NANDX1 G23188 (.A1(W24097), .A2(W15866), .ZN(O6070));
  NANDX1 G23189 (.A1(W30740), .A2(W1225), .ZN(O6068));
  NANDX1 G23190 (.A1(W24308), .A2(W27818), .ZN(W32040));
  NANDX1 G23191 (.A1(I1878), .A2(W30137), .ZN(W32036));
  NANDX1 G23192 (.A1(W4470), .A2(W30533), .ZN(O6063));
  NANDX1 G23193 (.A1(W29495), .A2(W8732), .ZN(W32028));
  NANDX1 G23194 (.A1(W14634), .A2(W24458), .ZN(O6061));
  NANDX1 G23195 (.A1(W20676), .A2(W26695), .ZN(O6105));
  NANDX1 G23196 (.A1(W11489), .A2(W14434), .ZN(O6135));
  NANDX1 G23197 (.A1(W31941), .A2(W24315), .ZN(O6134));
  NANDX1 G23198 (.A1(W16689), .A2(W32100), .ZN(W32177));
  NANDX1 G23199 (.A1(W7387), .A2(W23452), .ZN(O6131));
  NANDX1 G23200 (.A1(W16567), .A2(W7147), .ZN(O6130));
  NANDX1 G23201 (.A1(I220), .A2(W29010), .ZN(O6127));
  NANDX1 G23202 (.A1(W29405), .A2(W26292), .ZN(W32164));
  NANDX1 G23203 (.A1(W27318), .A2(W20618), .ZN(O6124));
  NANDX1 G23204 (.A1(W11298), .A2(W1467), .ZN(O6122));
  NANDX1 G23205 (.A1(W27203), .A2(W24098), .ZN(O6117));
  NANDX1 G23206 (.A1(W3781), .A2(W21615), .ZN(O6113));
  NANDX1 G23207 (.A1(W9666), .A2(W27072), .ZN(O6106));
  NANDX1 G23208 (.A1(W13629), .A2(W16833), .ZN(O6060));
  NANDX1 G23209 (.A1(I825), .A2(W13717), .ZN(W32131));
  NANDX1 G23210 (.A1(W26616), .A2(W19573), .ZN(O6103));
  NANDX1 G23211 (.A1(W13162), .A2(I1458), .ZN(O6099));
  NANDX1 G23212 (.A1(W31430), .A2(W31090), .ZN(O6098));
  NANDX1 G23213 (.A1(W6408), .A2(W16639), .ZN(W32114));
  NANDX1 G23214 (.A1(I1953), .A2(W16252), .ZN(O6095));
  NANDX1 G23215 (.A1(W15772), .A2(W13922), .ZN(W32109));
  NANDX1 G23216 (.A1(W4648), .A2(W14276), .ZN(O6093));
  NANDX1 G23217 (.A1(W17442), .A2(W16401), .ZN(W32106));
  NANDX1 G23218 (.A1(W3812), .A2(W10492), .ZN(W32104));
  NANDX1 G23219 (.A1(W29359), .A2(W3708), .ZN(O6091));
  NANDX1 G23220 (.A1(W9183), .A2(W6923), .ZN(O6002));
  NANDX1 G23221 (.A1(W10045), .A2(W28266), .ZN(O6014));
  NANDX1 G23222 (.A1(W22151), .A2(W3697), .ZN(W31927));
  NANDX1 G23223 (.A1(W7837), .A2(W28902), .ZN(W31925));
  NANDX1 G23224 (.A1(W11973), .A2(W16400), .ZN(W31917));
  NANDX1 G23225 (.A1(W30112), .A2(W10382), .ZN(W31914));
  NANDX1 G23226 (.A1(W5833), .A2(W401), .ZN(W31912));
  NANDX1 G23227 (.A1(W14524), .A2(W30619), .ZN(W31910));
  NANDX1 G23228 (.A1(W672), .A2(W4737), .ZN(O6007));
  NANDX1 G23229 (.A1(W127), .A2(W27083), .ZN(O6006));
  NANDX1 G23230 (.A1(W17572), .A2(W5650), .ZN(W31901));
  NANDX1 G23231 (.A1(W5901), .A2(W15956), .ZN(O6003));
  NANDX1 G23232 (.A1(W218), .A2(W8181), .ZN(W31899));
  NANDX1 G23233 (.A1(I626), .A2(W30364), .ZN(W31934));
  NANDX1 G23234 (.A1(W12695), .A2(W28849), .ZN(W31881));
  NANDX1 G23235 (.A1(W27206), .A2(W1753), .ZN(O5992));
  NANDX1 G23236 (.A1(W16250), .A2(W21707), .ZN(W31872));
  NANDX1 G23237 (.A1(W26914), .A2(W7387), .ZN(O5984));
  NANDX1 G23238 (.A1(W15954), .A2(W10935), .ZN(O5978));
  NANDX1 G23239 (.A1(W11966), .A2(W22365), .ZN(W31855));
  NANDX1 G23240 (.A1(W30307), .A2(W1975), .ZN(O5976));
  NANDX1 G23241 (.A1(W23957), .A2(W14765), .ZN(O5975));
  NANDX1 G23242 (.A1(W30868), .A2(W16380), .ZN(W31842));
  NANDX1 G23243 (.A1(W30384), .A2(W2950), .ZN(O5971));
  NANDX1 G23244 (.A1(W29953), .A2(W21473), .ZN(W31834));
  NANDX1 G23245 (.A1(W22764), .A2(W2901), .ZN(W31984));
  NANDX1 G23246 (.A1(I744), .A2(W30116), .ZN(O6059));
  NANDX1 G23247 (.A1(W15153), .A2(W20649), .ZN(O6055));
  NANDX1 G23248 (.A1(W27643), .A2(W19012), .ZN(W32015));
  NANDX1 G23249 (.A1(W16339), .A2(W15358), .ZN(O6053));
  NANDX1 G23250 (.A1(I1747), .A2(W13854), .ZN(O6048));
  NANDX1 G23251 (.A1(W19645), .A2(W23611), .ZN(O6047));
  NANDX1 G23252 (.A1(W895), .A2(W3447), .ZN(O6043));
  NANDX1 G23253 (.A1(W722), .A2(W26012), .ZN(W31995));
  NANDX1 G23254 (.A1(W19294), .A2(W11911), .ZN(O6040));
  NANDX1 G23255 (.A1(W20412), .A2(W28074), .ZN(O6039));
  NANDX1 G23256 (.A1(W7001), .A2(W2831), .ZN(W31987));
  NANDX1 G23257 (.A1(W14960), .A2(W28268), .ZN(W32188));
  NANDX1 G23258 (.A1(W18219), .A2(W3945), .ZN(W31982));
  NANDX1 G23259 (.A1(W26415), .A2(W25241), .ZN(W31981));
  NANDX1 G23260 (.A1(W16273), .A2(W30930), .ZN(W31978));
  NANDX1 G23261 (.A1(W20901), .A2(W5821), .ZN(W31976));
  NANDX1 G23262 (.A1(W14444), .A2(W11245), .ZN(O6028));
  NANDX1 G23263 (.A1(W5338), .A2(W7206), .ZN(W31963));
  NANDX1 G23264 (.A1(W18678), .A2(W7726), .ZN(W31959));
  NANDX1 G23265 (.A1(W18166), .A2(W9259), .ZN(O6022));
  NANDX1 G23266 (.A1(W10), .A2(W29929), .ZN(O6021));
  NANDX1 G23267 (.A1(W26339), .A2(W28883), .ZN(W31938));
  NANDX1 G23268 (.A1(W5445), .A2(W3117), .ZN(O6016));
  NANDX1 G23269 (.A1(W17416), .A2(W30899), .ZN(O6204));
  NANDX1 G23270 (.A1(W7366), .A2(W32052), .ZN(W32390));
  NANDX1 G23271 (.A1(W30765), .A2(W15163), .ZN(W32386));
  NANDX1 G23272 (.A1(W5884), .A2(W5619), .ZN(W32383));
  NANDX1 G23273 (.A1(W28586), .A2(W20233), .ZN(O6215));
  NANDX1 G23274 (.A1(W10760), .A2(W13770), .ZN(W32379));
  NANDX1 G23275 (.A1(W4801), .A2(W29559), .ZN(O6214));
  NANDX1 G23276 (.A1(W16593), .A2(W24726), .ZN(O6212));
  NANDX1 G23277 (.A1(W15976), .A2(W4566), .ZN(W32374));
  NANDX1 G23278 (.A1(W1223), .A2(W3340), .ZN(W32367));
  NANDX1 G23279 (.A1(I498), .A2(W12710), .ZN(W32364));
  NANDX1 G23280 (.A1(W26640), .A2(W4777), .ZN(W32363));
  NANDX1 G23281 (.A1(W12446), .A2(W25661), .ZN(O6205));
  NANDX1 G23282 (.A1(W17380), .A2(W27247), .ZN(W32397));
  NANDX1 G23283 (.A1(W27096), .A2(W3532), .ZN(W32351));
  NANDX1 G23284 (.A1(W22264), .A2(W30084), .ZN(W32347));
  NANDX1 G23285 (.A1(W20889), .A2(W24401), .ZN(W32344));
  NANDX1 G23286 (.A1(W5646), .A2(W16910), .ZN(W32343));
  NANDX1 G23287 (.A1(W29387), .A2(W21087), .ZN(O6200));
  NANDX1 G23288 (.A1(W22788), .A2(W9777), .ZN(O6197));
  NANDX1 G23289 (.A1(W19704), .A2(W30427), .ZN(O6196));
  NANDX1 G23290 (.A1(W7070), .A2(W1506), .ZN(W32334));
  NANDX1 G23291 (.A1(W27388), .A2(W6263), .ZN(O6195));
  NANDX1 G23292 (.A1(W27854), .A2(I1014), .ZN(O6194));
  NANDX1 G23293 (.A1(W27549), .A2(W16273), .ZN(W32330));
  NANDX1 G23294 (.A1(W18463), .A2(W21406), .ZN(W32423));
  NANDX1 G23295 (.A1(W11144), .A2(W23879), .ZN(W32448));
  NANDX1 G23296 (.A1(W18222), .A2(W20879), .ZN(O6240));
  NANDX1 G23297 (.A1(W32294), .A2(W29806), .ZN(W32443));
  NANDX1 G23298 (.A1(W22003), .A2(W6641), .ZN(O6239));
  NANDX1 G23299 (.A1(W30591), .A2(W3205), .ZN(W32440));
  NANDX1 G23300 (.A1(W32406), .A2(W3652), .ZN(W32436));
  NANDX1 G23301 (.A1(W4423), .A2(W13322), .ZN(W32434));
  NANDX1 G23302 (.A1(W18144), .A2(W4038), .ZN(O6235));
  NANDX1 G23303 (.A1(W24209), .A2(W21870), .ZN(W32426));
  NANDX1 G23304 (.A1(W29236), .A2(W20625), .ZN(W32425));
  NANDX1 G23305 (.A1(W20029), .A2(W31454), .ZN(W32424));
  NANDX1 G23306 (.A1(I815), .A2(W16582), .ZN(W32324));
  NANDX1 G23307 (.A1(W18954), .A2(I1277), .ZN(W32422));
  NANDX1 G23308 (.A1(W21403), .A2(W8070), .ZN(O6232));
  NANDX1 G23309 (.A1(W8697), .A2(I1248), .ZN(W32416));
  NANDX1 G23310 (.A1(W30626), .A2(W25330), .ZN(O6230));
  NANDX1 G23311 (.A1(W4378), .A2(W9866), .ZN(O6228));
  NANDX1 G23312 (.A1(W31864), .A2(W5347), .ZN(O6227));
  NANDX1 G23313 (.A1(W1260), .A2(W6216), .ZN(O6226));
  NANDX1 G23314 (.A1(W20497), .A2(W32305), .ZN(W32402));
  NANDX1 G23315 (.A1(W21340), .A2(W12153), .ZN(W32400));
  NANDX1 G23316 (.A1(W21803), .A2(W2208), .ZN(W32399));
  NANDX1 G23317 (.A1(W955), .A2(W26734), .ZN(O6223));
  NANDX1 G23318 (.A1(W6553), .A2(W609), .ZN(O6154));
  NANDX1 G23319 (.A1(W28206), .A2(W27051), .ZN(O6165));
  NANDX1 G23320 (.A1(W5487), .A2(W4983), .ZN(O6164));
  NANDX1 G23321 (.A1(W17996), .A2(I1265), .ZN(W32254));
  NANDX1 G23322 (.A1(W7034), .A2(W4506), .ZN(O6162));
  NANDX1 G23323 (.A1(W31880), .A2(W22337), .ZN(W32250));
  NANDX1 G23324 (.A1(I754), .A2(W4053), .ZN(W32248));
  NANDX1 G23325 (.A1(W20733), .A2(W26973), .ZN(O6159));
  NANDX1 G23326 (.A1(W5033), .A2(I1408), .ZN(W32242));
  NANDX1 G23327 (.A1(W13911), .A2(W31277), .ZN(O6157));
  NANDX1 G23328 (.A1(W1822), .A2(W18359), .ZN(W32236));
  NANDX1 G23329 (.A1(W19137), .A2(W2609), .ZN(W32235));
  NANDX1 G23330 (.A1(W15708), .A2(W27086), .ZN(W32232));
  NANDX1 G23331 (.A1(W17661), .A2(W4547), .ZN(W32258));
  NANDX1 G23332 (.A1(W72), .A2(W7570), .ZN(W32230));
  NANDX1 G23333 (.A1(W21111), .A2(W23027), .ZN(O6152));
  NANDX1 G23334 (.A1(W25134), .A2(W2341), .ZN(O6151));
  NANDX1 G23335 (.A1(W12163), .A2(W29836), .ZN(W32216));
  NANDX1 G23336 (.A1(W30060), .A2(W17856), .ZN(W32213));
  NANDX1 G23337 (.A1(W8850), .A2(W30312), .ZN(W32211));
  NANDX1 G23338 (.A1(W27279), .A2(W20566), .ZN(W32205));
  NANDX1 G23339 (.A1(W2756), .A2(W14638), .ZN(O6143));
  NANDX1 G23340 (.A1(W11798), .A2(W32106), .ZN(O6142));
  NANDX1 G23341 (.A1(W20460), .A2(W15610), .ZN(O6141));
  NANDX1 G23342 (.A1(W17812), .A2(W26539), .ZN(O6137));
  NANDX1 G23343 (.A1(W19065), .A2(W13769), .ZN(W32291));
  NANDX1 G23344 (.A1(I1091), .A2(W31697), .ZN(W32320));
  NANDX1 G23345 (.A1(W30465), .A2(W31884), .ZN(W32318));
  NANDX1 G23346 (.A1(W22104), .A2(W28532), .ZN(O6186));
  NANDX1 G23347 (.A1(W24335), .A2(W10592), .ZN(O6184));
  NANDX1 G23348 (.A1(W20932), .A2(W16187), .ZN(W32306));
  NANDX1 G23349 (.A1(W18869), .A2(W16991), .ZN(W32305));
  NANDX1 G23350 (.A1(W16302), .A2(W1650), .ZN(O6181));
  NANDX1 G23351 (.A1(W19831), .A2(W23219), .ZN(W32299));
  NANDX1 G23352 (.A1(W15124), .A2(W18780), .ZN(O6179));
  NANDX1 G23353 (.A1(W3208), .A2(I78), .ZN(W32293));
  NANDX1 G23354 (.A1(W72), .A2(W28614), .ZN(W32292));
  NANDX1 G23355 (.A1(W32185), .A2(W28221), .ZN(W33049));
  NANDX1 G23356 (.A1(W29627), .A2(W6949), .ZN(W32290));
  NANDX1 G23357 (.A1(W6380), .A2(W16843), .ZN(W32289));
  NANDX1 G23358 (.A1(W30464), .A2(W17627), .ZN(O6175));
  NANDX1 G23359 (.A1(W12157), .A2(W9118), .ZN(W32285));
  NANDX1 G23360 (.A1(W23485), .A2(W3731), .ZN(O6173));
  NANDX1 G23361 (.A1(W16103), .A2(W23097), .ZN(O6172));
  NANDX1 G23362 (.A1(W23493), .A2(W16002), .ZN(O6169));
  NANDX1 G23363 (.A1(W8584), .A2(W13019), .ZN(W32270));
  NANDX1 G23364 (.A1(W8648), .A2(W26871), .ZN(W32269));
  NANDX1 G23365 (.A1(W18231), .A2(W5207), .ZN(W32265));
  NANDX1 G23366 (.A1(W20282), .A2(I539), .ZN(W32263));
  NANDX1 G23367 (.A1(W244), .A2(I1164), .ZN(W33819));
  NANDX1 G23368 (.A1(W1016), .A2(W32323), .ZN(W33864));
  NANDX1 G23369 (.A1(W11960), .A2(W7466), .ZN(O6922));
  NANDX1 G23370 (.A1(W22584), .A2(W29222), .ZN(W33855));
  NANDX1 G23371 (.A1(W20010), .A2(W17253), .ZN(W33853));
  NANDX1 G23372 (.A1(W30376), .A2(W13071), .ZN(O6916));
  NANDX1 G23373 (.A1(W22440), .A2(W4916), .ZN(W33843));
  NANDX1 G23374 (.A1(W20427), .A2(W15012), .ZN(O6914));
  NANDX1 G23375 (.A1(W20531), .A2(W8612), .ZN(W33839));
  NANDX1 G23376 (.A1(W15207), .A2(W17236), .ZN(W33837));
  NANDX1 G23377 (.A1(W8026), .A2(W8661), .ZN(W33834));
  NANDX1 G23378 (.A1(W11680), .A2(W31957), .ZN(W33826));
  NANDX1 G23379 (.A1(W18878), .A2(W7673), .ZN(W33821));
  NANDX1 G23380 (.A1(W23569), .A2(W19563), .ZN(O6923));
  NANDX1 G23381 (.A1(W14418), .A2(I1287), .ZN(O6902));
  NANDX1 G23382 (.A1(W2596), .A2(W6330), .ZN(O6899));
  NANDX1 G23383 (.A1(W13807), .A2(W5915), .ZN(W33811));
  NANDX1 G23384 (.A1(W5891), .A2(W28112), .ZN(O6895));
  NANDX1 G23385 (.A1(W27131), .A2(W29331), .ZN(O6894));
  NANDX1 G23386 (.A1(W11340), .A2(W27027), .ZN(O6893));
  NANDX1 G23387 (.A1(W1407), .A2(W25149), .ZN(O6890));
  NANDX1 G23388 (.A1(W20467), .A2(W2041), .ZN(O6888));
  NANDX1 G23389 (.A1(W7104), .A2(W30173), .ZN(O6886));
  NANDX1 G23390 (.A1(W22558), .A2(W29300), .ZN(O6885));
  NANDX1 G23391 (.A1(W21351), .A2(I721), .ZN(O6883));
  NANDX1 G23392 (.A1(W31090), .A2(W2177), .ZN(O6940));
  NANDX1 G23393 (.A1(W17714), .A2(W23698), .ZN(O6964));
  NANDX1 G23394 (.A1(W26475), .A2(I20), .ZN(O6961));
  NANDX1 G23395 (.A1(W13087), .A2(W30016), .ZN(W33925));
  NANDX1 G23396 (.A1(W1090), .A2(W27640), .ZN(W33921));
  NANDX1 G23397 (.A1(W13467), .A2(W13882), .ZN(W33916));
  NANDX1 G23398 (.A1(W5797), .A2(W32795), .ZN(O6952));
  NANDX1 G23399 (.A1(W31067), .A2(W26350), .ZN(O6950));
  NANDX1 G23400 (.A1(W33005), .A2(W26960), .ZN(O6948));
  NANDX1 G23401 (.A1(W33159), .A2(I966), .ZN(O6947));
  NANDX1 G23402 (.A1(W5237), .A2(W24670), .ZN(W33903));
  NANDX1 G23403 (.A1(W29067), .A2(W5514), .ZN(O6943));
  NANDX1 G23404 (.A1(W15048), .A2(W8895), .ZN(O6942));
  NANDX1 G23405 (.A1(W30786), .A2(W15166), .ZN(O6882));
  NANDX1 G23406 (.A1(W1932), .A2(W22517), .ZN(O6939));
  NANDX1 G23407 (.A1(W13710), .A2(W5626), .ZN(W33887));
  NANDX1 G23408 (.A1(W10633), .A2(W14966), .ZN(O6934));
  NANDX1 G23409 (.A1(I1019), .A2(W12896), .ZN(O6933));
  NANDX1 G23410 (.A1(W20952), .A2(W4082), .ZN(O6932));
  NANDX1 G23411 (.A1(W2413), .A2(W22397), .ZN(O6931));
  NANDX1 G23412 (.A1(W32510), .A2(W12043), .ZN(O6930));
  NANDX1 G23413 (.A1(W17289), .A2(W17917), .ZN(O6927));
  NANDX1 G23414 (.A1(W29375), .A2(W5361), .ZN(O6926));
  NANDX1 G23415 (.A1(W16509), .A2(W15700), .ZN(O6925));
  NANDX1 G23416 (.A1(W1449), .A2(W22132), .ZN(O6924));
  NANDX1 G23417 (.A1(W10359), .A2(W22959), .ZN(O6833));
  NANDX1 G23418 (.A1(W7820), .A2(W26856), .ZN(O6848));
  NANDX1 G23419 (.A1(W27832), .A2(W13642), .ZN(W33714));
  NANDX1 G23420 (.A1(W14118), .A2(W21809), .ZN(O6847));
  NANDX1 G23421 (.A1(W799), .A2(W25519), .ZN(O6845));
  NANDX1 G23422 (.A1(W15684), .A2(W3304), .ZN(O6844));
  NANDX1 G23423 (.A1(W3396), .A2(W10684), .ZN(O6841));
  NANDX1 G23424 (.A1(W8897), .A2(W28342), .ZN(O6840));
  NANDX1 G23425 (.A1(W2373), .A2(W12881), .ZN(W33704));
  NANDX1 G23426 (.A1(W13437), .A2(W2103), .ZN(W33702));
  NANDX1 G23427 (.A1(W31141), .A2(W3891), .ZN(W33701));
  NANDX1 G23428 (.A1(W29231), .A2(W7097), .ZN(W33699));
  NANDX1 G23429 (.A1(W15813), .A2(W23219), .ZN(W33695));
  NANDX1 G23430 (.A1(W18306), .A2(W13973), .ZN(O6849));
  NANDX1 G23431 (.A1(W7675), .A2(W10723), .ZN(W33685));
  NANDX1 G23432 (.A1(W8372), .A2(W16905), .ZN(O6829));
  NANDX1 G23433 (.A1(I108), .A2(W13647), .ZN(O6826));
  NANDX1 G23434 (.A1(W21588), .A2(W9279), .ZN(O6823));
  NANDX1 G23435 (.A1(W16905), .A2(W25992), .ZN(W33671));
  NANDX1 G23436 (.A1(W27064), .A2(W10479), .ZN(W33669));
  NANDX1 G23437 (.A1(W10167), .A2(W5164), .ZN(O6821));
  NANDX1 G23438 (.A1(W30194), .A2(W7122), .ZN(O6819));
  NANDX1 G23439 (.A1(W28645), .A2(W6539), .ZN(O6817));
  NANDX1 G23440 (.A1(W28413), .A2(W25364), .ZN(O6816));
  NANDX1 G23441 (.A1(W10986), .A2(W8516), .ZN(O6815));
  NANDX1 G23442 (.A1(W33256), .A2(W1978), .ZN(O6864));
  NANDX1 G23443 (.A1(W3858), .A2(W6423), .ZN(W33781));
  NANDX1 G23444 (.A1(W5198), .A2(W15093), .ZN(O6876));
  NANDX1 G23445 (.A1(W27290), .A2(W12548), .ZN(W33774));
  NANDX1 G23446 (.A1(I1918), .A2(W13546), .ZN(O6873));
  NANDX1 G23447 (.A1(W32745), .A2(W3771), .ZN(O6872));
  NANDX1 G23448 (.A1(W11624), .A2(W993), .ZN(W33764));
  NANDX1 G23449 (.A1(W11477), .A2(W2090), .ZN(O6868));
  NANDX1 G23450 (.A1(W17182), .A2(W1755), .ZN(W33761));
  NANDX1 G23451 (.A1(W10648), .A2(W4030), .ZN(W33755));
  NANDX1 G23452 (.A1(I277), .A2(W28707), .ZN(W33754));
  NANDX1 G23453 (.A1(W1244), .A2(W27438), .ZN(O6865));
  NANDX1 G23454 (.A1(W19324), .A2(I413), .ZN(W33934));
  NANDX1 G23455 (.A1(W2705), .A2(W5589), .ZN(W33742));
  NANDX1 G23456 (.A1(W26567), .A2(I1324), .ZN(W33741));
  NANDX1 G23457 (.A1(W26083), .A2(W25740), .ZN(O6862));
  NANDX1 G23458 (.A1(W18731), .A2(W5623), .ZN(O6860));
  NANDX1 G23459 (.A1(W3879), .A2(W2421), .ZN(O6856));
  NANDX1 G23460 (.A1(W25724), .A2(W24732), .ZN(O6855));
  NANDX1 G23461 (.A1(W14004), .A2(W31), .ZN(W33728));
  NANDX1 G23462 (.A1(W7459), .A2(W6606), .ZN(W33726));
  NANDX1 G23463 (.A1(W425), .A2(W2242), .ZN(O6852));
  NANDX1 G23464 (.A1(W29066), .A2(W31230), .ZN(W33722));
  NANDX1 G23465 (.A1(I1503), .A2(W26575), .ZN(O6851));
  NANDX1 G23466 (.A1(W14733), .A2(I1949), .ZN(O7062));
  NANDX1 G23467 (.A1(W22424), .A2(W3100), .ZN(W34120));
  NANDX1 G23468 (.A1(W14249), .A2(W11), .ZN(O7074));
  NANDX1 G23469 (.A1(W30544), .A2(W6813), .ZN(O7070));
  NANDX1 G23470 (.A1(W21337), .A2(W17316), .ZN(W34106));
  NANDX1 G23471 (.A1(W10641), .A2(W8309), .ZN(O7068));
  NANDX1 G23472 (.A1(W14331), .A2(W29041), .ZN(O7067));
  NANDX1 G23473 (.A1(W14475), .A2(W15070), .ZN(W34100));
  NANDX1 G23474 (.A1(W10169), .A2(W24221), .ZN(W34099));
  NANDX1 G23475 (.A1(W13638), .A2(W326), .ZN(O7064));
  NANDX1 G23476 (.A1(W29569), .A2(W21079), .ZN(O7063));
  NANDX1 G23477 (.A1(W1363), .A2(W26975), .ZN(W34094));
  NANDX1 G23478 (.A1(W30596), .A2(W15274), .ZN(W34092));
  NANDX1 G23479 (.A1(I1149), .A2(W30382), .ZN(W34128));
  NANDX1 G23480 (.A1(W1815), .A2(W6411), .ZN(W34088));
  NANDX1 G23481 (.A1(W11535), .A2(W8716), .ZN(O7061));
  NANDX1 G23482 (.A1(W28154), .A2(W30172), .ZN(W34083));
  NANDX1 G23483 (.A1(W17332), .A2(I594), .ZN(O7058));
  NANDX1 G23484 (.A1(W5176), .A2(W20698), .ZN(O7055));
  NANDX1 G23485 (.A1(W1736), .A2(W12053), .ZN(W34075));
  NANDX1 G23486 (.A1(W23607), .A2(W12118), .ZN(O7053));
  NANDX1 G23487 (.A1(I1374), .A2(W26428), .ZN(O7050));
  NANDX1 G23488 (.A1(W22005), .A2(I48), .ZN(W34066));
  NANDX1 G23489 (.A1(W25362), .A2(W2745), .ZN(O7047));
  NANDX1 G23490 (.A1(W16466), .A2(W16919), .ZN(O7042));
  NANDX1 G23491 (.A1(W3173), .A2(W13050), .ZN(W34167));
  NANDX1 G23492 (.A1(W14494), .A2(W6597), .ZN(O7117));
  NANDX1 G23493 (.A1(W18791), .A2(W26606), .ZN(W34195));
  NANDX1 G23494 (.A1(W10777), .A2(W7491), .ZN(W34194));
  NANDX1 G23495 (.A1(W11421), .A2(W18692), .ZN(W34186));
  NANDX1 G23496 (.A1(W10037), .A2(W33399), .ZN(O7113));
  NANDX1 G23497 (.A1(W23554), .A2(W18503), .ZN(W34183));
  NANDX1 G23498 (.A1(W33403), .A2(W4556), .ZN(W34179));
  NANDX1 G23499 (.A1(W32457), .A2(W22450), .ZN(O7109));
  NANDX1 G23500 (.A1(W16234), .A2(W6354), .ZN(O7105));
  NANDX1 G23501 (.A1(W23121), .A2(W32766), .ZN(O7104));
  NANDX1 G23502 (.A1(I1569), .A2(W20251), .ZN(W34170));
  NANDX1 G23503 (.A1(W31959), .A2(W23516), .ZN(W34168));
  NANDX1 G23504 (.A1(W16823), .A2(W28879), .ZN(O7040));
  NANDX1 G23505 (.A1(W21931), .A2(W10410), .ZN(W34165));
  NANDX1 G23506 (.A1(W33039), .A2(W19682), .ZN(O7102));
  NANDX1 G23507 (.A1(W12782), .A2(W31698), .ZN(O7094));
  NANDX1 G23508 (.A1(W15777), .A2(W13390), .ZN(O7093));
  NANDX1 G23509 (.A1(W28002), .A2(W24733), .ZN(W34144));
  NANDX1 G23510 (.A1(W32199), .A2(W23871), .ZN(O7088));
  NANDX1 G23511 (.A1(W29358), .A2(W12076), .ZN(O7087));
  NANDX1 G23512 (.A1(W20631), .A2(W24028), .ZN(W34136));
  NANDX1 G23513 (.A1(W23395), .A2(W14868), .ZN(O7084));
  NANDX1 G23514 (.A1(W24551), .A2(W29790), .ZN(O7082));
  NANDX1 G23515 (.A1(W15633), .A2(I61), .ZN(W34129));
  NANDX1 G23516 (.A1(W25985), .A2(W12408), .ZN(W33967));
  NANDX1 G23517 (.A1(W22048), .A2(W11175), .ZN(O7006));
  NANDX1 G23518 (.A1(I1120), .A2(I1221), .ZN(W34000));
  NANDX1 G23519 (.A1(W17283), .A2(W6687), .ZN(O7004));
  NANDX1 G23520 (.A1(W21441), .A2(W6114), .ZN(O7003));
  NANDX1 G23521 (.A1(W3354), .A2(W19552), .ZN(W33994));
  NANDX1 G23522 (.A1(W32177), .A2(W26618), .ZN(W33992));
  NANDX1 G23523 (.A1(W338), .A2(I71), .ZN(O6998));
  NANDX1 G23524 (.A1(W6070), .A2(W590), .ZN(O6996));
  NANDX1 G23525 (.A1(W24996), .A2(W27005), .ZN(W33983));
  NANDX1 G23526 (.A1(W14564), .A2(W25583), .ZN(O6993));
  NANDX1 G23527 (.A1(W4029), .A2(W28586), .ZN(O6991));
  NANDX1 G23528 (.A1(W1542), .A2(W32781), .ZN(O6987));
  NANDX1 G23529 (.A1(W11814), .A2(W15281), .ZN(W34004));
  NANDX1 G23530 (.A1(W11404), .A2(W12683), .ZN(W33966));
  NANDX1 G23531 (.A1(W241), .A2(W33177), .ZN(W33961));
  NANDX1 G23532 (.A1(W7863), .A2(W19595), .ZN(O6980));
  NANDX1 G23533 (.A1(W2812), .A2(W955), .ZN(W33958));
  NANDX1 G23534 (.A1(W11149), .A2(W11367), .ZN(O6973));
  NANDX1 G23535 (.A1(W25080), .A2(W33117), .ZN(O6971));
  NANDX1 G23536 (.A1(W2518), .A2(W10194), .ZN(O6970));
  NANDX1 G23537 (.A1(W14452), .A2(W26205), .ZN(W33944));
  NANDX1 G23538 (.A1(W3028), .A2(W22353), .ZN(W33942));
  NANDX1 G23539 (.A1(W29092), .A2(W26706), .ZN(W33938));
  NANDX1 G23540 (.A1(W5432), .A2(W9236), .ZN(W33936));
  NANDX1 G23541 (.A1(W10102), .A2(I128), .ZN(W34035));
  NANDX1 G23542 (.A1(W27248), .A2(W4709), .ZN(O7039));
  NANDX1 G23543 (.A1(W252), .A2(W7048), .ZN(O7038));
  NANDX1 G23544 (.A1(W7543), .A2(I282), .ZN(W34053));
  NANDX1 G23545 (.A1(W13164), .A2(W18944), .ZN(W34048));
  NANDX1 G23546 (.A1(W28441), .A2(W19379), .ZN(W34047));
  NANDX1 G23547 (.A1(W6923), .A2(W1263), .ZN(O7034));
  NANDX1 G23548 (.A1(W24466), .A2(W13786), .ZN(O7031));
  NANDX1 G23549 (.A1(W13295), .A2(W626), .ZN(W34040));
  NANDX1 G23550 (.A1(I1256), .A2(W931), .ZN(O7030));
  NANDX1 G23551 (.A1(W9942), .A2(W20818), .ZN(W34037));
  NANDX1 G23552 (.A1(W14349), .A2(W15541), .ZN(O7028));
  NANDX1 G23553 (.A1(W15982), .A2(W31462), .ZN(O6811));
  NANDX1 G23554 (.A1(W27024), .A2(W10540), .ZN(W34032));
  NANDX1 G23555 (.A1(W8581), .A2(W33810), .ZN(O7026));
  NANDX1 G23556 (.A1(W4017), .A2(W7621), .ZN(W34030));
  NANDX1 G23557 (.A1(W5501), .A2(W8751), .ZN(W34024));
  NANDX1 G23558 (.A1(W8613), .A2(W9291), .ZN(O7020));
  NANDX1 G23559 (.A1(W15902), .A2(I1222), .ZN(O7018));
  NANDX1 G23560 (.A1(W20247), .A2(W33434), .ZN(W34014));
  NANDX1 G23561 (.A1(W4698), .A2(W29939), .ZN(O7011));
  NANDX1 G23562 (.A1(W13886), .A2(W957), .ZN(O7010));
  NANDX1 G23563 (.A1(I583), .A2(W31492), .ZN(O7009));
  NANDX1 G23564 (.A1(W24262), .A2(W27152), .ZN(O7008));
  NANDX1 G23565 (.A1(W4154), .A2(I416), .ZN(W33262));
  NANDX1 G23566 (.A1(W1375), .A2(W8450), .ZN(O6631));
  NANDX1 G23567 (.A1(W8163), .A2(W1767), .ZN(W33281));
  NANDX1 G23568 (.A1(W5340), .A2(W1649), .ZN(W33280));
  NANDX1 G23569 (.A1(W29496), .A2(W4949), .ZN(O6630));
  NANDX1 G23570 (.A1(W21343), .A2(W26114), .ZN(W33276));
  NANDX1 G23571 (.A1(I1557), .A2(W6712), .ZN(W33274));
  NANDX1 G23572 (.A1(W27643), .A2(W14646), .ZN(W33273));
  NANDX1 G23573 (.A1(W24108), .A2(W9037), .ZN(W33272));
  NANDX1 G23574 (.A1(W21367), .A2(W14903), .ZN(W33271));
  NANDX1 G23575 (.A1(W7499), .A2(W6985), .ZN(O6629));
  NANDX1 G23576 (.A1(W28461), .A2(W673), .ZN(W33268));
  NANDX1 G23577 (.A1(W15625), .A2(W19004), .ZN(W33264));
  NANDX1 G23578 (.A1(W2003), .A2(W12589), .ZN(O6632));
  NANDX1 G23579 (.A1(W7976), .A2(W30268), .ZN(O6626));
  NANDX1 G23580 (.A1(W32280), .A2(W22125), .ZN(O6625));
  NANDX1 G23581 (.A1(W30281), .A2(W27893), .ZN(W33256));
  NANDX1 G23582 (.A1(W2711), .A2(W20962), .ZN(O6622));
  NANDX1 G23583 (.A1(W17001), .A2(W875), .ZN(W33254));
  NANDX1 G23584 (.A1(W11453), .A2(I1672), .ZN(W33242));
  NANDX1 G23585 (.A1(I825), .A2(I418), .ZN(O6614));
  NANDX1 G23586 (.A1(W30028), .A2(W22978), .ZN(W33238));
  NANDX1 G23587 (.A1(W11490), .A2(W25941), .ZN(O6608));
  NANDX1 G23588 (.A1(W15828), .A2(W22985), .ZN(O6605));
  NANDX1 G23589 (.A1(I1116), .A2(W18291), .ZN(O6604));
  NANDX1 G23590 (.A1(W22575), .A2(W24206), .ZN(W33311));
  NANDX1 G23591 (.A1(W9918), .A2(W16881), .ZN(O6663));
  NANDX1 G23592 (.A1(W16565), .A2(W23568), .ZN(W33348));
  NANDX1 G23593 (.A1(W10340), .A2(W21775), .ZN(O6662));
  NANDX1 G23594 (.A1(W8130), .A2(W33073), .ZN(O6659));
  NANDX1 G23595 (.A1(W22391), .A2(W27920), .ZN(W33338));
  NANDX1 G23596 (.A1(W7347), .A2(W3949), .ZN(O6654));
  NANDX1 G23597 (.A1(W16006), .A2(W2170), .ZN(O6650));
  NANDX1 G23598 (.A1(W19518), .A2(W6867), .ZN(W33323));
  NANDX1 G23599 (.A1(W6610), .A2(W16506), .ZN(O6643));
  NANDX1 G23600 (.A1(W28696), .A2(W233), .ZN(W33314));
  NANDX1 G23601 (.A1(W2980), .A2(W589), .ZN(O6642));
  NANDX1 G23602 (.A1(W11832), .A2(W1834), .ZN(W33312));
  NANDX1 G23603 (.A1(W13627), .A2(W971), .ZN(O6602));
  NANDX1 G23604 (.A1(W12043), .A2(W19454), .ZN(O6641));
  NANDX1 G23605 (.A1(W22014), .A2(W31518), .ZN(W33308));
  NANDX1 G23606 (.A1(W15425), .A2(W18237), .ZN(O6640));
  NANDX1 G23607 (.A1(W25256), .A2(W21667), .ZN(O6638));
  NANDX1 G23608 (.A1(W7316), .A2(W30991), .ZN(W33301));
  NANDX1 G23609 (.A1(W33170), .A2(W22440), .ZN(W33300));
  NANDX1 G23610 (.A1(W14578), .A2(W19641), .ZN(W33299));
  NANDX1 G23611 (.A1(W4488), .A2(W3600), .ZN(W33291));
  NANDX1 G23612 (.A1(W27252), .A2(W1075), .ZN(W33288));
  NANDX1 G23613 (.A1(W11250), .A2(W24699), .ZN(O6634));
  NANDX1 G23614 (.A1(W21848), .A2(W3720), .ZN(O6633));
  NANDX1 G23615 (.A1(W3426), .A2(W15115), .ZN(W33086));
  NANDX1 G23616 (.A1(W15628), .A2(W28363), .ZN(W33122));
  NANDX1 G23617 (.A1(W6526), .A2(W20416), .ZN(O6555));
  NANDX1 G23618 (.A1(W2140), .A2(W11561), .ZN(W33117));
  NANDX1 G23619 (.A1(W27833), .A2(W10799), .ZN(O6552));
  NANDX1 G23620 (.A1(W24176), .A2(W28491), .ZN(O6548));
  NANDX1 G23621 (.A1(W7662), .A2(W3364), .ZN(O6547));
  NANDX1 G23622 (.A1(W6151), .A2(W1562), .ZN(O6545));
  NANDX1 G23623 (.A1(W17847), .A2(W29928), .ZN(W33105));
  NANDX1 G23624 (.A1(W31771), .A2(W25891), .ZN(W33101));
  NANDX1 G23625 (.A1(I734), .A2(W4910), .ZN(O6541));
  NANDX1 G23626 (.A1(W20526), .A2(W17393), .ZN(O6540));
  NANDX1 G23627 (.A1(W16400), .A2(W22803), .ZN(W33093));
  NANDX1 G23628 (.A1(W31197), .A2(W31587), .ZN(W33128));
  NANDX1 G23629 (.A1(W31504), .A2(W16174), .ZN(W33085));
  NANDX1 G23630 (.A1(W2298), .A2(W19146), .ZN(W33078));
  NANDX1 G23631 (.A1(W19186), .A2(W9197), .ZN(W33077));
  NANDX1 G23632 (.A1(I1750), .A2(W9295), .ZN(O6529));
  NANDX1 G23633 (.A1(W11440), .A2(W989), .ZN(O6528));
  NANDX1 G23634 (.A1(W5906), .A2(W5308), .ZN(W33070));
  NANDX1 G23635 (.A1(W4752), .A2(W20200), .ZN(W33064));
  NANDX1 G23636 (.A1(W11185), .A2(W18679), .ZN(W33060));
  NANDX1 G23637 (.A1(W13743), .A2(W3792), .ZN(O6524));
  NANDX1 G23638 (.A1(W18075), .A2(W22851), .ZN(O6522));
  NANDX1 G23639 (.A1(I712), .A2(W16723), .ZN(W33055));
  NANDX1 G23640 (.A1(W10127), .A2(I1935), .ZN(W33161));
  NANDX1 G23641 (.A1(W16893), .A2(W18157), .ZN(W33211));
  NANDX1 G23642 (.A1(W28622), .A2(W7849), .ZN(W33205));
  NANDX1 G23643 (.A1(W19855), .A2(W14854), .ZN(W33200));
  NANDX1 G23644 (.A1(W2076), .A2(W4929), .ZN(O6586));
  NANDX1 G23645 (.A1(W4573), .A2(W16463), .ZN(W33186));
  NANDX1 G23646 (.A1(W27340), .A2(W28596), .ZN(O6578));
  NANDX1 G23647 (.A1(W28217), .A2(W7968), .ZN(W33174));
  NANDX1 G23648 (.A1(W16993), .A2(W15674), .ZN(W33172));
  NANDX1 G23649 (.A1(W10986), .A2(W21168), .ZN(O6577));
  NANDX1 G23650 (.A1(W10644), .A2(W27648), .ZN(O6576));
  NANDX1 G23651 (.A1(W26929), .A2(W1965), .ZN(O6575));
  NANDX1 G23652 (.A1(W18913), .A2(W27107), .ZN(O6665));
  NANDX1 G23653 (.A1(W20545), .A2(W29630), .ZN(W33159));
  NANDX1 G23654 (.A1(W25951), .A2(W29571), .ZN(O6570));
  NANDX1 G23655 (.A1(W25800), .A2(W22644), .ZN(W33154));
  NANDX1 G23656 (.A1(W10877), .A2(W28647), .ZN(O6568));
  NANDX1 G23657 (.A1(W13924), .A2(W28375), .ZN(O6567));
  NANDX1 G23658 (.A1(W30321), .A2(W26095), .ZN(W33147));
  NANDX1 G23659 (.A1(W583), .A2(W22931), .ZN(O6564));
  NANDX1 G23660 (.A1(W22776), .A2(W31113), .ZN(W33137));
  NANDX1 G23661 (.A1(W21910), .A2(W20719), .ZN(O6562));
  NANDX1 G23662 (.A1(W1502), .A2(W15739), .ZN(W33133));
  NANDX1 G23663 (.A1(W7954), .A2(W16402), .ZN(O6559));
  NANDX1 G23664 (.A1(W26714), .A2(W23753), .ZN(O6754));
  NANDX1 G23665 (.A1(W31120), .A2(W16571), .ZN(W33575));
  NANDX1 G23666 (.A1(W10655), .A2(W7182), .ZN(W33574));
  NANDX1 G23667 (.A1(W2671), .A2(W23470), .ZN(O6763));
  NANDX1 G23668 (.A1(W805), .A2(W1644), .ZN(W33558));
  NANDX1 G23669 (.A1(W17190), .A2(W18159), .ZN(W33557));
  NANDX1 G23670 (.A1(W20055), .A2(W3881), .ZN(O6760));
  NANDX1 G23671 (.A1(W14658), .A2(W23091), .ZN(O6759));
  NANDX1 G23672 (.A1(W280), .A2(W29600), .ZN(O6758));
  NANDX1 G23673 (.A1(W495), .A2(W19028), .ZN(W33551));
  NANDX1 G23674 (.A1(W23306), .A2(W11520), .ZN(O6757));
  NANDX1 G23675 (.A1(W25379), .A2(W19427), .ZN(O6756));
  NANDX1 G23676 (.A1(W24744), .A2(W7396), .ZN(W33547));
  NANDX1 G23677 (.A1(W1555), .A2(W19609), .ZN(W33577));
  NANDX1 G23678 (.A1(W8745), .A2(W26251), .ZN(O6752));
  NANDX1 G23679 (.A1(W32388), .A2(W33266), .ZN(O6749));
  NANDX1 G23680 (.A1(W19259), .A2(W2925), .ZN(W33535));
  NANDX1 G23681 (.A1(W25874), .A2(W23242), .ZN(O6747));
  NANDX1 G23682 (.A1(W30376), .A2(W33457), .ZN(W33527));
  NANDX1 G23683 (.A1(W14599), .A2(W344), .ZN(O6744));
  NANDX1 G23684 (.A1(W13114), .A2(W16161), .ZN(W33525));
  NANDX1 G23685 (.A1(W10390), .A2(W9558), .ZN(O6742));
  NANDX1 G23686 (.A1(W23000), .A2(W4764), .ZN(W33518));
  NANDX1 G23687 (.A1(W29039), .A2(W13490), .ZN(O6740));
  NANDX1 G23688 (.A1(W10908), .A2(W5705), .ZN(O6738));
  NANDX1 G23689 (.A1(W13827), .A2(W10719), .ZN(W33613));
  NANDX1 G23690 (.A1(W24588), .A2(W25040), .ZN(O6808));
  NANDX1 G23691 (.A1(W16675), .A2(W33332), .ZN(O6806));
  NANDX1 G23692 (.A1(W3278), .A2(W22239), .ZN(W33645));
  NANDX1 G23693 (.A1(W19358), .A2(W11652), .ZN(W33644));
  NANDX1 G23694 (.A1(W19904), .A2(I202), .ZN(O6804));
  NANDX1 G23695 (.A1(W16264), .A2(W11896), .ZN(W33635));
  NANDX1 G23696 (.A1(W23074), .A2(W9892), .ZN(O6797));
  NANDX1 G23697 (.A1(W23756), .A2(W15242), .ZN(W33624));
  NANDX1 G23698 (.A1(W19924), .A2(W13595), .ZN(W33623));
  NANDX1 G23699 (.A1(W10901), .A2(W11677), .ZN(W33619));
  NANDX1 G23700 (.A1(W7073), .A2(W16851), .ZN(O6788));
  NANDX1 G23701 (.A1(W23921), .A2(W8218), .ZN(O6737));
  NANDX1 G23702 (.A1(W25065), .A2(W15166), .ZN(W33612));
  NANDX1 G23703 (.A1(W24), .A2(W11878), .ZN(W33609));
  NANDX1 G23704 (.A1(W19019), .A2(W21605), .ZN(O6782));
  NANDX1 G23705 (.A1(W2947), .A2(W16166), .ZN(O6781));
  NANDX1 G23706 (.A1(W11695), .A2(W1539), .ZN(O6780));
  NANDX1 G23707 (.A1(W7825), .A2(W5532), .ZN(O6775));
  NANDX1 G23708 (.A1(W16959), .A2(I1069), .ZN(O6771));
  NANDX1 G23709 (.A1(W9364), .A2(W32762), .ZN(O6770));
  NANDX1 G23710 (.A1(W16670), .A2(W14096), .ZN(W33584));
  NANDX1 G23711 (.A1(W24811), .A2(W150), .ZN(O6769));
  NANDX1 G23712 (.A1(W8910), .A2(W2224), .ZN(O6768));
  NANDX1 G23713 (.A1(W15726), .A2(W5168), .ZN(W33399));
  NANDX1 G23714 (.A1(W24906), .A2(W10445), .ZN(O6701));
  NANDX1 G23715 (.A1(W11517), .A2(W21157), .ZN(O6700));
  NANDX1 G23716 (.A1(W13306), .A2(W5708), .ZN(O6698));
  NANDX1 G23717 (.A1(W15581), .A2(W11339), .ZN(W33425));
  NANDX1 G23718 (.A1(W12347), .A2(W21712), .ZN(W33424));
  NANDX1 G23719 (.A1(W32006), .A2(W4585), .ZN(W33422));
  NANDX1 G23720 (.A1(W25972), .A2(W28808), .ZN(O6690));
  NANDX1 G23721 (.A1(W7661), .A2(W10640), .ZN(W33411));
  NANDX1 G23722 (.A1(W7441), .A2(W33172), .ZN(O6686));
  NANDX1 G23723 (.A1(W28650), .A2(W31357), .ZN(W33409));
  NANDX1 G23724 (.A1(W29809), .A2(W4066), .ZN(W33407));
  NANDX1 G23725 (.A1(W29509), .A2(W7433), .ZN(W33401));
  NANDX1 G23726 (.A1(W3770), .A2(W14372), .ZN(O6703));
  NANDX1 G23727 (.A1(W1312), .A2(W16690), .ZN(O6684));
  NANDX1 G23728 (.A1(W26355), .A2(W15791), .ZN(W33394));
  NANDX1 G23729 (.A1(I1994), .A2(W23416), .ZN(W33389));
  NANDX1 G23730 (.A1(I112), .A2(W2072), .ZN(O6677));
  NANDX1 G23731 (.A1(W513), .A2(W11391), .ZN(W33379));
  NANDX1 G23732 (.A1(W7446), .A2(W4044), .ZN(W33375));
  NANDX1 G23733 (.A1(W21237), .A2(W10513), .ZN(W33373));
  NANDX1 G23734 (.A1(W12363), .A2(W6053), .ZN(W33369));
  NANDX1 G23735 (.A1(W17053), .A2(W8651), .ZN(W33365));
  NANDX1 G23736 (.A1(W29695), .A2(I489), .ZN(W33364));
  NANDX1 G23737 (.A1(W8983), .A2(W2320), .ZN(O6666));
  NANDX1 G23738 (.A1(W8825), .A2(W12495), .ZN(O6718));
  NANDX1 G23739 (.A1(W30183), .A2(W20874), .ZN(O6733));
  NANDX1 G23740 (.A1(W18206), .A2(I40), .ZN(W33499));
  NANDX1 G23741 (.A1(W29669), .A2(W14660), .ZN(W33498));
  NANDX1 G23742 (.A1(W25251), .A2(W15982), .ZN(W33497));
  NANDX1 G23743 (.A1(W7224), .A2(W14482), .ZN(O6732));
  NANDX1 G23744 (.A1(W251), .A2(W32575), .ZN(W33488));
  NANDX1 G23745 (.A1(W9396), .A2(W2479), .ZN(O6728));
  NANDX1 G23746 (.A1(W16207), .A2(W6247), .ZN(W33486));
  NANDX1 G23747 (.A1(W15389), .A2(W31811), .ZN(W33485));
  NANDX1 G23748 (.A1(I808), .A2(W22356), .ZN(O6726));
  NANDX1 G23749 (.A1(W32725), .A2(W6793), .ZN(O6723));
  NANDX1 G23750 (.A1(W10119), .A2(W9786), .ZN(O8430));
  NANDX1 G23751 (.A1(W29624), .A2(W31072), .ZN(O6717));
  NANDX1 G23752 (.A1(W11547), .A2(W10424), .ZN(O6716));
  NANDX1 G23753 (.A1(W18283), .A2(W10989), .ZN(W33466));
  NANDX1 G23754 (.A1(W19531), .A2(W31496), .ZN(O6714));
  NANDX1 G23755 (.A1(W14735), .A2(W14640), .ZN(W33463));
  NANDX1 G23756 (.A1(W4137), .A2(W19025), .ZN(W33461));
  NANDX1 G23757 (.A1(I1337), .A2(W9427), .ZN(O6712));
  NANDX1 G23758 (.A1(W24633), .A2(W12303), .ZN(W33457));
  NANDX1 G23759 (.A1(W9283), .A2(W31052), .ZN(O6707));
  NANDX1 G23760 (.A1(W24203), .A2(W2858), .ZN(W33448));
  NANDX1 G23761 (.A1(W3492), .A2(W11710), .ZN(W33447));
  NANDX1 G23762 (.A1(W9441), .A2(W35767), .ZN(O10434));
  NANDX1 G23763 (.A1(W30472), .A2(W33900), .ZN(W39790));
  NANDX1 G23764 (.A1(W39397), .A2(W9533), .ZN(W39785));
  NANDX1 G23765 (.A1(W7230), .A2(W21713), .ZN(O10446));
  NANDX1 G23766 (.A1(W20456), .A2(W17037), .ZN(O10445));
  NANDX1 G23767 (.A1(W31927), .A2(W9306), .ZN(O10443));
  NANDX1 G23768 (.A1(I1378), .A2(W12008), .ZN(W39778));
  NANDX1 G23769 (.A1(W26166), .A2(W39545), .ZN(O10442));
  NANDX1 G23770 (.A1(W35981), .A2(W31901), .ZN(O10440));
  NANDX1 G23771 (.A1(W20283), .A2(W31216), .ZN(O10439));
  NANDX1 G23772 (.A1(W11260), .A2(W3136), .ZN(O10437));
  NANDX1 G23773 (.A1(W2819), .A2(W14377), .ZN(W39764));
  NANDX1 G23774 (.A1(W12187), .A2(W20224), .ZN(W39762));
  NANDX1 G23775 (.A1(W8338), .A2(W12762), .ZN(O10450));
  NANDX1 G23776 (.A1(W9674), .A2(W18273), .ZN(O10424));
  NANDX1 G23777 (.A1(W4829), .A2(W29836), .ZN(O10422));
  NANDX1 G23778 (.A1(W5464), .A2(W21942), .ZN(O10419));
  NANDX1 G23779 (.A1(W2394), .A2(W30432), .ZN(O10418));
  NANDX1 G23780 (.A1(W10416), .A2(W1059), .ZN(W39736));
  NANDX1 G23781 (.A1(I999), .A2(W22172), .ZN(O10412));
  NANDX1 G23782 (.A1(W30020), .A2(W19403), .ZN(O10411));
  NANDX1 G23783 (.A1(W27326), .A2(W13559), .ZN(O10410));
  NANDX1 G23784 (.A1(W39208), .A2(W16939), .ZN(W39728));
  NANDX1 G23785 (.A1(W4220), .A2(W683), .ZN(W39725));
  NANDX1 G23786 (.A1(W9937), .A2(W39133), .ZN(W39714));
  NANDX1 G23787 (.A1(W10704), .A2(W34305), .ZN(O10474));
  NANDX1 G23788 (.A1(W32256), .A2(W35247), .ZN(O10515));
  NANDX1 G23789 (.A1(W3557), .A2(W3509), .ZN(O10514));
  NANDX1 G23790 (.A1(W7429), .A2(W5544), .ZN(W39871));
  NANDX1 G23791 (.A1(W15856), .A2(W32740), .ZN(O10513));
  NANDX1 G23792 (.A1(W7963), .A2(W18100), .ZN(O10509));
  NANDX1 G23793 (.A1(W28653), .A2(W34041), .ZN(O10503));
  NANDX1 G23794 (.A1(W31761), .A2(W3605), .ZN(O10500));
  NANDX1 G23795 (.A1(W29757), .A2(W30172), .ZN(O10494));
  NANDX1 G23796 (.A1(W3948), .A2(W21453), .ZN(O10492));
  NANDX1 G23797 (.A1(W18837), .A2(W33473), .ZN(W39840));
  NANDX1 G23798 (.A1(W9625), .A2(W10579), .ZN(O10484));
  NANDX1 G23799 (.A1(W214), .A2(W23518), .ZN(O10475));
  NANDX1 G23800 (.A1(W21758), .A2(W19927), .ZN(O10399));
  NANDX1 G23801 (.A1(W4445), .A2(W24020), .ZN(O10472));
  NANDX1 G23802 (.A1(I844), .A2(W35227), .ZN(O10471));
  NANDX1 G23803 (.A1(W16110), .A2(W11236), .ZN(O10469));
  NANDX1 G23804 (.A1(W35105), .A2(W13591), .ZN(O10467));
  NANDX1 G23805 (.A1(W2564), .A2(W34866), .ZN(O10466));
  NANDX1 G23806 (.A1(W14961), .A2(W26749), .ZN(O10464));
  NANDX1 G23807 (.A1(W22272), .A2(W11772), .ZN(O10463));
  NANDX1 G23808 (.A1(W6618), .A2(W33934), .ZN(W39807));
  NANDX1 G23809 (.A1(W19081), .A2(W32619), .ZN(O10461));
  NANDX1 G23810 (.A1(W17894), .A2(W33517), .ZN(O10456));
  NANDX1 G23811 (.A1(W6463), .A2(W12583), .ZN(O10455));
  NANDX1 G23812 (.A1(W7834), .A2(W6903), .ZN(O10315));
  NANDX1 G23813 (.A1(W33161), .A2(W1940), .ZN(O10335));
  NANDX1 G23814 (.A1(W9428), .A2(W18017), .ZN(O10332));
  NANDX1 G23815 (.A1(W18339), .A2(W32122), .ZN(W39611));
  NANDX1 G23816 (.A1(W2876), .A2(W14806), .ZN(O10330));
  NANDX1 G23817 (.A1(W28727), .A2(W34838), .ZN(O10329));
  NANDX1 G23818 (.A1(W2823), .A2(W20578), .ZN(O10328));
  NANDX1 G23819 (.A1(W29916), .A2(W38932), .ZN(O10327));
  NANDX1 G23820 (.A1(W35755), .A2(W12455), .ZN(O10326));
  NANDX1 G23821 (.A1(W4135), .A2(W36453), .ZN(W39605));
  NANDX1 G23822 (.A1(W21635), .A2(W16535), .ZN(O10322));
  NANDX1 G23823 (.A1(W2820), .A2(W2523), .ZN(O10317));
  NANDX1 G23824 (.A1(W30094), .A2(W11465), .ZN(O10316));
  NANDX1 G23825 (.A1(W21073), .A2(W10788), .ZN(W39618));
  NANDX1 G23826 (.A1(W11078), .A2(W34766), .ZN(O10313));
  NANDX1 G23827 (.A1(W32217), .A2(W14567), .ZN(W39587));
  NANDX1 G23828 (.A1(W21951), .A2(W4699), .ZN(O10310));
  NANDX1 G23829 (.A1(I968), .A2(W20142), .ZN(O10309));
  NANDX1 G23830 (.A1(W39202), .A2(W12936), .ZN(O10307));
  NANDX1 G23831 (.A1(W8673), .A2(W20073), .ZN(W39574));
  NANDX1 G23832 (.A1(W17122), .A2(W16759), .ZN(W39572));
  NANDX1 G23833 (.A1(W26820), .A2(W16351), .ZN(O10299));
  NANDX1 G23834 (.A1(W11938), .A2(W17421), .ZN(W39566));
  NANDX1 G23835 (.A1(W31881), .A2(W32347), .ZN(O10296));
  NANDX1 G23836 (.A1(W11372), .A2(W7338), .ZN(O10294));
  NANDX1 G23837 (.A1(W28003), .A2(W19024), .ZN(O10373));
  NANDX1 G23838 (.A1(W25216), .A2(W6628), .ZN(O10398));
  NANDX1 G23839 (.A1(W21115), .A2(W16908), .ZN(O10395));
  NANDX1 G23840 (.A1(W31181), .A2(W26570), .ZN(O10393));
  NANDX1 G23841 (.A1(W3676), .A2(W7534), .ZN(O10387));
  NANDX1 G23842 (.A1(W34447), .A2(W37261), .ZN(O10386));
  NANDX1 G23843 (.A1(W2245), .A2(W33097), .ZN(W39693));
  NANDX1 G23844 (.A1(W38297), .A2(W18872), .ZN(W39691));
  NANDX1 G23845 (.A1(W25355), .A2(W1380), .ZN(O10381));
  NANDX1 G23846 (.A1(W30055), .A2(W10092), .ZN(W39686));
  NANDX1 G23847 (.A1(W19049), .A2(W37027), .ZN(O10380));
  NANDX1 G23848 (.A1(W16746), .A2(W30945), .ZN(W39680));
  NANDX1 G23849 (.A1(W29756), .A2(W31796), .ZN(W39880));
  NANDX1 G23850 (.A1(W18000), .A2(W27071), .ZN(O10372));
  NANDX1 G23851 (.A1(W35754), .A2(W15603), .ZN(O10370));
  NANDX1 G23852 (.A1(W20501), .A2(W27056), .ZN(W39661));
  NANDX1 G23853 (.A1(W10571), .A2(W9005), .ZN(W39660));
  NANDX1 G23854 (.A1(W13413), .A2(W2855), .ZN(O10363));
  NANDX1 G23855 (.A1(W28836), .A2(W38746), .ZN(O10361));
  NANDX1 G23856 (.A1(W30071), .A2(W32860), .ZN(O10354));
  NANDX1 G23857 (.A1(W21275), .A2(W14198), .ZN(O10349));
  NANDX1 G23858 (.A1(W18123), .A2(W11396), .ZN(W39636));
  NANDX1 G23859 (.A1(W22053), .A2(W9682), .ZN(O10343));
  NANDX1 G23860 (.A1(W16093), .A2(W31587), .ZN(W39625));
  NANDX1 G23861 (.A1(W30187), .A2(W12119), .ZN(O10652));
  NANDX1 G23862 (.A1(W34459), .A2(W25683), .ZN(O10667));
  NANDX1 G23863 (.A1(W4011), .A2(I548), .ZN(O10666));
  NANDX1 G23864 (.A1(W15148), .A2(W8150), .ZN(O10662));
  NANDX1 G23865 (.A1(W31266), .A2(I572), .ZN(O10661));
  NANDX1 G23866 (.A1(W37935), .A2(W755), .ZN(O10660));
  NANDX1 G23867 (.A1(W1617), .A2(W16641), .ZN(O10659));
  NANDX1 G23868 (.A1(W11967), .A2(I1310), .ZN(O10658));
  NANDX1 G23869 (.A1(W29622), .A2(W4143), .ZN(O10657));
  NANDX1 G23870 (.A1(W21914), .A2(W12647), .ZN(O10656));
  NANDX1 G23871 (.A1(W2930), .A2(W21042), .ZN(W40080));
  NANDX1 G23872 (.A1(W24293), .A2(W15869), .ZN(W40079));
  NANDX1 G23873 (.A1(W462), .A2(W11379), .ZN(W40078));
  NANDX1 G23874 (.A1(W10059), .A2(W26513), .ZN(O10674));
  NANDX1 G23875 (.A1(W5035), .A2(W15035), .ZN(O10649));
  NANDX1 G23876 (.A1(W22244), .A2(W438), .ZN(O10647));
  NANDX1 G23877 (.A1(W11531), .A2(W24194), .ZN(O10643));
  NANDX1 G23878 (.A1(W36735), .A2(W23499), .ZN(O10639));
  NANDX1 G23879 (.A1(W32104), .A2(W22471), .ZN(O10636));
  NANDX1 G23880 (.A1(W12913), .A2(W18891), .ZN(O10635));
  NANDX1 G23881 (.A1(W3555), .A2(W28168), .ZN(W40048));
  NANDX1 G23882 (.A1(W2874), .A2(I1768), .ZN(W40047));
  NANDX1 G23883 (.A1(W4181), .A2(W6849), .ZN(W40045));
  NANDX1 G23884 (.A1(W16431), .A2(W8079), .ZN(W40039));
  NANDX1 G23885 (.A1(W12495), .A2(I1621), .ZN(W40032));
  NANDX1 G23886 (.A1(I1161), .A2(W29144), .ZN(W40160));
  NANDX1 G23887 (.A1(W10651), .A2(W29700), .ZN(W40194));
  NANDX1 G23888 (.A1(W1280), .A2(W25903), .ZN(O10732));
  NANDX1 G23889 (.A1(W34447), .A2(W34238), .ZN(O10731));
  NANDX1 G23890 (.A1(W30780), .A2(W29064), .ZN(W40190));
  NANDX1 G23891 (.A1(W3819), .A2(W11924), .ZN(O10729));
  NANDX1 G23892 (.A1(W23130), .A2(W36797), .ZN(O10728));
  NANDX1 G23893 (.A1(W33921), .A2(W19045), .ZN(W40180));
  NANDX1 G23894 (.A1(W33290), .A2(W2172), .ZN(W40179));
  NANDX1 G23895 (.A1(W26416), .A2(W35839), .ZN(W40174));
  NANDX1 G23896 (.A1(W11231), .A2(W11061), .ZN(O10722));
  NANDX1 G23897 (.A1(W12226), .A2(W24517), .ZN(O10721));
  NANDX1 G23898 (.A1(W26112), .A2(W2351), .ZN(W40167));
  NANDX1 G23899 (.A1(W34808), .A2(W23524), .ZN(O10621));
  NANDX1 G23900 (.A1(W17220), .A2(W21959), .ZN(W40158));
  NANDX1 G23901 (.A1(W21342), .A2(W38757), .ZN(O10711));
  NANDX1 G23902 (.A1(W27275), .A2(W10774), .ZN(W40156));
  NANDX1 G23903 (.A1(W36254), .A2(W8151), .ZN(O10707));
  NANDX1 G23904 (.A1(W7347), .A2(W32436), .ZN(W40148));
  NANDX1 G23905 (.A1(W7871), .A2(W31448), .ZN(O10693));
  NANDX1 G23906 (.A1(W29647), .A2(W22424), .ZN(O10692));
  NANDX1 G23907 (.A1(W33146), .A2(W4024), .ZN(O10688));
  NANDX1 G23908 (.A1(W18395), .A2(W3760), .ZN(O10686));
  NANDX1 G23909 (.A1(W34710), .A2(W19658), .ZN(O10685));
  NANDX1 G23910 (.A1(W11388), .A2(W4327), .ZN(O10683));
  NANDX1 G23911 (.A1(W37682), .A2(W7482), .ZN(O10550));
  NANDX1 G23912 (.A1(W857), .A2(W5785), .ZN(O10582));
  NANDX1 G23913 (.A1(W11373), .A2(W1941), .ZN(O10579));
  NANDX1 G23914 (.A1(W35802), .A2(W38757), .ZN(O10576));
  NANDX1 G23915 (.A1(W25169), .A2(W12329), .ZN(O10575));
  NANDX1 G23916 (.A1(W18872), .A2(W12686), .ZN(W39958));
  NANDX1 G23917 (.A1(W26043), .A2(W2810), .ZN(O10572));
  NANDX1 G23918 (.A1(W27894), .A2(W11537), .ZN(O10571));
  NANDX1 G23919 (.A1(W19105), .A2(W36326), .ZN(W39944));
  NANDX1 G23920 (.A1(W422), .A2(W7597), .ZN(O10564));
  NANDX1 G23921 (.A1(W25783), .A2(W34937), .ZN(W39936));
  NANDX1 G23922 (.A1(W22834), .A2(W36237), .ZN(O10558));
  NANDX1 G23923 (.A1(W29140), .A2(W26445), .ZN(O10553));
  NANDX1 G23924 (.A1(W34264), .A2(W14455), .ZN(W39971));
  NANDX1 G23925 (.A1(W37579), .A2(W23726), .ZN(W39921));
  NANDX1 G23926 (.A1(W16961), .A2(W17788), .ZN(O10542));
  NANDX1 G23927 (.A1(W18167), .A2(W2197), .ZN(O10540));
  NANDX1 G23928 (.A1(W355), .A2(W6505), .ZN(O10539));
  NANDX1 G23929 (.A1(W11334), .A2(W7128), .ZN(O10531));
  NANDX1 G23930 (.A1(W28698), .A2(W125), .ZN(O10530));
  NANDX1 G23931 (.A1(W12649), .A2(W23098), .ZN(W39895));
  NANDX1 G23932 (.A1(W18700), .A2(W38072), .ZN(O10529));
  NANDX1 G23933 (.A1(I608), .A2(W9214), .ZN(W39893));
  NANDX1 G23934 (.A1(W27553), .A2(W35043), .ZN(O10528));
  NANDX1 G23935 (.A1(W37217), .A2(W5946), .ZN(O10522));
  NANDX1 G23936 (.A1(W26100), .A2(W23583), .ZN(O10600));
  NANDX1 G23937 (.A1(W28687), .A2(W8916), .ZN(O10619));
  NANDX1 G23938 (.A1(W17106), .A2(W29739), .ZN(W40026));
  NANDX1 G23939 (.A1(W5319), .A2(W918), .ZN(O10613));
  NANDX1 G23940 (.A1(W39432), .A2(W39788), .ZN(O10611));
  NANDX1 G23941 (.A1(W32095), .A2(W3363), .ZN(W40009));
  NANDX1 G23942 (.A1(W20914), .A2(W39196), .ZN(W40008));
  NANDX1 G23943 (.A1(W13414), .A2(W23557), .ZN(O10606));
  NANDX1 G23944 (.A1(W11955), .A2(W6502), .ZN(O10604));
  NANDX1 G23945 (.A1(W35209), .A2(I126), .ZN(O10602));
  NANDX1 G23946 (.A1(W30835), .A2(W32661), .ZN(W40000));
  NANDX1 G23947 (.A1(W34049), .A2(I714), .ZN(O10601));
  NANDX1 G23948 (.A1(W20746), .A2(W5216), .ZN(O10293));
  NANDX1 G23949 (.A1(W12572), .A2(W31500), .ZN(O10598));
  NANDX1 G23950 (.A1(W2303), .A2(W8358), .ZN(O10597));
  NANDX1 G23951 (.A1(W1184), .A2(I557), .ZN(O10595));
  NANDX1 G23952 (.A1(W8478), .A2(W26970), .ZN(O10594));
  NANDX1 G23953 (.A1(W12183), .A2(W13499), .ZN(O10593));
  NANDX1 G23954 (.A1(I1401), .A2(W6132), .ZN(W39988));
  NANDX1 G23955 (.A1(W39550), .A2(W2522), .ZN(W39978));
  NANDX1 G23956 (.A1(W27572), .A2(W12844), .ZN(O10584));
  NANDX1 G23957 (.A1(W14564), .A2(W1564), .ZN(W39974));
  NANDX1 G23958 (.A1(W31387), .A2(W9179), .ZN(W39973));
  NANDX1 G23959 (.A1(W13740), .A2(W19219), .ZN(O10583));
  NANDX1 G23960 (.A1(W27108), .A2(W25421), .ZN(O9990));
  NANDX1 G23961 (.A1(W31768), .A2(W31463), .ZN(O10008));
  NANDX1 G23962 (.A1(W7819), .A2(W26198), .ZN(O10007));
  NANDX1 G23963 (.A1(W15684), .A2(W25177), .ZN(O10005));
  NANDX1 G23964 (.A1(W35260), .A2(W29875), .ZN(O10004));
  NANDX1 G23965 (.A1(I1558), .A2(W2879), .ZN(O10002));
  NANDX1 G23966 (.A1(W15419), .A2(W24281), .ZN(O10001));
  NANDX1 G23967 (.A1(W3593), .A2(W19623), .ZN(W39138));
  NANDX1 G23968 (.A1(W27910), .A2(W22871), .ZN(W39137));
  NANDX1 G23969 (.A1(W32960), .A2(W6794), .ZN(O9998));
  NANDX1 G23970 (.A1(W9240), .A2(W4444), .ZN(O9996));
  NANDX1 G23971 (.A1(W4930), .A2(W25621), .ZN(W39129));
  NANDX1 G23972 (.A1(W2017), .A2(W7979), .ZN(O9991));
  NANDX1 G23973 (.A1(W18640), .A2(W31730), .ZN(W39154));
  NANDX1 G23974 (.A1(W7421), .A2(W33834), .ZN(O9989));
  NANDX1 G23975 (.A1(W11046), .A2(W20148), .ZN(O9986));
  NANDX1 G23976 (.A1(W8759), .A2(W27829), .ZN(O9983));
  NANDX1 G23977 (.A1(W3530), .A2(W20563), .ZN(W39114));
  NANDX1 G23978 (.A1(W23446), .A2(W24139), .ZN(O9974));
  NANDX1 G23979 (.A1(I760), .A2(W6207), .ZN(W39101));
  NANDX1 G23980 (.A1(W27242), .A2(W26461), .ZN(O9972));
  NANDX1 G23981 (.A1(W14086), .A2(W37200), .ZN(W39099));
  NANDX1 G23982 (.A1(W6585), .A2(W4510), .ZN(W39098));
  NANDX1 G23983 (.A1(W10565), .A2(W17451), .ZN(O9969));
  NANDX1 G23984 (.A1(W31404), .A2(W18761), .ZN(O9968));
  NANDX1 G23985 (.A1(W34388), .A2(W29682), .ZN(W39193));
  NANDX1 G23986 (.A1(W550), .A2(W22372), .ZN(O10064));
  NANDX1 G23987 (.A1(W21742), .A2(W38672), .ZN(O10063));
  NANDX1 G23988 (.A1(W18325), .A2(W37395), .ZN(O10059));
  NANDX1 G23989 (.A1(W32751), .A2(W19342), .ZN(O10057));
  NANDX1 G23990 (.A1(W20881), .A2(W14779), .ZN(W39216));
  NANDX1 G23991 (.A1(W2084), .A2(W10146), .ZN(O10056));
  NANDX1 G23992 (.A1(W28453), .A2(W32695), .ZN(W39208));
  NANDX1 G23993 (.A1(W29230), .A2(W32543), .ZN(O10048));
  NANDX1 G23994 (.A1(W8975), .A2(W33581), .ZN(W39202));
  NANDX1 G23995 (.A1(W11361), .A2(W3750), .ZN(W39196));
  NANDX1 G23996 (.A1(W10421), .A2(W24389), .ZN(O10042));
  NANDX1 G23997 (.A1(W7579), .A2(W22254), .ZN(O10041));
  NANDX1 G23998 (.A1(W32811), .A2(W10408), .ZN(W39089));
  NANDX1 G23999 (.A1(W32473), .A2(W19259), .ZN(W39181));
  NANDX1 G24000 (.A1(W23934), .A2(W35352), .ZN(O10033));
  NANDX1 G24001 (.A1(W13932), .A2(W13765), .ZN(O10030));
  NANDX1 G24002 (.A1(W1424), .A2(W30067), .ZN(W39176));
  NANDX1 G24003 (.A1(W10568), .A2(W34797), .ZN(O10026));
  NANDX1 G24004 (.A1(W26132), .A2(W23594), .ZN(W39171));
  NANDX1 G24005 (.A1(W38349), .A2(W21631), .ZN(O10024));
  NANDX1 G24006 (.A1(W31330), .A2(I499), .ZN(O10023));
  NANDX1 G24007 (.A1(W18054), .A2(W23843), .ZN(O10019));
  NANDX1 G24008 (.A1(W12447), .A2(W7790), .ZN(O10016));
  NANDX1 G24009 (.A1(W6726), .A2(W3044), .ZN(O10015));
  NANDX1 G24010 (.A1(W8071), .A2(W18597), .ZN(W38979));
  NANDX1 G24011 (.A1(W26662), .A2(W30025), .ZN(W39025));
  NANDX1 G24012 (.A1(W18890), .A2(W33644), .ZN(W39024));
  NANDX1 G24013 (.A1(W4949), .A2(W35677), .ZN(W39021));
  NANDX1 G24014 (.A1(W32512), .A2(I957), .ZN(O9923));
  NANDX1 G24015 (.A1(W30320), .A2(W9659), .ZN(W39015));
  NANDX1 G24016 (.A1(W37745), .A2(W6241), .ZN(W39013));
  NANDX1 G24017 (.A1(W36255), .A2(W35356), .ZN(O9920));
  NANDX1 G24018 (.A1(W4735), .A2(W32505), .ZN(W39009));
  NANDX1 G24019 (.A1(W4199), .A2(W2473), .ZN(O9918));
  NANDX1 G24020 (.A1(W23913), .A2(W22164), .ZN(W38995));
  NANDX1 G24021 (.A1(W6350), .A2(W8266), .ZN(W38992));
  NANDX1 G24022 (.A1(W610), .A2(W12876), .ZN(W38982));
  NANDX1 G24023 (.A1(W13948), .A2(W11584), .ZN(O9928));
  NANDX1 G24024 (.A1(W32864), .A2(W28633), .ZN(O9901));
  NANDX1 G24025 (.A1(W5357), .A2(W16715), .ZN(O9900));
  NANDX1 G24026 (.A1(W25319), .A2(W12016), .ZN(O9897));
  NANDX1 G24027 (.A1(W18797), .A2(W23706), .ZN(O9896));
  NANDX1 G24028 (.A1(W27243), .A2(W8452), .ZN(W38962));
  NANDX1 G24029 (.A1(W8578), .A2(W24842), .ZN(O9888));
  NANDX1 G24030 (.A1(W25207), .A2(W32493), .ZN(O9887));
  NANDX1 G24031 (.A1(W6066), .A2(W1648), .ZN(W38952));
  NANDX1 G24032 (.A1(W18788), .A2(W2643), .ZN(W38951));
  NANDX1 G24033 (.A1(W10256), .A2(W14646), .ZN(O9886));
  NANDX1 G24034 (.A1(W36125), .A2(W18268), .ZN(O9881));
  NANDX1 G24035 (.A1(W31283), .A2(W5220), .ZN(W39065));
  NANDX1 G24036 (.A1(W18920), .A2(W31328), .ZN(W39088));
  NANDX1 G24037 (.A1(W13054), .A2(W28712), .ZN(O9965));
  NANDX1 G24038 (.A1(W33026), .A2(W7630), .ZN(W39086));
  NANDX1 G24039 (.A1(W17142), .A2(W20744), .ZN(O9964));
  NANDX1 G24040 (.A1(W21264), .A2(W5123), .ZN(O9962));
  NANDX1 G24041 (.A1(W12283), .A2(W7087), .ZN(O9960));
  NANDX1 G24042 (.A1(W21824), .A2(W8264), .ZN(O9958));
  NANDX1 G24043 (.A1(W16032), .A2(W14044), .ZN(O9954));
  NANDX1 G24044 (.A1(W6118), .A2(W3393), .ZN(O9953));
  NANDX1 G24045 (.A1(W13795), .A2(W26946), .ZN(O9952));
  NANDX1 G24046 (.A1(W3862), .A2(W16433), .ZN(O9951));
  NANDX1 G24047 (.A1(W24780), .A2(W24696), .ZN(O10065));
  NANDX1 G24048 (.A1(W25845), .A2(W16126), .ZN(W39059));
  NANDX1 G24049 (.A1(W29873), .A2(W23211), .ZN(O9944));
  NANDX1 G24050 (.A1(W7559), .A2(W23011), .ZN(W39055));
  NANDX1 G24051 (.A1(I357), .A2(W30490), .ZN(O9940));
  NANDX1 G24052 (.A1(W38162), .A2(W36982), .ZN(W39050));
  NANDX1 G24053 (.A1(W10997), .A2(W26418), .ZN(O9939));
  NANDX1 G24054 (.A1(W38062), .A2(W18380), .ZN(O9937));
  NANDX1 G24055 (.A1(W33406), .A2(W30114), .ZN(O9936));
  NANDX1 G24056 (.A1(W24868), .A2(W14666), .ZN(W39042));
  NANDX1 G24057 (.A1(W10624), .A2(W24585), .ZN(O9932));
  NANDX1 G24058 (.A1(W29211), .A2(W30436), .ZN(W39034));
  NANDX1 G24059 (.A1(I852), .A2(W20759), .ZN(O10195));
  NANDX1 G24060 (.A1(W2525), .A2(W36337), .ZN(O10236));
  NANDX1 G24061 (.A1(W30353), .A2(W37036), .ZN(O10235));
  NANDX1 G24062 (.A1(W36325), .A2(W32826), .ZN(O10232));
  NANDX1 G24063 (.A1(W7094), .A2(W4801), .ZN(O10229));
  NANDX1 G24064 (.A1(W2044), .A2(W36859), .ZN(O10228));
  NANDX1 G24065 (.A1(W26209), .A2(W12824), .ZN(W39465));
  NANDX1 G24066 (.A1(W34084), .A2(W33466), .ZN(W39459));
  NANDX1 G24067 (.A1(W20323), .A2(W6077), .ZN(O10222));
  NANDX1 G24068 (.A1(W24429), .A2(W33761), .ZN(O10211));
  NANDX1 G24069 (.A1(W9683), .A2(W1331), .ZN(O10208));
  NANDX1 G24070 (.A1(W25977), .A2(W35369), .ZN(O10206));
  NANDX1 G24071 (.A1(W12879), .A2(W27223), .ZN(W39432));
  NANDX1 G24072 (.A1(W31636), .A2(W21945), .ZN(W39479));
  NANDX1 G24073 (.A1(W34891), .A2(W4881), .ZN(W39415));
  NANDX1 G24074 (.A1(W38915), .A2(W34583), .ZN(O10192));
  NANDX1 G24075 (.A1(I731), .A2(W34797), .ZN(O10190));
  NANDX1 G24076 (.A1(W31255), .A2(W32392), .ZN(O10188));
  NANDX1 G24077 (.A1(W32046), .A2(W35982), .ZN(W39406));
  NANDX1 G24078 (.A1(W14179), .A2(W3081), .ZN(W39403));
  NANDX1 G24079 (.A1(W38491), .A2(W26675), .ZN(O10176));
  NANDX1 G24080 (.A1(W2092), .A2(W30766), .ZN(O10172));
  NANDX1 G24081 (.A1(W4119), .A2(W14234), .ZN(W39379));
  NANDX1 G24082 (.A1(W25304), .A2(W26690), .ZN(O10165));
  NANDX1 G24083 (.A1(W276), .A2(W19624), .ZN(O10161));
  NANDX1 G24084 (.A1(W36403), .A2(W20), .ZN(O10262));
  NANDX1 G24085 (.A1(W27095), .A2(W865), .ZN(O10292));
  NANDX1 G24086 (.A1(W22839), .A2(W37590), .ZN(W39555));
  NANDX1 G24087 (.A1(W37308), .A2(W3665), .ZN(O10289));
  NANDX1 G24088 (.A1(W38141), .A2(W37457), .ZN(W39550));
  NANDX1 G24089 (.A1(W1937), .A2(W20576), .ZN(O10285));
  NANDX1 G24090 (.A1(W5187), .A2(W18590), .ZN(W39547));
  NANDX1 G24091 (.A1(W36796), .A2(W32925), .ZN(O10281));
  NANDX1 G24092 (.A1(W26702), .A2(W21871), .ZN(O10278));
  NANDX1 G24093 (.A1(W3536), .A2(W23054), .ZN(O10277));
  NANDX1 G24094 (.A1(W25463), .A2(W788), .ZN(O10274));
  NANDX1 G24095 (.A1(W32155), .A2(W31944), .ZN(W39528));
  NANDX1 G24096 (.A1(W14299), .A2(W37165), .ZN(O10263));
  NANDX1 G24097 (.A1(W16661), .A2(W5704), .ZN(O10160));
  NANDX1 G24098 (.A1(W1619), .A2(W20861), .ZN(W39514));
  NANDX1 G24099 (.A1(W25330), .A2(W26655), .ZN(O10260));
  NANDX1 G24100 (.A1(W6699), .A2(W104), .ZN(O10258));
  NANDX1 G24101 (.A1(W10178), .A2(W26095), .ZN(W39505));
  NANDX1 G24102 (.A1(W26875), .A2(W17671), .ZN(O10250));
  NANDX1 G24103 (.A1(W10779), .A2(W35251), .ZN(W39491));
  NANDX1 G24104 (.A1(W28871), .A2(W39261), .ZN(O10241));
  NANDX1 G24105 (.A1(W34548), .A2(W5986), .ZN(W39484));
  NANDX1 G24106 (.A1(W4849), .A2(W25096), .ZN(O10240));
  NANDX1 G24107 (.A1(W8549), .A2(W543), .ZN(O10239));
  NANDX1 G24108 (.A1(I171), .A2(W15998), .ZN(O10238));
  NANDX1 G24109 (.A1(W28815), .A2(W2612), .ZN(W39257));
  NANDX1 G24110 (.A1(W29217), .A2(W38361), .ZN(W39289));
  NANDX1 G24111 (.A1(W35793), .A2(W36599), .ZN(W39288));
  NANDX1 G24112 (.A1(W34958), .A2(W18691), .ZN(O10102));
  NANDX1 G24113 (.A1(W23692), .A2(W30679), .ZN(O10100));
  NANDX1 G24114 (.A1(W33244), .A2(W29001), .ZN(O10099));
  NANDX1 G24115 (.A1(W878), .A2(W4713), .ZN(O10096));
  NANDX1 G24116 (.A1(W1741), .A2(W145), .ZN(O10095));
  NANDX1 G24117 (.A1(W10435), .A2(W6755), .ZN(O10094));
  NANDX1 G24118 (.A1(W25241), .A2(W5546), .ZN(W39267));
  NANDX1 G24119 (.A1(W10677), .A2(W9395), .ZN(W39264));
  NANDX1 G24120 (.A1(W13499), .A2(W30), .ZN(O10088));
  NANDX1 G24121 (.A1(W20751), .A2(I1738), .ZN(W39260));
  NANDX1 G24122 (.A1(W34921), .A2(W2005), .ZN(O10106));
  NANDX1 G24123 (.A1(W4410), .A2(W7287), .ZN(W39256));
  NANDX1 G24124 (.A1(W18792), .A2(W5945), .ZN(O10085));
  NANDX1 G24125 (.A1(W12771), .A2(W14089), .ZN(O10081));
  NANDX1 G24126 (.A1(W4886), .A2(W38354), .ZN(O10080));
  NANDX1 G24127 (.A1(W32453), .A2(W12351), .ZN(O10077));
  NANDX1 G24128 (.A1(W30767), .A2(W31303), .ZN(W39242));
  NANDX1 G24129 (.A1(W29278), .A2(W21797), .ZN(W39241));
  NANDX1 G24130 (.A1(W27177), .A2(W38916), .ZN(O10071));
  NANDX1 G24131 (.A1(W22516), .A2(W11342), .ZN(W39235));
  NANDX1 G24132 (.A1(W26499), .A2(W26662), .ZN(W39233));
  NANDX1 G24133 (.A1(W27302), .A2(W11589), .ZN(O10069));
  NANDX1 G24134 (.A1(W12656), .A2(W25003), .ZN(O10135));
  NANDX1 G24135 (.A1(W34004), .A2(W28440), .ZN(O10152));
  NANDX1 G24136 (.A1(W376), .A2(W4483), .ZN(O10148));
  NANDX1 G24137 (.A1(W38479), .A2(W36809), .ZN(O10147));
  NANDX1 G24138 (.A1(W20694), .A2(W4381), .ZN(O10145));
  NANDX1 G24139 (.A1(W30360), .A2(W16736), .ZN(W39354));
  NANDX1 G24140 (.A1(W33086), .A2(W24605), .ZN(W39352));
  NANDX1 G24141 (.A1(W26763), .A2(W29730), .ZN(O10144));
  NANDX1 G24142 (.A1(W13987), .A2(W14400), .ZN(O10140));
  NANDX1 G24143 (.A1(W11996), .A2(W9475), .ZN(W39344));
  NANDX1 G24144 (.A1(W28368), .A2(W25755), .ZN(O10139));
  NANDX1 G24145 (.A1(W24974), .A2(I1688), .ZN(W39341));
  NANDX1 G24146 (.A1(W32901), .A2(W20836), .ZN(O10733));
  NANDX1 G24147 (.A1(I1639), .A2(W23194), .ZN(O10130));
  NANDX1 G24148 (.A1(W10980), .A2(W3082), .ZN(O10128));
  NANDX1 G24149 (.A1(W25537), .A2(W33821), .ZN(W39328));
  NANDX1 G24150 (.A1(W36237), .A2(W24362), .ZN(O10120));
  NANDX1 G24151 (.A1(W11435), .A2(W32980), .ZN(O10117));
  NANDX1 G24152 (.A1(W7609), .A2(W11781), .ZN(O10116));
  NANDX1 G24153 (.A1(W27457), .A2(W5041), .ZN(O10114));
  NANDX1 G24154 (.A1(W23453), .A2(W2499), .ZN(W39304));
  NANDX1 G24155 (.A1(W28180), .A2(W38090), .ZN(O10111));
  NANDX1 G24156 (.A1(W36608), .A2(W35219), .ZN(O10108));
  NANDX1 G24157 (.A1(W38989), .A2(W7726), .ZN(O10107));
  NANDX1 G24158 (.A1(W39397), .A2(W3338), .ZN(O11333));
  NANDX1 G24159 (.A1(W9127), .A2(W15210), .ZN(O11389));
  NANDX1 G24160 (.A1(W6543), .A2(W7106), .ZN(W41128));
  NANDX1 G24161 (.A1(W5116), .A2(W23256), .ZN(O11384));
  NANDX1 G24162 (.A1(W11154), .A2(W9004), .ZN(O11380));
  NANDX1 G24163 (.A1(W28539), .A2(W11962), .ZN(O11376));
  NANDX1 G24164 (.A1(W10360), .A2(W35852), .ZN(O11366));
  NANDX1 G24165 (.A1(W3232), .A2(W23425), .ZN(O11347));
  NANDX1 G24166 (.A1(W33551), .A2(W36386), .ZN(W41071));
  NANDX1 G24167 (.A1(W27394), .A2(W24851), .ZN(O11343));
  NANDX1 G24168 (.A1(W13906), .A2(W23292), .ZN(O11338));
  NANDX1 G24169 (.A1(W23633), .A2(W16208), .ZN(O11336));
  NANDX1 G24170 (.A1(W26295), .A2(W7991), .ZN(O11334));
  NANDX1 G24171 (.A1(W33221), .A2(W28707), .ZN(O11390));
  NANDX1 G24172 (.A1(W35982), .A2(W23908), .ZN(O11329));
  NANDX1 G24173 (.A1(I163), .A2(W15182), .ZN(O11326));
  NANDX1 G24174 (.A1(W20974), .A2(W35706), .ZN(O11325));
  NANDX1 G24175 (.A1(W40202), .A2(W22931), .ZN(O11324));
  NANDX1 G24176 (.A1(W4671), .A2(W30592), .ZN(O11323));
  NANDX1 G24177 (.A1(W28622), .A2(W19791), .ZN(O11322));
  NANDX1 G24178 (.A1(W21090), .A2(W23720), .ZN(O11321));
  NANDX1 G24179 (.A1(W22293), .A2(W34142), .ZN(W41035));
  NANDX1 G24180 (.A1(W32250), .A2(W34865), .ZN(O11316));
  NANDX1 G24181 (.A1(W4106), .A2(W20953), .ZN(W41031));
  NANDX1 G24182 (.A1(W27510), .A2(W33870), .ZN(O11314));
  NANDX1 G24183 (.A1(W22933), .A2(W2915), .ZN(O11427));
  NANDX1 G24184 (.A1(W6932), .A2(W11926), .ZN(O11450));
  NANDX1 G24185 (.A1(W23441), .A2(W9504), .ZN(O11447));
  NANDX1 G24186 (.A1(W37778), .A2(W39877), .ZN(O11445));
  NANDX1 G24187 (.A1(W33149), .A2(W6754), .ZN(O11441));
  NANDX1 G24188 (.A1(W13244), .A2(W33518), .ZN(O11440));
  NANDX1 G24189 (.A1(W3951), .A2(I22), .ZN(O11439));
  NANDX1 G24190 (.A1(W63), .A2(W5988), .ZN(O11437));
  NANDX1 G24191 (.A1(W35862), .A2(W11143), .ZN(W41198));
  NANDX1 G24192 (.A1(W27575), .A2(I960), .ZN(O11434));
  NANDX1 G24193 (.A1(W29045), .A2(W36999), .ZN(O11433));
  NANDX1 G24194 (.A1(W2161), .A2(W3703), .ZN(O11430));
  NANDX1 G24195 (.A1(W18933), .A2(W37522), .ZN(O11428));
  NANDX1 G24196 (.A1(W21484), .A2(W29003), .ZN(O11311));
  NANDX1 G24197 (.A1(W37787), .A2(W36239), .ZN(O11425));
  NANDX1 G24198 (.A1(W38287), .A2(W15218), .ZN(W41176));
  NANDX1 G24199 (.A1(W5093), .A2(W26385), .ZN(O11424));
  NANDX1 G24200 (.A1(W25108), .A2(W4381), .ZN(O11423));
  NANDX1 G24201 (.A1(W30346), .A2(W23625), .ZN(W41173));
  NANDX1 G24202 (.A1(W40999), .A2(W6910), .ZN(O11418));
  NANDX1 G24203 (.A1(W13257), .A2(W19989), .ZN(W41165));
  NANDX1 G24204 (.A1(W12170), .A2(W593), .ZN(O11417));
  NANDX1 G24205 (.A1(W18079), .A2(W15700), .ZN(O11413));
  NANDX1 G24206 (.A1(W8525), .A2(W9489), .ZN(O11410));
  NANDX1 G24207 (.A1(W8017), .A2(W21323), .ZN(W41142));
  NANDX1 G24208 (.A1(W35638), .A2(W17327), .ZN(O11225));
  NANDX1 G24209 (.A1(W22981), .A2(W37126), .ZN(O11249));
  NANDX1 G24210 (.A1(W30689), .A2(W26702), .ZN(W40927));
  NANDX1 G24211 (.A1(W12369), .A2(W18605), .ZN(O11245));
  NANDX1 G24212 (.A1(W17496), .A2(W11915), .ZN(O11240));
  NANDX1 G24213 (.A1(W7246), .A2(W39686), .ZN(O11239));
  NANDX1 G24214 (.A1(W38345), .A2(W18889), .ZN(O11237));
  NANDX1 G24215 (.A1(W3386), .A2(W16099), .ZN(W40911));
  NANDX1 G24216 (.A1(W3214), .A2(W22314), .ZN(O11233));
  NANDX1 G24217 (.A1(W35387), .A2(W6092), .ZN(O11231));
  NANDX1 G24218 (.A1(W12830), .A2(W36031), .ZN(O11230));
  NANDX1 G24219 (.A1(W14399), .A2(W37447), .ZN(W40905));
  NANDX1 G24220 (.A1(W12731), .A2(W17147), .ZN(W40904));
  NANDX1 G24221 (.A1(W19020), .A2(W36175), .ZN(O11252));
  NANDX1 G24222 (.A1(W681), .A2(W13742), .ZN(O11222));
  NANDX1 G24223 (.A1(W33623), .A2(W32034), .ZN(O11217));
  NANDX1 G24224 (.A1(I921), .A2(W38180), .ZN(W40889));
  NANDX1 G24225 (.A1(W12505), .A2(W37055), .ZN(W40885));
  NANDX1 G24226 (.A1(W24996), .A2(W9814), .ZN(O11214));
  NANDX1 G24227 (.A1(W12498), .A2(W35551), .ZN(O11209));
  NANDX1 G24228 (.A1(W23293), .A2(W14878), .ZN(O11207));
  NANDX1 G24229 (.A1(W37096), .A2(W1860), .ZN(W40866));
  NANDX1 G24230 (.A1(W25724), .A2(W7421), .ZN(O11198));
  NANDX1 G24231 (.A1(W9603), .A2(W38240), .ZN(W40860));
  NANDX1 G24232 (.A1(W32864), .A2(W17899), .ZN(W40848));
  NANDX1 G24233 (.A1(W900), .A2(W17079), .ZN(W40992));
  NANDX1 G24234 (.A1(W35354), .A2(W33492), .ZN(W41018));
  NANDX1 G24235 (.A1(W26020), .A2(W26337), .ZN(O11307));
  NANDX1 G24236 (.A1(W28563), .A2(W22509), .ZN(O11305));
  NANDX1 G24237 (.A1(W15390), .A2(W27512), .ZN(W41009));
  NANDX1 G24238 (.A1(W35899), .A2(W3327), .ZN(O11302));
  NANDX1 G24239 (.A1(W795), .A2(I1535), .ZN(O11301));
  NANDX1 G24240 (.A1(W33036), .A2(W27400), .ZN(O11300));
  NANDX1 G24241 (.A1(W14272), .A2(W2792), .ZN(W41002));
  NANDX1 G24242 (.A1(I430), .A2(W40148), .ZN(O11299));
  NANDX1 G24243 (.A1(W26716), .A2(W21081), .ZN(O11296));
  NANDX1 G24244 (.A1(W5383), .A2(W5712), .ZN(O11295));
  NANDX1 G24245 (.A1(W39974), .A2(W19876), .ZN(O11451));
  NANDX1 G24246 (.A1(W30782), .A2(I687), .ZN(W40986));
  NANDX1 G24247 (.A1(W26894), .A2(W3398), .ZN(O11290));
  NANDX1 G24248 (.A1(W22959), .A2(I1381), .ZN(O11282));
  NANDX1 G24249 (.A1(W5255), .A2(W6347), .ZN(W40970));
  NANDX1 G24250 (.A1(I1932), .A2(W17011), .ZN(O11273));
  NANDX1 G24251 (.A1(W33312), .A2(W28687), .ZN(O11267));
  NANDX1 G24252 (.A1(W39465), .A2(W37109), .ZN(W40952));
  NANDX1 G24253 (.A1(W16243), .A2(I1556), .ZN(W40951));
  NANDX1 G24254 (.A1(W33499), .A2(W36168), .ZN(W40945));
  NANDX1 G24255 (.A1(W1385), .A2(W36267), .ZN(O11255));
  NANDX1 G24256 (.A1(W31899), .A2(W17319), .ZN(O11254));
  NANDX1 G24257 (.A1(W19649), .A2(W36351), .ZN(O11585));
  NANDX1 G24258 (.A1(W24930), .A2(W23438), .ZN(O11602));
  NANDX1 G24259 (.A1(W41209), .A2(W9284), .ZN(O11600));
  NANDX1 G24260 (.A1(W7841), .A2(W19598), .ZN(O11599));
  NANDX1 G24261 (.A1(W9469), .A2(W2056), .ZN(O11597));
  NANDX1 G24262 (.A1(W22544), .A2(W8614), .ZN(O11595));
  NANDX1 G24263 (.A1(W28755), .A2(W550), .ZN(O11594));
  NANDX1 G24264 (.A1(W24220), .A2(W22193), .ZN(O11593));
  NANDX1 G24265 (.A1(W28662), .A2(W21289), .ZN(O11592));
  NANDX1 G24266 (.A1(W7799), .A2(W6143), .ZN(O11590));
  NANDX1 G24267 (.A1(W3553), .A2(W28087), .ZN(O11588));
  NANDX1 G24268 (.A1(W15210), .A2(W10787), .ZN(O11587));
  NANDX1 G24269 (.A1(W13467), .A2(W34561), .ZN(O11586));
  NANDX1 G24270 (.A1(W24025), .A2(W24374), .ZN(O11603));
  NANDX1 G24271 (.A1(W15141), .A2(W18164), .ZN(O11584));
  NANDX1 G24272 (.A1(W11414), .A2(W31227), .ZN(W41410));
  NANDX1 G24273 (.A1(W15852), .A2(W21863), .ZN(O11577));
  NANDX1 G24274 (.A1(W38566), .A2(W29682), .ZN(O11576));
  NANDX1 G24275 (.A1(W16270), .A2(W34693), .ZN(W41403));
  NANDX1 G24276 (.A1(W38963), .A2(W3551), .ZN(W41400));
  NANDX1 G24277 (.A1(W35662), .A2(W23106), .ZN(W41397));
  NANDX1 G24278 (.A1(W11781), .A2(W30899), .ZN(O11569));
  NANDX1 G24279 (.A1(W2924), .A2(W13332), .ZN(W41393));
  NANDX1 G24280 (.A1(W21994), .A2(W13585), .ZN(O11565));
  NANDX1 G24281 (.A1(W6814), .A2(W5789), .ZN(O11564));
  NANDX1 G24282 (.A1(W23491), .A2(W6185), .ZN(O11630));
  NANDX1 G24283 (.A1(W35782), .A2(W21319), .ZN(W41523));
  NANDX1 G24284 (.A1(W20648), .A2(W28973), .ZN(O11662));
  NANDX1 G24285 (.A1(W10240), .A2(W38029), .ZN(O11661));
  NANDX1 G24286 (.A1(W25847), .A2(W1331), .ZN(O11658));
  NANDX1 G24287 (.A1(W32283), .A2(I1264), .ZN(W41512));
  NANDX1 G24288 (.A1(W21180), .A2(W3417), .ZN(O11652));
  NANDX1 G24289 (.A1(W16513), .A2(W27960), .ZN(W41497));
  NANDX1 G24290 (.A1(W9219), .A2(W39849), .ZN(O11642));
  NANDX1 G24291 (.A1(W987), .A2(W429), .ZN(O11639));
  NANDX1 G24292 (.A1(W31466), .A2(I1579), .ZN(O11634));
  NANDX1 G24293 (.A1(W27267), .A2(W27083), .ZN(O11632));
  NANDX1 G24294 (.A1(W41281), .A2(W37713), .ZN(O11631));
  NANDX1 G24295 (.A1(W24300), .A2(W16585), .ZN(W41387));
  NANDX1 G24296 (.A1(W27661), .A2(W32949), .ZN(W41475));
  NANDX1 G24297 (.A1(W41465), .A2(W21580), .ZN(W41473));
  NANDX1 G24298 (.A1(W20858), .A2(W16065), .ZN(W41469));
  NANDX1 G24299 (.A1(W30379), .A2(I1614), .ZN(O11622));
  NANDX1 G24300 (.A1(W7752), .A2(I1602), .ZN(W41463));
  NANDX1 G24301 (.A1(W32097), .A2(W3496), .ZN(O11617));
  NANDX1 G24302 (.A1(W14374), .A2(W10897), .ZN(W41454));
  NANDX1 G24303 (.A1(W26669), .A2(W15181), .ZN(W41453));
  NANDX1 G24304 (.A1(W5682), .A2(W38435), .ZN(O11609));
  NANDX1 G24305 (.A1(W35477), .A2(W16011), .ZN(O11608));
  NANDX1 G24306 (.A1(W17777), .A2(W27756), .ZN(O11607));
  NANDX1 G24307 (.A1(W35059), .A2(I1352), .ZN(W41265));
  NANDX1 G24308 (.A1(I1837), .A2(W6135), .ZN(O11510));
  NANDX1 G24309 (.A1(W5413), .A2(W32224), .ZN(O11502));
  NANDX1 G24310 (.A1(W24640), .A2(W28271), .ZN(O11499));
  NANDX1 G24311 (.A1(W31486), .A2(W12870), .ZN(O11498));
  NANDX1 G24312 (.A1(W6488), .A2(W2307), .ZN(W41298));
  NANDX1 G24313 (.A1(W22973), .A2(W24481), .ZN(O11493));
  NANDX1 G24314 (.A1(W37982), .A2(W32051), .ZN(O11492));
  NANDX1 G24315 (.A1(I638), .A2(W14068), .ZN(O11491));
  NANDX1 G24316 (.A1(W4421), .A2(W10898), .ZN(W41282));
  NANDX1 G24317 (.A1(W24652), .A2(W19122), .ZN(W41276));
  NANDX1 G24318 (.A1(W26894), .A2(W34170), .ZN(W41270));
  NANDX1 G24319 (.A1(W32722), .A2(W13531), .ZN(O11481));
  NANDX1 G24320 (.A1(W39655), .A2(I885), .ZN(O11511));
  NANDX1 G24321 (.A1(W1313), .A2(W5302), .ZN(O11476));
  NANDX1 G24322 (.A1(W26183), .A2(I522), .ZN(O11472));
  NANDX1 G24323 (.A1(W31451), .A2(W15414), .ZN(W41252));
  NANDX1 G24324 (.A1(W13289), .A2(W37380), .ZN(O11470));
  NANDX1 G24325 (.A1(W22609), .A2(W7810), .ZN(O11467));
  NANDX1 G24326 (.A1(W30803), .A2(W40860), .ZN(W41245));
  NANDX1 G24327 (.A1(W17528), .A2(W19417), .ZN(O11463));
  NANDX1 G24328 (.A1(W40364), .A2(W4846), .ZN(W41236));
  NANDX1 G24329 (.A1(W28471), .A2(W23041), .ZN(W41234));
  NANDX1 G24330 (.A1(W366), .A2(I485), .ZN(W41233));
  NANDX1 G24331 (.A1(W12652), .A2(W1081), .ZN(W41229));
  NANDX1 G24332 (.A1(I1154), .A2(W32919), .ZN(W41342));
  NANDX1 G24333 (.A1(W21136), .A2(W6654), .ZN(O11562));
  NANDX1 G24334 (.A1(W12376), .A2(W29876), .ZN(W41382));
  NANDX1 G24335 (.A1(W22234), .A2(I433), .ZN(W41380));
  NANDX1 G24336 (.A1(W25131), .A2(W13733), .ZN(O11558));
  NANDX1 G24337 (.A1(W2711), .A2(W36233), .ZN(W41374));
  NANDX1 G24338 (.A1(W30071), .A2(W7), .ZN(O11555));
  NANDX1 G24339 (.A1(W19844), .A2(W11938), .ZN(W41363));
  NANDX1 G24340 (.A1(W16033), .A2(W6367), .ZN(O11548));
  NANDX1 G24341 (.A1(W32259), .A2(W34557), .ZN(O11544));
  NANDX1 G24342 (.A1(W25787), .A2(W10738), .ZN(O11537));
  NANDX1 G24343 (.A1(W3369), .A2(W17840), .ZN(O11536));
  NANDX1 G24344 (.A1(W10816), .A2(W4037), .ZN(O11186));
  NANDX1 G24345 (.A1(W17510), .A2(W15639), .ZN(O11530));
  NANDX1 G24346 (.A1(W22700), .A2(W30308), .ZN(O11524));
  NANDX1 G24347 (.A1(W37767), .A2(W38533), .ZN(O11523));
  NANDX1 G24348 (.A1(W29466), .A2(W10920), .ZN(O11522));
  NANDX1 G24349 (.A1(W23803), .A2(W15472), .ZN(O11521));
  NANDX1 G24350 (.A1(W7961), .A2(I628), .ZN(O11520));
  NANDX1 G24351 (.A1(W22613), .A2(W16713), .ZN(O11519));
  NANDX1 G24352 (.A1(W28324), .A2(W13470), .ZN(O11516));
  NANDX1 G24353 (.A1(W5231), .A2(W5423), .ZN(O11515));
  NANDX1 G24354 (.A1(W35580), .A2(W31492), .ZN(O11513));
  NANDX1 G24355 (.A1(W14928), .A2(W18372), .ZN(O11512));
  NANDX1 G24356 (.A1(W36524), .A2(W28931), .ZN(O10852));
  NANDX1 G24357 (.A1(W22575), .A2(W30397), .ZN(O10888));
  NANDX1 G24358 (.A1(W1903), .A2(W33685), .ZN(O10885));
  NANDX1 G24359 (.A1(W25172), .A2(W31234), .ZN(O10882));
  NANDX1 G24360 (.A1(W9399), .A2(W30529), .ZN(O10878));
  NANDX1 G24361 (.A1(W9743), .A2(W28713), .ZN(O10876));
  NANDX1 G24362 (.A1(W19676), .A2(W23713), .ZN(W40412));
  NANDX1 G24363 (.A1(W2782), .A2(W12957), .ZN(O10872));
  NANDX1 G24364 (.A1(W17329), .A2(W36990), .ZN(O10871));
  NANDX1 G24365 (.A1(W11032), .A2(W29844), .ZN(O10862));
  NANDX1 G24366 (.A1(W1080), .A2(W1403), .ZN(O10860));
  NANDX1 G24367 (.A1(W13814), .A2(W17234), .ZN(W40386));
  NANDX1 G24368 (.A1(W36332), .A2(W22651), .ZN(O10855));
  NANDX1 G24369 (.A1(W1446), .A2(W28036), .ZN(O10904));
  NANDX1 G24370 (.A1(W13704), .A2(W796), .ZN(O10851));
  NANDX1 G24371 (.A1(W18500), .A2(W7275), .ZN(W40377));
  NANDX1 G24372 (.A1(W10399), .A2(W38724), .ZN(O10848));
  NANDX1 G24373 (.A1(W1211), .A2(W5772), .ZN(O10847));
  NANDX1 G24374 (.A1(W5283), .A2(W27988), .ZN(W40371));
  NANDX1 G24375 (.A1(W10411), .A2(W25656), .ZN(O10845));
  NANDX1 G24376 (.A1(W13144), .A2(I102), .ZN(O10842));
  NANDX1 G24377 (.A1(W27388), .A2(W30303), .ZN(O10841));
  NANDX1 G24378 (.A1(I267), .A2(W32582), .ZN(O10840));
  NANDX1 G24379 (.A1(W22246), .A2(W1479), .ZN(O10839));
  NANDX1 G24380 (.A1(I863), .A2(W14714), .ZN(O10835));
  NANDX1 G24381 (.A1(W31257), .A2(W15674), .ZN(W40484));
  NANDX1 G24382 (.A1(W13098), .A2(W11755), .ZN(W40519));
  NANDX1 G24383 (.A1(W32383), .A2(W39667), .ZN(O10957));
  NANDX1 G24384 (.A1(W30570), .A2(W36848), .ZN(W40516));
  NANDX1 G24385 (.A1(W11821), .A2(W3422), .ZN(W40514));
  NANDX1 G24386 (.A1(W18832), .A2(W33013), .ZN(W40513));
  NANDX1 G24387 (.A1(W38220), .A2(W4482), .ZN(O10953));
  NANDX1 G24388 (.A1(W14855), .A2(W7763), .ZN(O10952));
  NANDX1 G24389 (.A1(W28659), .A2(W38143), .ZN(O10948));
  NANDX1 G24390 (.A1(W135), .A2(W7085), .ZN(O10945));
  NANDX1 G24391 (.A1(W25975), .A2(W31004), .ZN(O10944));
  NANDX1 G24392 (.A1(W37107), .A2(W38674), .ZN(O10940));
  NANDX1 G24393 (.A1(W35313), .A2(W23261), .ZN(O10939));
  NANDX1 G24394 (.A1(W36440), .A2(W4231), .ZN(O10831));
  NANDX1 G24395 (.A1(W15801), .A2(W14416), .ZN(O10932));
  NANDX1 G24396 (.A1(W2502), .A2(W29117), .ZN(W40479));
  NANDX1 G24397 (.A1(W17337), .A2(W32885), .ZN(W40478));
  NANDX1 G24398 (.A1(W2730), .A2(W15378), .ZN(O10928));
  NANDX1 G24399 (.A1(I947), .A2(W36506), .ZN(O10925));
  NANDX1 G24400 (.A1(I1112), .A2(W28113), .ZN(O10924));
  NANDX1 G24401 (.A1(W4134), .A2(I1639), .ZN(W40470));
  NANDX1 G24402 (.A1(W8839), .A2(W6965), .ZN(O10923));
  NANDX1 G24403 (.A1(W18695), .A2(W10589), .ZN(O10918));
  NANDX1 G24404 (.A1(W15692), .A2(W19590), .ZN(W40461));
  NANDX1 G24405 (.A1(I786), .A2(W14272), .ZN(O10908));
  NANDX1 G24406 (.A1(W14612), .A2(W33038), .ZN(O10769));
  NANDX1 G24407 (.A1(W2085), .A2(W22442), .ZN(O10790));
  NANDX1 G24408 (.A1(W10489), .A2(W37187), .ZN(O10789));
  NANDX1 G24409 (.A1(W13871), .A2(W38904), .ZN(W40266));
  NANDX1 G24410 (.A1(W15551), .A2(I382), .ZN(O10780));
  NANDX1 G24411 (.A1(W17147), .A2(W31597), .ZN(O10779));
  NANDX1 G24412 (.A1(W28961), .A2(W17543), .ZN(O10778));
  NANDX1 G24413 (.A1(W20675), .A2(W32795), .ZN(W40257));
  NANDX1 G24414 (.A1(W32444), .A2(W2298), .ZN(W40256));
  NANDX1 G24415 (.A1(W11815), .A2(W5305), .ZN(O10777));
  NANDX1 G24416 (.A1(W27648), .A2(W31573), .ZN(O10776));
  NANDX1 G24417 (.A1(W23001), .A2(W24244), .ZN(W40249));
  NANDX1 G24418 (.A1(W17603), .A2(W6450), .ZN(O10770));
  NANDX1 G24419 (.A1(I787), .A2(W17632), .ZN(O10791));
  NANDX1 G24420 (.A1(I1170), .A2(W39301), .ZN(O10766));
  NANDX1 G24421 (.A1(W930), .A2(W26260), .ZN(O10761));
  NANDX1 G24422 (.A1(W38598), .A2(W7595), .ZN(O10760));
  NANDX1 G24423 (.A1(W35160), .A2(W4951), .ZN(W40225));
  NANDX1 G24424 (.A1(W14606), .A2(W21972), .ZN(O10752));
  NANDX1 G24425 (.A1(W31951), .A2(W26659), .ZN(W40216));
  NANDX1 G24426 (.A1(W39450), .A2(W19254), .ZN(O10747));
  NANDX1 G24427 (.A1(W23908), .A2(W17553), .ZN(O10739));
  NANDX1 G24428 (.A1(W26694), .A2(I1222), .ZN(O10735));
  NANDX1 G24429 (.A1(W18025), .A2(W19404), .ZN(O10734));
  NANDX1 G24430 (.A1(W36533), .A2(W24322), .ZN(W40196));
  NANDX1 G24431 (.A1(W2810), .A2(W27735), .ZN(O10811));
  NANDX1 G24432 (.A1(W35854), .A2(W20464), .ZN(O10827));
  NANDX1 G24433 (.A1(W27415), .A2(W23002), .ZN(O10826));
  NANDX1 G24434 (.A1(W21661), .A2(W750), .ZN(O10825));
  NANDX1 G24435 (.A1(W37877), .A2(W19702), .ZN(O10823));
  NANDX1 G24436 (.A1(W15946), .A2(W39188), .ZN(O10822));
  NANDX1 G24437 (.A1(W35172), .A2(I1608), .ZN(W40336));
  NANDX1 G24438 (.A1(W21310), .A2(W9011), .ZN(O10818));
  NANDX1 G24439 (.A1(W38868), .A2(W32947), .ZN(W40326));
  NANDX1 G24440 (.A1(W39028), .A2(W20710), .ZN(W40324));
  NANDX1 G24441 (.A1(I1380), .A2(W20661), .ZN(W40322));
  NANDX1 G24442 (.A1(W16247), .A2(W7029), .ZN(W40319));
  NANDX1 G24443 (.A1(W15834), .A2(W29986), .ZN(O10959));
  NANDX1 G24444 (.A1(W5090), .A2(W27096), .ZN(W40315));
  NANDX1 G24445 (.A1(W19937), .A2(W21624), .ZN(O10808));
  NANDX1 G24446 (.A1(W31863), .A2(W13872), .ZN(W40308));
  NANDX1 G24447 (.A1(W20608), .A2(W25917), .ZN(W40303));
  NANDX1 G24448 (.A1(W29892), .A2(W32077), .ZN(O10801));
  NANDX1 G24449 (.A1(W26983), .A2(W31490), .ZN(O10798));
  NANDX1 G24450 (.A1(W33971), .A2(W12593), .ZN(W40292));
  NANDX1 G24451 (.A1(W10794), .A2(W39752), .ZN(W40291));
  NANDX1 G24452 (.A1(W12888), .A2(W16918), .ZN(O10794));
  NANDX1 G24453 (.A1(W17499), .A2(W23092), .ZN(W40285));
  NANDX1 G24454 (.A1(W6511), .A2(W32315), .ZN(O10792));
  NANDX1 G24455 (.A1(W29189), .A2(W27946), .ZN(O11111));
  NANDX1 G24456 (.A1(W24186), .A2(W5685), .ZN(O11139));
  NANDX1 G24457 (.A1(W4992), .A2(W36878), .ZN(O11131));
  NANDX1 G24458 (.A1(W9676), .A2(W11601), .ZN(W40764));
  NANDX1 G24459 (.A1(W28416), .A2(W23479), .ZN(O11130));
  NANDX1 G24460 (.A1(W13011), .A2(W3960), .ZN(O11129));
  NANDX1 G24461 (.A1(W13732), .A2(W38842), .ZN(W40758));
  NANDX1 G24462 (.A1(W26136), .A2(W16598), .ZN(O11124));
  NANDX1 G24463 (.A1(W12103), .A2(W31659), .ZN(O11123));
  NANDX1 G24464 (.A1(W39971), .A2(W2125), .ZN(O11122));
  NANDX1 G24465 (.A1(W19139), .A2(W24889), .ZN(O11120));
  NANDX1 G24466 (.A1(W3956), .A2(W13804), .ZN(O11116));
  NANDX1 G24467 (.A1(I755), .A2(W24551), .ZN(O11114));
  NANDX1 G24468 (.A1(W40114), .A2(W18263), .ZN(W40776));
  NANDX1 G24469 (.A1(W15187), .A2(W13174), .ZN(W40737));
  NANDX1 G24470 (.A1(W24316), .A2(W27870), .ZN(O11110));
  NANDX1 G24471 (.A1(W34574), .A2(W34272), .ZN(O11109));
  NANDX1 G24472 (.A1(I977), .A2(W16144), .ZN(O11101));
  NANDX1 G24473 (.A1(W16454), .A2(W22512), .ZN(O11099));
  NANDX1 G24474 (.A1(W30993), .A2(W2217), .ZN(O11098));
  NANDX1 G24475 (.A1(W38756), .A2(W4956), .ZN(O11094));
  NANDX1 G24476 (.A1(W27833), .A2(W333), .ZN(O11093));
  NANDX1 G24477 (.A1(W22273), .A2(W28438), .ZN(O11084));
  NANDX1 G24478 (.A1(W14200), .A2(W32842), .ZN(O11083));
  NANDX1 G24479 (.A1(W35141), .A2(W13680), .ZN(O11079));
  NANDX1 G24480 (.A1(W6927), .A2(W17114), .ZN(O11165));
  NANDX1 G24481 (.A1(W18941), .A2(W23342), .ZN(O11185));
  NANDX1 G24482 (.A1(W32642), .A2(W17565), .ZN(W40839));
  NANDX1 G24483 (.A1(W3926), .A2(W36764), .ZN(O11181));
  NANDX1 G24484 (.A1(W26468), .A2(W20113), .ZN(O11178));
  NANDX1 G24485 (.A1(W34858), .A2(W24446), .ZN(O11176));
  NANDX1 G24486 (.A1(W9446), .A2(W13977), .ZN(W40830));
  NANDX1 G24487 (.A1(W28203), .A2(W21967), .ZN(O11172));
  NANDX1 G24488 (.A1(W32545), .A2(W10352), .ZN(O11171));
  NANDX1 G24489 (.A1(W19679), .A2(W9008), .ZN(O11170));
  NANDX1 G24490 (.A1(W18339), .A2(W19575), .ZN(O11169));
  NANDX1 G24491 (.A1(W31443), .A2(W3476), .ZN(O11166));
  NANDX1 G24492 (.A1(W21981), .A2(W10230), .ZN(O11077));
  NANDX1 G24493 (.A1(W7619), .A2(W37857), .ZN(O11164));
  NANDX1 G24494 (.A1(W22951), .A2(W36412), .ZN(O11163));
  NANDX1 G24495 (.A1(W36004), .A2(W37904), .ZN(O11162));
  NANDX1 G24496 (.A1(W12019), .A2(I494), .ZN(W40800));
  NANDX1 G24497 (.A1(W27508), .A2(W4250), .ZN(W40797));
  NANDX1 G24498 (.A1(W2823), .A2(W32212), .ZN(O11151));
  NANDX1 G24499 (.A1(W25855), .A2(W30115), .ZN(O11149));
  NANDX1 G24500 (.A1(W28475), .A2(W15179), .ZN(W40787));
  NANDX1 G24501 (.A1(W16872), .A2(W1933), .ZN(W40783));
  NANDX1 G24502 (.A1(W39775), .A2(W34128), .ZN(O11142));
  NANDX1 G24503 (.A1(W21092), .A2(W26254), .ZN(O11140));
  NANDX1 G24504 (.A1(W725), .A2(W27166), .ZN(O10981));
  NANDX1 G24505 (.A1(W39648), .A2(W10420), .ZN(O11021));
  NANDX1 G24506 (.A1(W33344), .A2(W15002), .ZN(W40608));
  NANDX1 G24507 (.A1(W22877), .A2(W27350), .ZN(W40604));
  NANDX1 G24508 (.A1(W32421), .A2(W16887), .ZN(O11017));
  NANDX1 G24509 (.A1(W11800), .A2(W23120), .ZN(O11012));
  NANDX1 G24510 (.A1(W32546), .A2(W18141), .ZN(W40577));
  NANDX1 G24511 (.A1(W11137), .A2(W15312), .ZN(O10995));
  NANDX1 G24512 (.A1(W19536), .A2(W35419), .ZN(O10992));
  NANDX1 G24513 (.A1(W19297), .A2(W38867), .ZN(W40565));
  NANDX1 G24514 (.A1(W18743), .A2(W23369), .ZN(O10987));
  NANDX1 G24515 (.A1(I44), .A2(W18322), .ZN(O10986));
  NANDX1 G24516 (.A1(W29756), .A2(W11378), .ZN(O10984));
  NANDX1 G24517 (.A1(W38272), .A2(W23775), .ZN(W40616));
  NANDX1 G24518 (.A1(W8528), .A2(W34880), .ZN(O10980));
  NANDX1 G24519 (.A1(W17657), .A2(W9917), .ZN(O10975));
  NANDX1 G24520 (.A1(W40291), .A2(W17926), .ZN(O10974));
  NANDX1 G24521 (.A1(W33607), .A2(W36649), .ZN(O10971));
  NANDX1 G24522 (.A1(W5660), .A2(W28637), .ZN(O10968));
  NANDX1 G24523 (.A1(I318), .A2(W2582), .ZN(W40532));
  NANDX1 G24524 (.A1(W31270), .A2(W12346), .ZN(O10966));
  NANDX1 G24525 (.A1(W19832), .A2(W20050), .ZN(O10963));
  NANDX1 G24526 (.A1(W16266), .A2(W39705), .ZN(W40526));
  NANDX1 G24527 (.A1(W22419), .A2(W26759), .ZN(O10961));
  NANDX1 G24528 (.A1(W31727), .A2(W1673), .ZN(O10960));
  NANDX1 G24529 (.A1(W25114), .A2(W19820), .ZN(O11055));
  NANDX1 G24530 (.A1(I861), .A2(W34024), .ZN(W40687));
  NANDX1 G24531 (.A1(W31370), .A2(W17722), .ZN(W40686));
  NANDX1 G24532 (.A1(W11740), .A2(W33839), .ZN(W40680));
  NANDX1 G24533 (.A1(W9452), .A2(W29588), .ZN(O11071));
  NANDX1 G24534 (.A1(W37431), .A2(W25004), .ZN(O11070));
  NANDX1 G24535 (.A1(W4687), .A2(W20248), .ZN(W40675));
  NANDX1 G24536 (.A1(W22809), .A2(I1912), .ZN(W40673));
  NANDX1 G24537 (.A1(W37914), .A2(W14530), .ZN(O11068));
  NANDX1 G24538 (.A1(I64), .A2(W3620), .ZN(O11062));
  NANDX1 G24539 (.A1(W32355), .A2(W29934), .ZN(O11061));
  NANDX1 G24540 (.A1(W30325), .A2(W31513), .ZN(O11056));
  NANDX1 G24541 (.A1(W21724), .A2(W34298), .ZN(W38939));
  NANDX1 G24542 (.A1(W20769), .A2(W27095), .ZN(O11051));
  NANDX1 G24543 (.A1(W19604), .A2(W3938), .ZN(O11050));
  NANDX1 G24544 (.A1(W34254), .A2(W35563), .ZN(W40646));
  NANDX1 G24545 (.A1(W14702), .A2(W9201), .ZN(W40639));
  NANDX1 G24546 (.A1(W21745), .A2(W33271), .ZN(O11039));
  NANDX1 G24547 (.A1(W27444), .A2(W10762), .ZN(W40630));
  NANDX1 G24548 (.A1(I18), .A2(W32270), .ZN(O11037));
  NANDX1 G24549 (.A1(W21989), .A2(W34265), .ZN(O11036));
  NANDX1 G24550 (.A1(W8672), .A2(W13712), .ZN(O11031));
  NANDX1 G24551 (.A1(W24787), .A2(W35596), .ZN(O11030));
  NANDX1 G24552 (.A1(W39527), .A2(I752), .ZN(O11029));
  NANDX1 G24553 (.A1(W11608), .A2(W2715), .ZN(W37321));
  NANDX1 G24554 (.A1(W33591), .A2(W4678), .ZN(W37364));
  NANDX1 G24555 (.A1(W5568), .A2(W6107), .ZN(W37362));
  NANDX1 G24556 (.A1(W9169), .A2(W6128), .ZN(O8935));
  NANDX1 G24557 (.A1(W25099), .A2(W5214), .ZN(O8934));
  NANDX1 G24558 (.A1(W12007), .A2(W22886), .ZN(O8932));
  NANDX1 G24559 (.A1(W32165), .A2(W26553), .ZN(O8929));
  NANDX1 G24560 (.A1(W17432), .A2(W24979), .ZN(W37341));
  NANDX1 G24561 (.A1(W21845), .A2(W7878), .ZN(O8919));
  NANDX1 G24562 (.A1(W12564), .A2(W1904), .ZN(O8917));
  NANDX1 G24563 (.A1(W25681), .A2(W2854), .ZN(O8916));
  NANDX1 G24564 (.A1(W13728), .A2(W14734), .ZN(W37324));
  NANDX1 G24565 (.A1(W19128), .A2(I1247), .ZN(W37323));
  NANDX1 G24566 (.A1(W36539), .A2(W405), .ZN(O8944));
  NANDX1 G24567 (.A1(W9154), .A2(W32055), .ZN(O8908));
  NANDX1 G24568 (.A1(W8524), .A2(W1251), .ZN(W37313));
  NANDX1 G24569 (.A1(W21603), .A2(W35201), .ZN(O8905));
  NANDX1 G24570 (.A1(W3026), .A2(W64), .ZN(O8904));
  NANDX1 G24571 (.A1(W10522), .A2(W4492), .ZN(O8895));
  NANDX1 G24572 (.A1(W35869), .A2(W21670), .ZN(O8893));
  NANDX1 G24573 (.A1(W8229), .A2(W9940), .ZN(O8891));
  NANDX1 G24574 (.A1(W19823), .A2(W6283), .ZN(O8885));
  NANDX1 G24575 (.A1(I1092), .A2(W24337), .ZN(W37280));
  NANDX1 G24576 (.A1(I736), .A2(W34367), .ZN(O8882));
  NANDX1 G24577 (.A1(W31792), .A2(W23354), .ZN(W37266));
  NANDX1 G24578 (.A1(W21779), .A2(W24306), .ZN(O8971));
  NANDX1 G24579 (.A1(W9602), .A2(W7520), .ZN(W37455));
  NANDX1 G24580 (.A1(W5685), .A2(W20232), .ZN(W37453));
  NANDX1 G24581 (.A1(W5363), .A2(W15265), .ZN(O8987));
  NANDX1 G24582 (.A1(W17416), .A2(W26605), .ZN(O8986));
  NANDX1 G24583 (.A1(W18953), .A2(W20667), .ZN(W37448));
  NANDX1 G24584 (.A1(W23948), .A2(W23050), .ZN(O8984));
  NANDX1 G24585 (.A1(W15675), .A2(W32269), .ZN(O8983));
  NANDX1 G24586 (.A1(W445), .A2(W14239), .ZN(W37440));
  NANDX1 G24587 (.A1(I337), .A2(W5948), .ZN(O8977));
  NANDX1 G24588 (.A1(W31335), .A2(W177), .ZN(O8976));
  NANDX1 G24589 (.A1(W26808), .A2(W5801), .ZN(W37425));
  NANDX1 G24590 (.A1(W9339), .A2(W4076), .ZN(O8972));
  NANDX1 G24591 (.A1(W32204), .A2(W36480), .ZN(O8874));
  NANDX1 G24592 (.A1(W19409), .A2(W31269), .ZN(W37405));
  NANDX1 G24593 (.A1(W17193), .A2(W2386), .ZN(W37404));
  NANDX1 G24594 (.A1(W32291), .A2(W29496), .ZN(O8962));
  NANDX1 G24595 (.A1(W14341), .A2(W24967), .ZN(O8960));
  NANDX1 G24596 (.A1(W37071), .A2(W20453), .ZN(O8958));
  NANDX1 G24597 (.A1(W8192), .A2(W8991), .ZN(W37392));
  NANDX1 G24598 (.A1(W26757), .A2(W17431), .ZN(O8955));
  NANDX1 G24599 (.A1(W15506), .A2(W13185), .ZN(W37388));
  NANDX1 G24600 (.A1(W11461), .A2(W25131), .ZN(O8951));
  NANDX1 G24601 (.A1(W29041), .A2(W31091), .ZN(W37373));
  NANDX1 G24602 (.A1(W28689), .A2(W4765), .ZN(O8945));
  NANDX1 G24603 (.A1(W9005), .A2(W414), .ZN(W37151));
  NANDX1 G24604 (.A1(W30937), .A2(W28868), .ZN(O8828));
  NANDX1 G24605 (.A1(W3192), .A2(W17004), .ZN(O8826));
  NANDX1 G24606 (.A1(W17368), .A2(W4494), .ZN(O8824));
  NANDX1 G24607 (.A1(W13586), .A2(W17377), .ZN(O8823));
  NANDX1 G24608 (.A1(W30781), .A2(W8052), .ZN(W37174));
  NANDX1 G24609 (.A1(W27484), .A2(W4348), .ZN(W37165));
  NANDX1 G24610 (.A1(W29500), .A2(W24254), .ZN(W37164));
  NANDX1 G24611 (.A1(W20443), .A2(W16826), .ZN(W37162));
  NANDX1 G24612 (.A1(W7595), .A2(W14123), .ZN(W37158));
  NANDX1 G24613 (.A1(W14877), .A2(W28729), .ZN(O8810));
  NANDX1 G24614 (.A1(W18456), .A2(W4426), .ZN(O8809));
  NANDX1 G24615 (.A1(W7738), .A2(W6412), .ZN(O8808));
  NANDX1 G24616 (.A1(W26411), .A2(W22315), .ZN(O8829));
  NANDX1 G24617 (.A1(W4138), .A2(W4675), .ZN(O8803));
  NANDX1 G24618 (.A1(W21613), .A2(W5616), .ZN(W37140));
  NANDX1 G24619 (.A1(W27011), .A2(W27299), .ZN(O8802));
  NANDX1 G24620 (.A1(W29018), .A2(W36206), .ZN(O8801));
  NANDX1 G24621 (.A1(W23323), .A2(W21183), .ZN(O8800));
  NANDX1 G24622 (.A1(W23729), .A2(W7174), .ZN(O8794));
  NANDX1 G24623 (.A1(W34111), .A2(W37002), .ZN(O8793));
  NANDX1 G24624 (.A1(W3821), .A2(W8135), .ZN(O8791));
  NANDX1 G24625 (.A1(W34615), .A2(W9117), .ZN(O8790));
  NANDX1 G24626 (.A1(W26633), .A2(W36821), .ZN(O8789));
  NANDX1 G24627 (.A1(W1331), .A2(W1639), .ZN(W37112));
  NANDX1 G24628 (.A1(W2349), .A2(W1658), .ZN(W37220));
  NANDX1 G24629 (.A1(I1318), .A2(W11346), .ZN(W37263));
  NANDX1 G24630 (.A1(W26185), .A2(W11025), .ZN(O8873));
  NANDX1 G24631 (.A1(W8094), .A2(W1102), .ZN(W37257));
  NANDX1 G24632 (.A1(W22264), .A2(W20690), .ZN(W37256));
  NANDX1 G24633 (.A1(W17894), .A2(W2223), .ZN(O8872));
  NANDX1 G24634 (.A1(W18201), .A2(W4351), .ZN(W37253));
  NANDX1 G24635 (.A1(W18412), .A2(W9774), .ZN(O8869));
  NANDX1 G24636 (.A1(W18800), .A2(W8762), .ZN(O8865));
  NANDX1 G24637 (.A1(W13656), .A2(W19881), .ZN(O8860));
  NANDX1 G24638 (.A1(W20165), .A2(W29302), .ZN(O8856));
  NANDX1 G24639 (.A1(W1907), .A2(W24921), .ZN(O8849));
  NANDX1 G24640 (.A1(W27422), .A2(W1887), .ZN(O8992));
  NANDX1 G24641 (.A1(W11536), .A2(W24656), .ZN(O8848));
  NANDX1 G24642 (.A1(W15262), .A2(W8927), .ZN(O8847));
  NANDX1 G24643 (.A1(W22007), .A2(W10227), .ZN(O8840));
  NANDX1 G24644 (.A1(W21294), .A2(I1478), .ZN(O8837));
  NANDX1 G24645 (.A1(W35701), .A2(W32334), .ZN(W37200));
  NANDX1 G24646 (.A1(W10263), .A2(I428), .ZN(W37197));
  NANDX1 G24647 (.A1(W8401), .A2(W33449), .ZN(O8836));
  NANDX1 G24648 (.A1(W413), .A2(W26290), .ZN(O8834));
  NANDX1 G24649 (.A1(W6395), .A2(W36914), .ZN(W37190));
  NANDX1 G24650 (.A1(W26823), .A2(I737), .ZN(O8831));
  NANDX1 G24651 (.A1(W1654), .A2(W11969), .ZN(W37183));
  NANDX1 G24652 (.A1(W5355), .A2(W2838), .ZN(W37628));
  NANDX1 G24653 (.A1(W6469), .A2(W5452), .ZN(W37680));
  NANDX1 G24654 (.A1(W37049), .A2(W9251), .ZN(W37679));
  NANDX1 G24655 (.A1(W31917), .A2(W20020), .ZN(O9124));
  NANDX1 G24656 (.A1(W10635), .A2(W30528), .ZN(O9115));
  NANDX1 G24657 (.A1(W8468), .A2(W21450), .ZN(O9111));
  NANDX1 G24658 (.A1(W6647), .A2(W24133), .ZN(O9108));
  NANDX1 G24659 (.A1(W1629), .A2(W15491), .ZN(O9106));
  NANDX1 G24660 (.A1(W14892), .A2(W31119), .ZN(W37657));
  NANDX1 G24661 (.A1(W33803), .A2(W36999), .ZN(W37651));
  NANDX1 G24662 (.A1(W25624), .A2(W917), .ZN(O9098));
  NANDX1 G24663 (.A1(W2961), .A2(W20030), .ZN(O9095));
  NANDX1 G24664 (.A1(W14052), .A2(W18989), .ZN(O9094));
  NANDX1 G24665 (.A1(I1022), .A2(W1764), .ZN(O9126));
  NANDX1 G24666 (.A1(W8002), .A2(W14574), .ZN(O9085));
  NANDX1 G24667 (.A1(W13676), .A2(W35284), .ZN(O9083));
  NANDX1 G24668 (.A1(W30682), .A2(W858), .ZN(W37621));
  NANDX1 G24669 (.A1(I390), .A2(W27395), .ZN(O9081));
  NANDX1 G24670 (.A1(W18100), .A2(W12013), .ZN(O9080));
  NANDX1 G24671 (.A1(W22491), .A2(W32416), .ZN(W37611));
  NANDX1 G24672 (.A1(W20256), .A2(W36617), .ZN(W37610));
  NANDX1 G24673 (.A1(W18561), .A2(W2459), .ZN(O9077));
  NANDX1 G24674 (.A1(W4193), .A2(W23298), .ZN(O9072));
  NANDX1 G24675 (.A1(W2639), .A2(W34723), .ZN(O9071));
  NANDX1 G24676 (.A1(W10192), .A2(W12162), .ZN(O9070));
  NANDX1 G24677 (.A1(W7132), .A2(W24113), .ZN(W37713));
  NANDX1 G24678 (.A1(W20938), .A2(W18847), .ZN(W37744));
  NANDX1 G24679 (.A1(W25674), .A2(W11761), .ZN(O9160));
  NANDX1 G24680 (.A1(W34564), .A2(W30885), .ZN(O9158));
  NANDX1 G24681 (.A1(W8163), .A2(W27749), .ZN(W37738));
  NANDX1 G24682 (.A1(W12578), .A2(W9600), .ZN(W37737));
  NANDX1 G24683 (.A1(W27525), .A2(W14462), .ZN(O9156));
  NANDX1 G24684 (.A1(W11914), .A2(W23636), .ZN(O9154));
  NANDX1 G24685 (.A1(W35711), .A2(W27880), .ZN(O9150));
  NANDX1 G24686 (.A1(W23763), .A2(W35826), .ZN(O9149));
  NANDX1 G24687 (.A1(W13084), .A2(W4137), .ZN(W37726));
  NANDX1 G24688 (.A1(W37037), .A2(W20979), .ZN(W37723));
  NANDX1 G24689 (.A1(W8057), .A2(W17529), .ZN(W37715));
  NANDX1 G24690 (.A1(W1995), .A2(W13248), .ZN(W37588));
  NANDX1 G24691 (.A1(W36616), .A2(W27584), .ZN(W37712));
  NANDX1 G24692 (.A1(W32966), .A2(W35022), .ZN(O9140));
  NANDX1 G24693 (.A1(W2202), .A2(W29155), .ZN(W37706));
  NANDX1 G24694 (.A1(W15993), .A2(W4783), .ZN(W37703));
  NANDX1 G24695 (.A1(W34875), .A2(W14624), .ZN(W37702));
  NANDX1 G24696 (.A1(W23680), .A2(W12053), .ZN(O9136));
  NANDX1 G24697 (.A1(W37387), .A2(W23864), .ZN(W37698));
  NANDX1 G24698 (.A1(I1684), .A2(W16516), .ZN(O9134));
  NANDX1 G24699 (.A1(W30918), .A2(W2655), .ZN(W37694));
  NANDX1 G24700 (.A1(W17276), .A2(W37489), .ZN(O9128));
  NANDX1 G24701 (.A1(W1558), .A2(W3073), .ZN(O9127));
  NANDX1 G24702 (.A1(W14243), .A2(W3066), .ZN(O9009));
  NANDX1 G24703 (.A1(W12484), .A2(W3043), .ZN(W37518));
  NANDX1 G24704 (.A1(W18972), .A2(W485), .ZN(W37515));
  NANDX1 G24705 (.A1(W10314), .A2(W9907), .ZN(W37514));
  NANDX1 G24706 (.A1(W845), .A2(W28322), .ZN(O9023));
  NANDX1 G24707 (.A1(W25255), .A2(W20152), .ZN(O9022));
  NANDX1 G24708 (.A1(W9258), .A2(W4680), .ZN(O9021));
  NANDX1 G24709 (.A1(W26698), .A2(W1835), .ZN(W37506));
  NANDX1 G24710 (.A1(W25235), .A2(W34484), .ZN(O9019));
  NANDX1 G24711 (.A1(W16936), .A2(W26631), .ZN(O9017));
  NANDX1 G24712 (.A1(W23707), .A2(W5974), .ZN(W37499));
  NANDX1 G24713 (.A1(W33751), .A2(W20640), .ZN(O9015));
  NANDX1 G24714 (.A1(W25254), .A2(W25693), .ZN(O9011));
  NANDX1 G24715 (.A1(W29133), .A2(W36825), .ZN(W37524));
  NANDX1 G24716 (.A1(W4719), .A2(W7182), .ZN(O9008));
  NANDX1 G24717 (.A1(W24609), .A2(W23881), .ZN(O9006));
  NANDX1 G24718 (.A1(W36584), .A2(W31940), .ZN(W37483));
  NANDX1 G24719 (.A1(W21972), .A2(W12269), .ZN(O9005));
  NANDX1 G24720 (.A1(W34714), .A2(W26222), .ZN(O9002));
  NANDX1 G24721 (.A1(W30047), .A2(W16334), .ZN(O8999));
  NANDX1 G24722 (.A1(W27153), .A2(W20843), .ZN(O8997));
  NANDX1 G24723 (.A1(W29739), .A2(W2548), .ZN(W37469));
  NANDX1 G24724 (.A1(W4528), .A2(W22288), .ZN(W37466));
  NANDX1 G24725 (.A1(W9203), .A2(W20656), .ZN(W37465));
  NANDX1 G24726 (.A1(W29912), .A2(W1087), .ZN(W37464));
  NANDX1 G24727 (.A1(W31915), .A2(W6429), .ZN(O9046));
  NANDX1 G24728 (.A1(W29181), .A2(W24707), .ZN(O9065));
  NANDX1 G24729 (.A1(W37212), .A2(W5434), .ZN(W37586));
  NANDX1 G24730 (.A1(W24781), .A2(W9809), .ZN(W37585));
  NANDX1 G24731 (.A1(W22663), .A2(W20244), .ZN(O9064));
  NANDX1 G24732 (.A1(W31642), .A2(W33856), .ZN(O9062));
  NANDX1 G24733 (.A1(W6560), .A2(W21009), .ZN(O9057));
  NANDX1 G24734 (.A1(W26977), .A2(W34807), .ZN(W37567));
  NANDX1 G24735 (.A1(W1346), .A2(W307), .ZN(O9052));
  NANDX1 G24736 (.A1(W676), .A2(W23581), .ZN(O9048));
  NANDX1 G24737 (.A1(W25135), .A2(W22254), .ZN(O9047));
  NANDX1 G24738 (.A1(W24516), .A2(W29895), .ZN(W37553));
  NANDX1 G24739 (.A1(W36365), .A2(W2760), .ZN(W37106));
  NANDX1 G24740 (.A1(W15395), .A2(W15434), .ZN(W37551));
  NANDX1 G24741 (.A1(I843), .A2(W10497), .ZN(W37543));
  NANDX1 G24742 (.A1(W18171), .A2(W9530), .ZN(W37542));
  NANDX1 G24743 (.A1(W3764), .A2(W32426), .ZN(W37541));
  NANDX1 G24744 (.A1(W11833), .A2(W31684), .ZN(W37540));
  NANDX1 G24745 (.A1(I1703), .A2(W11604), .ZN(O9038));
  NANDX1 G24746 (.A1(W25411), .A2(W23930), .ZN(O9036));
  NANDX1 G24747 (.A1(W11662), .A2(W13513), .ZN(O9035));
  NANDX1 G24748 (.A1(W1532), .A2(W18971), .ZN(O9034));
  NANDX1 G24749 (.A1(W28073), .A2(I1390), .ZN(W37527));
  NANDX1 G24750 (.A1(W12100), .A2(W19263), .ZN(O9029));
  NANDX1 G24751 (.A1(W35166), .A2(W332), .ZN(W36664));
  NANDX1 G24752 (.A1(W8873), .A2(W34106), .ZN(O8554));
  NANDX1 G24753 (.A1(I914), .A2(W18671), .ZN(O8553));
  NANDX1 G24754 (.A1(W6150), .A2(W12676), .ZN(O8550));
  NANDX1 G24755 (.A1(W35177), .A2(W8632), .ZN(O8549));
  NANDX1 G24756 (.A1(W29259), .A2(W24072), .ZN(O8546));
  NANDX1 G24757 (.A1(I1727), .A2(W8043), .ZN(O8544));
  NANDX1 G24758 (.A1(W28905), .A2(W11331), .ZN(O8539));
  NANDX1 G24759 (.A1(W17973), .A2(W27232), .ZN(O8537));
  NANDX1 G24760 (.A1(W1159), .A2(W29027), .ZN(O8536));
  NANDX1 G24761 (.A1(W5226), .A2(W19665), .ZN(O8533));
  NANDX1 G24762 (.A1(W17863), .A2(W6326), .ZN(W36666));
  NANDX1 G24763 (.A1(W24500), .A2(W35259), .ZN(W36665));
  NANDX1 G24764 (.A1(W13852), .A2(W9504), .ZN(W36710));
  NANDX1 G24765 (.A1(W31449), .A2(W16722), .ZN(O8530));
  NANDX1 G24766 (.A1(W29995), .A2(W20236), .ZN(W36659));
  NANDX1 G24767 (.A1(W4368), .A2(W7977), .ZN(O8528));
  NANDX1 G24768 (.A1(W30135), .A2(W28242), .ZN(O8525));
  NANDX1 G24769 (.A1(W20679), .A2(W28682), .ZN(W36654));
  NANDX1 G24770 (.A1(W34262), .A2(W29740), .ZN(W36652));
  NANDX1 G24771 (.A1(W15428), .A2(W34507), .ZN(W36650));
  NANDX1 G24772 (.A1(W26224), .A2(W5589), .ZN(W36648));
  NANDX1 G24773 (.A1(W26769), .A2(W22798), .ZN(W36640));
  NANDX1 G24774 (.A1(W8811), .A2(W3447), .ZN(O8518));
  NANDX1 G24775 (.A1(W29104), .A2(W2182), .ZN(O8517));
  NANDX1 G24776 (.A1(W28205), .A2(W19463), .ZN(O8573));
  NANDX1 G24777 (.A1(W6627), .A2(W28084), .ZN(O8584));
  NANDX1 G24778 (.A1(W4201), .A2(W28960), .ZN(W36764));
  NANDX1 G24779 (.A1(W30159), .A2(W28038), .ZN(O8583));
  NANDX1 G24780 (.A1(I574), .A2(W11569), .ZN(O8582));
  NANDX1 G24781 (.A1(W16148), .A2(W18896), .ZN(O8581));
  NANDX1 G24782 (.A1(W11622), .A2(W31533), .ZN(O8580));
  NANDX1 G24783 (.A1(I552), .A2(W71), .ZN(O8576));
  NANDX1 G24784 (.A1(W23403), .A2(W11691), .ZN(O8575));
  NANDX1 G24785 (.A1(W35143), .A2(W7153), .ZN(W36749));
  NANDX1 G24786 (.A1(W22178), .A2(I430), .ZN(O8574));
  NANDX1 G24787 (.A1(W36154), .A2(W15167), .ZN(W36746));
  NANDX1 G24788 (.A1(W13435), .A2(W8147), .ZN(W36745));
  NANDX1 G24789 (.A1(W28298), .A2(W21489), .ZN(O8516));
  NANDX1 G24790 (.A1(W11097), .A2(W2413), .ZN(O8571));
  NANDX1 G24791 (.A1(W12661), .A2(W12690), .ZN(O8568));
  NANDX1 G24792 (.A1(I846), .A2(W32715), .ZN(W36733));
  NANDX1 G24793 (.A1(W33576), .A2(W16901), .ZN(O8564));
  NANDX1 G24794 (.A1(W3218), .A2(W28101), .ZN(W36726));
  NANDX1 G24795 (.A1(W1942), .A2(W10060), .ZN(O8563));
  NANDX1 G24796 (.A1(W25697), .A2(W23695), .ZN(W36723));
  NANDX1 G24797 (.A1(W28553), .A2(W1795), .ZN(W36717));
  NANDX1 G24798 (.A1(W7045), .A2(W24774), .ZN(O8560));
  NANDX1 G24799 (.A1(W30851), .A2(W337), .ZN(O8559));
  NANDX1 G24800 (.A1(W5401), .A2(W28488), .ZN(O8557));
  NANDX1 G24801 (.A1(W6273), .A2(W13410), .ZN(O8454));
  NANDX1 G24802 (.A1(W4346), .A2(W6391), .ZN(O8478));
  NANDX1 G24803 (.A1(W18300), .A2(W596), .ZN(O8477));
  NANDX1 G24804 (.A1(W26562), .A2(W11335), .ZN(O8475));
  NANDX1 G24805 (.A1(W12586), .A2(W34815), .ZN(O8474));
  NANDX1 G24806 (.A1(W23967), .A2(W24861), .ZN(O8472));
  NANDX1 G24807 (.A1(W15509), .A2(W6451), .ZN(W36556));
  NANDX1 G24808 (.A1(W10759), .A2(W23910), .ZN(O8466));
  NANDX1 G24809 (.A1(W25503), .A2(W7461), .ZN(O8464));
  NANDX1 G24810 (.A1(W735), .A2(W18601), .ZN(O8462));
  NANDX1 G24811 (.A1(W13076), .A2(W5381), .ZN(O8461));
  NANDX1 G24812 (.A1(W20943), .A2(W34887), .ZN(W36539));
  NANDX1 G24813 (.A1(W36021), .A2(W29043), .ZN(O8457));
  NANDX1 G24814 (.A1(W13981), .A2(W35528), .ZN(W36572));
  NANDX1 G24815 (.A1(W1327), .A2(W3264), .ZN(W36524));
  NANDX1 G24816 (.A1(W12590), .A2(W32951), .ZN(O8449));
  NANDX1 G24817 (.A1(W9849), .A2(W6517), .ZN(O8446));
  NANDX1 G24818 (.A1(W15635), .A2(W18404), .ZN(O8443));
  NANDX1 G24819 (.A1(W14930), .A2(W34232), .ZN(O8442));
  NANDX1 G24820 (.A1(W21382), .A2(W32945), .ZN(O8440));
  NANDX1 G24821 (.A1(W17464), .A2(W31402), .ZN(W36502));
  NANDX1 G24822 (.A1(W14041), .A2(W19804), .ZN(W36501));
  NANDX1 G24823 (.A1(W503), .A2(W17007), .ZN(O8436));
  NANDX1 G24824 (.A1(W28527), .A2(W5836), .ZN(W36499));
  NANDX1 G24825 (.A1(W19108), .A2(W14250), .ZN(O8431));
  NANDX1 G24826 (.A1(W27068), .A2(I1300), .ZN(W36598));
  NANDX1 G24827 (.A1(W22547), .A2(W15996), .ZN(W36634));
  NANDX1 G24828 (.A1(W3700), .A2(W32755), .ZN(W36630));
  NANDX1 G24829 (.A1(W27826), .A2(W26960), .ZN(O8513));
  NANDX1 G24830 (.A1(W7431), .A2(W7158), .ZN(O8510));
  NANDX1 G24831 (.A1(W1676), .A2(W30244), .ZN(W36617));
  NANDX1 G24832 (.A1(W17354), .A2(W25305), .ZN(O8504));
  NANDX1 G24833 (.A1(W18467), .A2(W19722), .ZN(O8503));
  NANDX1 G24834 (.A1(W12035), .A2(W36599), .ZN(O8501));
  NANDX1 G24835 (.A1(W3754), .A2(W14212), .ZN(O8500));
  NANDX1 G24836 (.A1(W6002), .A2(W32976), .ZN(O8499));
  NANDX1 G24837 (.A1(W8512), .A2(W32900), .ZN(O8495));
  NANDX1 G24838 (.A1(W5917), .A2(W7835), .ZN(W36770));
  NANDX1 G24839 (.A1(W29154), .A2(W12922), .ZN(W36596));
  NANDX1 G24840 (.A1(W34083), .A2(W10909), .ZN(W36593));
  NANDX1 G24841 (.A1(W16205), .A2(W18150), .ZN(O8491));
  NANDX1 G24842 (.A1(W7993), .A2(W14074), .ZN(W36587));
  NANDX1 G24843 (.A1(W1071), .A2(W35508), .ZN(W36586));
  NANDX1 G24844 (.A1(W36341), .A2(W29227), .ZN(O8487));
  NANDX1 G24845 (.A1(W2377), .A2(I1604), .ZN(W36580));
  NANDX1 G24846 (.A1(W33212), .A2(W13481), .ZN(W36579));
  NANDX1 G24847 (.A1(W17782), .A2(W14610), .ZN(W36577));
  NANDX1 G24848 (.A1(W14446), .A2(W15365), .ZN(O8484));
  NANDX1 G24849 (.A1(W13028), .A2(W2561), .ZN(O8483));
  NANDX1 G24850 (.A1(W15062), .A2(W25621), .ZN(W37008));
  NANDX1 G24851 (.A1(W16287), .A2(W3750), .ZN(W37037));
  NANDX1 G24852 (.A1(W13366), .A2(W35714), .ZN(O8736));
  NANDX1 G24853 (.A1(W14563), .A2(W23090), .ZN(W37025));
  NANDX1 G24854 (.A1(W6646), .A2(W25372), .ZN(O8732));
  NANDX1 G24855 (.A1(W2789), .A2(W12149), .ZN(W37023));
  NANDX1 G24856 (.A1(W3540), .A2(W32525), .ZN(W37022));
  NANDX1 G24857 (.A1(W2544), .A2(W34140), .ZN(W37019));
  NANDX1 G24858 (.A1(W30789), .A2(W9283), .ZN(O8731));
  NANDX1 G24859 (.A1(W11618), .A2(W17801), .ZN(W37017));
  NANDX1 G24860 (.A1(W15464), .A2(W35765), .ZN(W37016));
  NANDX1 G24861 (.A1(W31118), .A2(W313), .ZN(O8729));
  NANDX1 G24862 (.A1(W30012), .A2(W28189), .ZN(O8727));
  NANDX1 G24863 (.A1(I1394), .A2(W6873), .ZN(O8740));
  NANDX1 G24864 (.A1(W22674), .A2(W35173), .ZN(W37003));
  NANDX1 G24865 (.A1(W33346), .A2(W27717), .ZN(W37000));
  NANDX1 G24866 (.A1(W26508), .A2(W1356), .ZN(O8723));
  NANDX1 G24867 (.A1(I1650), .A2(W36460), .ZN(W36995));
  NANDX1 G24868 (.A1(W905), .A2(W3121), .ZN(O8722));
  NANDX1 G24869 (.A1(W11668), .A2(W4512), .ZN(W36989));
  NANDX1 G24870 (.A1(W97), .A2(W29511), .ZN(W36988));
  NANDX1 G24871 (.A1(W33455), .A2(W166), .ZN(O8718));
  NANDX1 G24872 (.A1(W11061), .A2(W11971), .ZN(O8717));
  NANDX1 G24873 (.A1(W18532), .A2(W33780), .ZN(O8711));
  NANDX1 G24874 (.A1(W27887), .A2(W35489), .ZN(O8708));
  NANDX1 G24875 (.A1(W23978), .A2(W32180), .ZN(W37071));
  NANDX1 G24876 (.A1(W1937), .A2(W11491), .ZN(O8782));
  NANDX1 G24877 (.A1(W7491), .A2(W22417), .ZN(O8780));
  NANDX1 G24878 (.A1(W24067), .A2(I1463), .ZN(W37099));
  NANDX1 G24879 (.A1(W31847), .A2(W16640), .ZN(W37094));
  NANDX1 G24880 (.A1(W8181), .A2(W35884), .ZN(O8774));
  NANDX1 G24881 (.A1(W694), .A2(W22076), .ZN(O8772));
  NANDX1 G24882 (.A1(W23293), .A2(W18686), .ZN(O8770));
  NANDX1 G24883 (.A1(W35769), .A2(W5927), .ZN(O8768));
  NANDX1 G24884 (.A1(W25972), .A2(W28202), .ZN(O8766));
  NANDX1 G24885 (.A1(W6146), .A2(W35549), .ZN(O8763));
  NANDX1 G24886 (.A1(W13529), .A2(W8314), .ZN(W37073));
  NANDX1 G24887 (.A1(W34195), .A2(W4025), .ZN(O8706));
  NANDX1 G24888 (.A1(W12196), .A2(W17169), .ZN(O8759));
  NANDX1 G24889 (.A1(W29727), .A2(I1457), .ZN(O8758));
  NANDX1 G24890 (.A1(I1473), .A2(W35920), .ZN(O8757));
  NANDX1 G24891 (.A1(W21950), .A2(W14367), .ZN(O8752));
  NANDX1 G24892 (.A1(W9536), .A2(W22821), .ZN(O8751));
  NANDX1 G24893 (.A1(W29155), .A2(W35815), .ZN(W37056));
  NANDX1 G24894 (.A1(W26264), .A2(W8538), .ZN(O8750));
  NANDX1 G24895 (.A1(W30364), .A2(W13209), .ZN(O8747));
  NANDX1 G24896 (.A1(W29069), .A2(W4786), .ZN(O8743));
  NANDX1 G24897 (.A1(W5621), .A2(W20059), .ZN(O8742));
  NANDX1 G24898 (.A1(W20947), .A2(W1534), .ZN(O8741));
  NANDX1 G24899 (.A1(W10106), .A2(W28557), .ZN(O8600));
  NANDX1 G24900 (.A1(W27388), .A2(W6136), .ZN(O8620));
  NANDX1 G24901 (.A1(W20989), .A2(W1998), .ZN(W36824));
  NANDX1 G24902 (.A1(W4215), .A2(W9500), .ZN(O8613));
  NANDX1 G24903 (.A1(W5752), .A2(W33769), .ZN(W36819));
  NANDX1 G24904 (.A1(W12456), .A2(W1171), .ZN(O8612));
  NANDX1 G24905 (.A1(W3516), .A2(W26019), .ZN(O8610));
  NANDX1 G24906 (.A1(W5902), .A2(W32572), .ZN(O8607));
  NANDX1 G24907 (.A1(W9906), .A2(W7968), .ZN(W36806));
  NANDX1 G24908 (.A1(W21768), .A2(W6704), .ZN(W36804));
  NANDX1 G24909 (.A1(W32317), .A2(W19226), .ZN(O8603));
  NANDX1 G24910 (.A1(W34202), .A2(I540), .ZN(W36797));
  NANDX1 G24911 (.A1(W31517), .A2(W15781), .ZN(O8601));
  NANDX1 G24912 (.A1(W28358), .A2(W16844), .ZN(W36832));
  NANDX1 G24913 (.A1(W4285), .A2(W26842), .ZN(O8599));
  NANDX1 G24914 (.A1(W31108), .A2(W10197), .ZN(W36790));
  NANDX1 G24915 (.A1(W16209), .A2(W25172), .ZN(W36788));
  NANDX1 G24916 (.A1(W13797), .A2(W5539), .ZN(O8598));
  NANDX1 G24917 (.A1(W26848), .A2(W32921), .ZN(O8594));
  NANDX1 G24918 (.A1(W3704), .A2(W23901), .ZN(W36780));
  NANDX1 G24919 (.A1(W8817), .A2(W14978), .ZN(W36779));
  NANDX1 G24920 (.A1(W34340), .A2(W35921), .ZN(O8590));
  NANDX1 G24921 (.A1(W5930), .A2(W11783), .ZN(W36773));
  NANDX1 G24922 (.A1(W2752), .A2(W12008), .ZN(W36772));
  NANDX1 G24923 (.A1(W19226), .A2(W23331), .ZN(O8588));
  NANDX1 G24924 (.A1(W26542), .A2(W21076), .ZN(O8661));
  NANDX1 G24925 (.A1(W19196), .A2(W35371), .ZN(O8705));
  NANDX1 G24926 (.A1(W28602), .A2(W9821), .ZN(W36959));
  NANDX1 G24927 (.A1(W25402), .A2(W33715), .ZN(O8698));
  NANDX1 G24928 (.A1(W20624), .A2(W23297), .ZN(O8688));
  NANDX1 G24929 (.A1(W15132), .A2(W8699), .ZN(O8687));
  NANDX1 G24930 (.A1(W3472), .A2(W36788), .ZN(O8683));
  NANDX1 G24931 (.A1(W29077), .A2(W28841), .ZN(W36931));
  NANDX1 G24932 (.A1(W20804), .A2(W27075), .ZN(O8675));
  NANDX1 G24933 (.A1(W3905), .A2(W5159), .ZN(O8669));
  NANDX1 G24934 (.A1(W14728), .A2(W15444), .ZN(O8668));
  NANDX1 G24935 (.A1(W33457), .A2(W21753), .ZN(O8667));
  NANDX1 G24936 (.A1(W35987), .A2(W11746), .ZN(W37745));
  NANDX1 G24937 (.A1(W18385), .A2(W4524), .ZN(O8659));
  NANDX1 G24938 (.A1(W8697), .A2(W6937), .ZN(O8653));
  NANDX1 G24939 (.A1(W33532), .A2(W16396), .ZN(W36886));
  NANDX1 G24940 (.A1(W261), .A2(W28793), .ZN(W36884));
  NANDX1 G24941 (.A1(I687), .A2(W20337), .ZN(O8647));
  NANDX1 G24942 (.A1(W1169), .A2(W16757), .ZN(O8645));
  NANDX1 G24943 (.A1(W5111), .A2(W14575), .ZN(W36872));
  NANDX1 G24944 (.A1(W25504), .A2(W6805), .ZN(W36858));
  NANDX1 G24945 (.A1(W20587), .A2(I1877), .ZN(O8634));
  NANDX1 G24946 (.A1(W5591), .A2(W1174), .ZN(W36846));
  NANDX1 G24947 (.A1(W29692), .A2(W2027), .ZN(O8629));
  NANDX1 G24948 (.A1(W4835), .A2(W25618), .ZN(O9652));
  NANDX1 G24949 (.A1(W4971), .A2(W24834), .ZN(O9671));
  NANDX1 G24950 (.A1(W15015), .A2(W7480), .ZN(O9670));
  NANDX1 G24951 (.A1(W19154), .A2(W19808), .ZN(W38593));
  NANDX1 G24952 (.A1(W23318), .A2(W26371), .ZN(W38590));
  NANDX1 G24953 (.A1(W18155), .A2(W15427), .ZN(O9668));
  NANDX1 G24954 (.A1(W4740), .A2(W30594), .ZN(O9661));
  NANDX1 G24955 (.A1(W17036), .A2(W22863), .ZN(O9659));
  NANDX1 G24956 (.A1(W8047), .A2(W9605), .ZN(O9656));
  NANDX1 G24957 (.A1(W3491), .A2(W11590), .ZN(W38566));
  NANDX1 G24958 (.A1(W29208), .A2(W20219), .ZN(O9654));
  NANDX1 G24959 (.A1(W30787), .A2(W31280), .ZN(W38563));
  NANDX1 G24960 (.A1(W4401), .A2(W9436), .ZN(W38560));
  NANDX1 G24961 (.A1(W10729), .A2(W36599), .ZN(W38598));
  NANDX1 G24962 (.A1(W19045), .A2(W28050), .ZN(W38556));
  NANDX1 G24963 (.A1(W3069), .A2(W19052), .ZN(O9650));
  NANDX1 G24964 (.A1(W29512), .A2(W36561), .ZN(O9649));
  NANDX1 G24965 (.A1(W20418), .A2(W13669), .ZN(O9646));
  NANDX1 G24966 (.A1(W9240), .A2(I219), .ZN(O9641));
  NANDX1 G24967 (.A1(W4219), .A2(W28176), .ZN(O9640));
  NANDX1 G24968 (.A1(W12036), .A2(W22569), .ZN(O9637));
  NANDX1 G24969 (.A1(W6343), .A2(W7767), .ZN(O9636));
  NANDX1 G24970 (.A1(W16838), .A2(W20479), .ZN(O9634));
  NANDX1 G24971 (.A1(W9245), .A2(I49), .ZN(O9632));
  NANDX1 G24972 (.A1(W29855), .A2(W12398), .ZN(O9630));
  NANDX1 G24973 (.A1(W7566), .A2(I919), .ZN(W38631));
  NANDX1 G24974 (.A1(W6808), .A2(W2322), .ZN(O9724));
  NANDX1 G24975 (.A1(W11854), .A2(W28079), .ZN(W38681));
  NANDX1 G24976 (.A1(W10171), .A2(W26545), .ZN(W38680));
  NANDX1 G24977 (.A1(I250), .A2(W23704), .ZN(O9722));
  NANDX1 G24978 (.A1(W21918), .A2(W12826), .ZN(W38675));
  NANDX1 G24979 (.A1(W12158), .A2(W23061), .ZN(O9719));
  NANDX1 G24980 (.A1(W8951), .A2(W10531), .ZN(W38670));
  NANDX1 G24981 (.A1(W10964), .A2(W38524), .ZN(O9716));
  NANDX1 G24982 (.A1(W2600), .A2(W7335), .ZN(O9701));
  NANDX1 G24983 (.A1(I858), .A2(W22806), .ZN(O9697));
  NANDX1 G24984 (.A1(W6550), .A2(W5428), .ZN(W38640));
  NANDX1 G24985 (.A1(W6400), .A2(W2872), .ZN(O9694));
  NANDX1 G24986 (.A1(I257), .A2(W38371), .ZN(O9627));
  NANDX1 G24987 (.A1(W27964), .A2(W6308), .ZN(O9688));
  NANDX1 G24988 (.A1(W30908), .A2(W25591), .ZN(W38622));
  NANDX1 G24989 (.A1(W16882), .A2(W15544), .ZN(O9687));
  NANDX1 G24990 (.A1(W1055), .A2(W17491), .ZN(O9682));
  NANDX1 G24991 (.A1(W12514), .A2(W32017), .ZN(W38613));
  NANDX1 G24992 (.A1(W22238), .A2(W13066), .ZN(O9678));
  NANDX1 G24993 (.A1(W2652), .A2(W18444), .ZN(W38608));
  NANDX1 G24994 (.A1(W26613), .A2(W30082), .ZN(O9676));
  NANDX1 G24995 (.A1(W3654), .A2(W3581), .ZN(O9675));
  NANDX1 G24996 (.A1(W2068), .A2(W18034), .ZN(O9673));
  NANDX1 G24997 (.A1(W32439), .A2(W36819), .ZN(W38601));
  NANDX1 G24998 (.A1(W31925), .A2(W19056), .ZN(O9544));
  NANDX1 G24999 (.A1(I785), .A2(W9266), .ZN(O9564));
  NANDX1 G25000 (.A1(W6170), .A2(W34997), .ZN(O9563));
  NANDX1 G25001 (.A1(W20763), .A2(W24724), .ZN(W38424));
  NANDX1 G25002 (.A1(W2803), .A2(W16212), .ZN(O9560));
  NANDX1 G25003 (.A1(I500), .A2(W3593), .ZN(W38418));
  NANDX1 G25004 (.A1(W6699), .A2(W3916), .ZN(W38416));
  NANDX1 G25005 (.A1(W17960), .A2(W30121), .ZN(O9557));
  NANDX1 G25006 (.A1(W19490), .A2(W12734), .ZN(W38412));
  NANDX1 G25007 (.A1(W20168), .A2(W33347), .ZN(O9555));
  NANDX1 G25008 (.A1(W13585), .A2(W23232), .ZN(O9549));
  NANDX1 G25009 (.A1(W32177), .A2(W3185), .ZN(O9547));
  NANDX1 G25010 (.A1(W37866), .A2(W12119), .ZN(O9546));
  NANDX1 G25011 (.A1(W18820), .A2(W17673), .ZN(O9566));
  NANDX1 G25012 (.A1(W28315), .A2(W15682), .ZN(W38389));
  NANDX1 G25013 (.A1(W25513), .A2(W31613), .ZN(W38384));
  NANDX1 G25014 (.A1(W31171), .A2(W29728), .ZN(O9535));
  NANDX1 G25015 (.A1(W626), .A2(W18918), .ZN(W38381));
  NANDX1 G25016 (.A1(W16085), .A2(W8156), .ZN(O9534));
  NANDX1 G25017 (.A1(W7535), .A2(W1691), .ZN(W38377));
  NANDX1 G25018 (.A1(I1639), .A2(I692), .ZN(O9531));
  NANDX1 G25019 (.A1(W29757), .A2(W26970), .ZN(O9525));
  NANDX1 G25020 (.A1(W5853), .A2(W29525), .ZN(O9522));
  NANDX1 G25021 (.A1(W23604), .A2(W26183), .ZN(O9521));
  NANDX1 G25022 (.A1(W31750), .A2(W21851), .ZN(W38356));
  NANDX1 G25023 (.A1(W20069), .A2(W14236), .ZN(O9594));
  NANDX1 G25024 (.A1(W24881), .A2(W38062), .ZN(W38519));
  NANDX1 G25025 (.A1(W19191), .A2(W20410), .ZN(O9621));
  NANDX1 G25026 (.A1(W22465), .A2(W20607), .ZN(O9620));
  NANDX1 G25027 (.A1(W37878), .A2(W26064), .ZN(O9618));
  NANDX1 G25028 (.A1(W14602), .A2(W29118), .ZN(W38506));
  NANDX1 G25029 (.A1(W20190), .A2(W30549), .ZN(W38491));
  NANDX1 G25030 (.A1(W8266), .A2(W24039), .ZN(O9606));
  NANDX1 G25031 (.A1(W15584), .A2(W22866), .ZN(O9603));
  NANDX1 G25032 (.A1(W15593), .A2(W16220), .ZN(W38479));
  NANDX1 G25033 (.A1(W12252), .A2(W3753), .ZN(O9600));
  NANDX1 G25034 (.A1(W37071), .A2(W15988), .ZN(O9596));
  NANDX1 G25035 (.A1(W32946), .A2(W31314), .ZN(O9725));
  NANDX1 G25036 (.A1(W9579), .A2(W21466), .ZN(W38464));
  NANDX1 G25037 (.A1(W8969), .A2(W26838), .ZN(O9593));
  NANDX1 G25038 (.A1(W4132), .A2(W30391), .ZN(O9586));
  NANDX1 G25039 (.A1(W36537), .A2(W8240), .ZN(W38455));
  NANDX1 G25040 (.A1(W1962), .A2(W38264), .ZN(W38454));
  NANDX1 G25041 (.A1(W15157), .A2(W18343), .ZN(O9584));
  NANDX1 G25042 (.A1(W11463), .A2(W36537), .ZN(W38449));
  NANDX1 G25043 (.A1(W19998), .A2(W10786), .ZN(W38446));
  NANDX1 G25044 (.A1(W24654), .A2(W34519), .ZN(O9574));
  NANDX1 G25045 (.A1(W3187), .A2(W26019), .ZN(O9573));
  NANDX1 G25046 (.A1(W23834), .A2(W37068), .ZN(W38435));
  NANDX1 G25047 (.A1(W33052), .A2(W3451), .ZN(W38842));
  NANDX1 G25048 (.A1(W25116), .A2(W18449), .ZN(W38867));
  NANDX1 G25049 (.A1(W24748), .A2(W30736), .ZN(O9834));
  NANDX1 G25050 (.A1(W32862), .A2(W738), .ZN(O9833));
  NANDX1 G25051 (.A1(W35400), .A2(W408), .ZN(O9831));
  NANDX1 G25052 (.A1(W35306), .A2(W32355), .ZN(W38855));
  NANDX1 G25053 (.A1(W8598), .A2(I942), .ZN(O9829));
  NANDX1 G25054 (.A1(W33434), .A2(W13546), .ZN(W38851));
  NANDX1 G25055 (.A1(W4204), .A2(W26806), .ZN(O9827));
  NANDX1 G25056 (.A1(W14936), .A2(W31526), .ZN(O9825));
  NANDX1 G25057 (.A1(W35779), .A2(W28327), .ZN(O9824));
  NANDX1 G25058 (.A1(W5274), .A2(W37573), .ZN(W38845));
  NANDX1 G25059 (.A1(W14882), .A2(W18183), .ZN(W38844));
  NANDX1 G25060 (.A1(W8820), .A2(W27115), .ZN(W38869));
  NANDX1 G25061 (.A1(W31162), .A2(W14468), .ZN(O9821));
  NANDX1 G25062 (.A1(W21201), .A2(W21006), .ZN(O9820));
  NANDX1 G25063 (.A1(W16861), .A2(W15109), .ZN(O9816));
  NANDX1 G25064 (.A1(W8859), .A2(W4482), .ZN(W38824));
  NANDX1 G25065 (.A1(W23415), .A2(W16544), .ZN(W38821));
  NANDX1 G25066 (.A1(W38375), .A2(W28823), .ZN(O9808));
  NANDX1 G25067 (.A1(W20917), .A2(W11173), .ZN(W38816));
  NANDX1 G25068 (.A1(W27167), .A2(W27599), .ZN(O9805));
  NANDX1 G25069 (.A1(W36248), .A2(W3722), .ZN(O9803));
  NANDX1 G25070 (.A1(W11460), .A2(W37642), .ZN(O9801));
  NANDX1 G25071 (.A1(W38161), .A2(W16019), .ZN(W38809));
  NANDX1 G25072 (.A1(W22250), .A2(W21977), .ZN(O9854));
  NANDX1 G25073 (.A1(W36432), .A2(W890), .ZN(O9872));
  NANDX1 G25074 (.A1(W19299), .A2(W25143), .ZN(O9865));
  NANDX1 G25075 (.A1(W18793), .A2(W34753), .ZN(W38923));
  NANDX1 G25076 (.A1(W3397), .A2(W10681), .ZN(W38921));
  NANDX1 G25077 (.A1(W22097), .A2(W1910), .ZN(O9864));
  NANDX1 G25078 (.A1(I1392), .A2(W387), .ZN(W38915));
  NANDX1 G25079 (.A1(W19414), .A2(W38557), .ZN(W38912));
  NANDX1 G25080 (.A1(W13160), .A2(W28750), .ZN(O9859));
  NANDX1 G25081 (.A1(W25276), .A2(W5991), .ZN(W38908));
  NANDX1 G25082 (.A1(W23870), .A2(W26200), .ZN(W38907));
  NANDX1 G25083 (.A1(W1907), .A2(W24728), .ZN(O9857));
  NANDX1 G25084 (.A1(W3069), .A2(W22177), .ZN(O9855));
  NANDX1 G25085 (.A1(W3648), .A2(W26425), .ZN(W38807));
  NANDX1 G25086 (.A1(W6245), .A2(W2332), .ZN(O9852));
  NANDX1 G25087 (.A1(W8491), .A2(W31287), .ZN(W38893));
  NANDX1 G25088 (.A1(W37134), .A2(W8035), .ZN(O9848));
  NANDX1 G25089 (.A1(W12187), .A2(W32313), .ZN(O9847));
  NANDX1 G25090 (.A1(W10401), .A2(W13643), .ZN(W38887));
  NANDX1 G25091 (.A1(W35344), .A2(W33103), .ZN(O9845));
  NANDX1 G25092 (.A1(W21078), .A2(W29997), .ZN(O9843));
  NANDX1 G25093 (.A1(W20839), .A2(W32575), .ZN(W38879));
  NANDX1 G25094 (.A1(W19581), .A2(W2112), .ZN(W38878));
  NANDX1 G25095 (.A1(W10838), .A2(W1498), .ZN(W38872));
  NANDX1 G25096 (.A1(W20194), .A2(W27111), .ZN(O9839));
  NANDX1 G25097 (.A1(W15598), .A2(W31260), .ZN(W38708));
  NANDX1 G25098 (.A1(W14174), .A2(W38231), .ZN(W38735));
  NANDX1 G25099 (.A1(W22292), .A2(W9702), .ZN(O9756));
  NANDX1 G25100 (.A1(W20316), .A2(W32123), .ZN(O9755));
  NANDX1 G25101 (.A1(W27952), .A2(W32324), .ZN(O9753));
  NANDX1 G25102 (.A1(W1913), .A2(W29617), .ZN(W38724));
  NANDX1 G25103 (.A1(W7972), .A2(W15903), .ZN(O9749));
  NANDX1 G25104 (.A1(W11992), .A2(W29423), .ZN(O9747));
  NANDX1 G25105 (.A1(W28671), .A2(W27204), .ZN(W38717));
  NANDX1 G25106 (.A1(W35759), .A2(W34453), .ZN(O9746));
  NANDX1 G25107 (.A1(W20370), .A2(W38644), .ZN(O9745));
  NANDX1 G25108 (.A1(W2422), .A2(W13818), .ZN(O9743));
  NANDX1 G25109 (.A1(W31531), .A2(W21459), .ZN(O9741));
  NANDX1 G25110 (.A1(W24087), .A2(W28476), .ZN(W38744));
  NANDX1 G25111 (.A1(W1039), .A2(W36226), .ZN(W38707));
  NANDX1 G25112 (.A1(W15477), .A2(W7868), .ZN(O9740));
  NANDX1 G25113 (.A1(W15650), .A2(W15308), .ZN(O9739));
  NANDX1 G25114 (.A1(W2438), .A2(W4900), .ZN(W38703));
  NANDX1 G25115 (.A1(W23670), .A2(W11326), .ZN(W38702));
  NANDX1 G25116 (.A1(W30005), .A2(W7087), .ZN(O9738));
  NANDX1 G25117 (.A1(W17233), .A2(W15524), .ZN(O9737));
  NANDX1 G25118 (.A1(W30728), .A2(W8218), .ZN(W38698));
  NANDX1 G25119 (.A1(W7806), .A2(W19299), .ZN(W38695));
  NANDX1 G25120 (.A1(W32921), .A2(W38115), .ZN(O9729));
  NANDX1 G25121 (.A1(W32003), .A2(W7379), .ZN(O9728));
  NANDX1 G25122 (.A1(W25151), .A2(W36779), .ZN(W38770));
  NANDX1 G25123 (.A1(W23971), .A2(W27537), .ZN(W38805));
  NANDX1 G25124 (.A1(W27753), .A2(W34792), .ZN(O9799));
  NANDX1 G25125 (.A1(I1308), .A2(W547), .ZN(O9796));
  NANDX1 G25126 (.A1(W9225), .A2(W12112), .ZN(O9795));
  NANDX1 G25127 (.A1(W30735), .A2(W8871), .ZN(O9788));
  NANDX1 G25128 (.A1(W14115), .A2(W1556), .ZN(O9787));
  NANDX1 G25129 (.A1(W20381), .A2(W18105), .ZN(W38785));
  NANDX1 G25130 (.A1(W21331), .A2(W33729), .ZN(W38782));
  NANDX1 G25131 (.A1(W21789), .A2(W27046), .ZN(O9781));
  NANDX1 G25132 (.A1(W32069), .A2(W36493), .ZN(W38776));
  NANDX1 G25133 (.A1(W38124), .A2(W23031), .ZN(W38772));
  NANDX1 G25134 (.A1(W34324), .A2(W29143), .ZN(W38353));
  NANDX1 G25135 (.A1(W1143), .A2(W1516), .ZN(O9776));
  NANDX1 G25136 (.A1(W13637), .A2(W7389), .ZN(O9775));
  NANDX1 G25137 (.A1(W14999), .A2(W7148), .ZN(O9772));
  NANDX1 G25138 (.A1(W14161), .A2(I1777), .ZN(W38761));
  NANDX1 G25139 (.A1(W14208), .A2(W11371), .ZN(O9770));
  NANDX1 G25140 (.A1(W18519), .A2(W36734), .ZN(W38754));
  NANDX1 G25141 (.A1(W29977), .A2(W28962), .ZN(W38752));
  NANDX1 G25142 (.A1(W16138), .A2(W25953), .ZN(W38751));
  NANDX1 G25143 (.A1(W14043), .A2(W24523), .ZN(O9766));
  NANDX1 G25144 (.A1(W21004), .A2(W25370), .ZN(W38748));
  NANDX1 G25145 (.A1(W591), .A2(W31924), .ZN(O9765));
  NANDX1 G25146 (.A1(I1195), .A2(W11179), .ZN(O9290));
  NANDX1 G25147 (.A1(W15100), .A2(I981), .ZN(W37973));
  NANDX1 G25148 (.A1(I1666), .A2(W21150), .ZN(W37969));
  NANDX1 G25149 (.A1(W560), .A2(I10), .ZN(W37968));
  NANDX1 G25150 (.A1(W30719), .A2(I1189), .ZN(W37967));
  NANDX1 G25151 (.A1(W15940), .A2(W2295), .ZN(W37966));
  NANDX1 G25152 (.A1(W807), .A2(W27955), .ZN(W37964));
  NANDX1 G25153 (.A1(W4769), .A2(W11196), .ZN(W37961));
  NANDX1 G25154 (.A1(W811), .A2(W10818), .ZN(W37958));
  NANDX1 G25155 (.A1(W12787), .A2(W27621), .ZN(O9297));
  NANDX1 G25156 (.A1(W8000), .A2(W18125), .ZN(O9296));
  NANDX1 G25157 (.A1(W4553), .A2(W32040), .ZN(O9294));
  NANDX1 G25158 (.A1(W36220), .A2(W28945), .ZN(W37952));
  NANDX1 G25159 (.A1(W18050), .A2(W36580), .ZN(O9303));
  NANDX1 G25160 (.A1(W3431), .A2(W30557), .ZN(O9289));
  NANDX1 G25161 (.A1(W13698), .A2(W22990), .ZN(O9288));
  NANDX1 G25162 (.A1(W31848), .A2(W30028), .ZN(W37939));
  NANDX1 G25163 (.A1(W33064), .A2(W13067), .ZN(W37938));
  NANDX1 G25164 (.A1(W8591), .A2(W23602), .ZN(W37937));
  NANDX1 G25165 (.A1(I1860), .A2(W34488), .ZN(O9285));
  NANDX1 G25166 (.A1(I986), .A2(W31544), .ZN(O9280));
  NANDX1 G25167 (.A1(W15917), .A2(W18153), .ZN(W37917));
  NANDX1 G25168 (.A1(W24794), .A2(W7828), .ZN(O9274));
  NANDX1 G25169 (.A1(W7855), .A2(W30548), .ZN(O9271));
  NANDX1 G25170 (.A1(W21661), .A2(W4748), .ZN(O9269));
  NANDX1 G25171 (.A1(W4496), .A2(W16286), .ZN(O9322));
  NANDX1 G25172 (.A1(W2271), .A2(W36608), .ZN(O9340));
  NANDX1 G25173 (.A1(W24466), .A2(W4244), .ZN(O9338));
  NANDX1 G25174 (.A1(W20208), .A2(W18013), .ZN(W38037));
  NANDX1 G25175 (.A1(W23793), .A2(W2102), .ZN(W38034));
  NANDX1 G25176 (.A1(W6645), .A2(W3860), .ZN(W38033));
  NANDX1 G25177 (.A1(W24722), .A2(W26706), .ZN(O9334));
  NANDX1 G25178 (.A1(W705), .A2(W32738), .ZN(O9332));
  NANDX1 G25179 (.A1(W24719), .A2(W603), .ZN(W38022));
  NANDX1 G25180 (.A1(W5777), .A2(W35233), .ZN(O9327));
  NANDX1 G25181 (.A1(W304), .A2(W29298), .ZN(W38015));
  NANDX1 G25182 (.A1(W229), .A2(W4520), .ZN(O9326));
  NANDX1 G25183 (.A1(W37252), .A2(W26060), .ZN(W38006));
  NANDX1 G25184 (.A1(W5226), .A2(W13780), .ZN(O9268));
  NANDX1 G25185 (.A1(I1076), .A2(W33983), .ZN(W38004));
  NANDX1 G25186 (.A1(W37321), .A2(W5482), .ZN(W38002));
  NANDX1 G25187 (.A1(W21126), .A2(W12808), .ZN(O9320));
  NANDX1 G25188 (.A1(W1463), .A2(W31768), .ZN(O9316));
  NANDX1 G25189 (.A1(W1816), .A2(W16146), .ZN(O9315));
  NANDX1 G25190 (.A1(W37812), .A2(W19295), .ZN(O9314));
  NANDX1 G25191 (.A1(W31970), .A2(W32422), .ZN(O9313));
  NANDX1 G25192 (.A1(W15414), .A2(W23620), .ZN(O9310));
  NANDX1 G25193 (.A1(W15692), .A2(W10714), .ZN(O9305));
  NANDX1 G25194 (.A1(W17951), .A2(W23313), .ZN(O9304));
  NANDX1 G25195 (.A1(W13810), .A2(W22571), .ZN(W37977));
  NANDX1 G25196 (.A1(W26803), .A2(W14247), .ZN(O9198));
  NANDX1 G25197 (.A1(W17603), .A2(W4902), .ZN(O9220));
  NANDX1 G25198 (.A1(I23), .A2(W28833), .ZN(O9218));
  NANDX1 G25199 (.A1(W33811), .A2(W27035), .ZN(O9213));
  NANDX1 G25200 (.A1(W31829), .A2(W8706), .ZN(O9212));
  NANDX1 G25201 (.A1(W8025), .A2(W11315), .ZN(W37822));
  NANDX1 G25202 (.A1(W23722), .A2(W32667), .ZN(W37821));
  NANDX1 G25203 (.A1(W3655), .A2(W4732), .ZN(O9207));
  NANDX1 G25204 (.A1(W25013), .A2(W25180), .ZN(W37810));
  NANDX1 G25205 (.A1(W19932), .A2(W33841), .ZN(O9203));
  NANDX1 G25206 (.A1(W26882), .A2(W36463), .ZN(O9202));
  NANDX1 G25207 (.A1(W19061), .A2(W37071), .ZN(O9200));
  NANDX1 G25208 (.A1(W26538), .A2(W25749), .ZN(O9199));
  NANDX1 G25209 (.A1(W6859), .A2(W12300), .ZN(O9222));
  NANDX1 G25210 (.A1(W3424), .A2(W19451), .ZN(W37803));
  NANDX1 G25211 (.A1(I583), .A2(W7655), .ZN(O9196));
  NANDX1 G25212 (.A1(W3637), .A2(W20240), .ZN(W37798));
  NANDX1 G25213 (.A1(W35646), .A2(W8569), .ZN(O9194));
  NANDX1 G25214 (.A1(W3678), .A2(W33715), .ZN(W37779));
  NANDX1 G25215 (.A1(W5993), .A2(W14145), .ZN(O9182));
  NANDX1 G25216 (.A1(W32240), .A2(W13328), .ZN(O9181));
  NANDX1 G25217 (.A1(W1008), .A2(W7259), .ZN(W37773));
  NANDX1 G25218 (.A1(W24191), .A2(W37557), .ZN(O9178));
  NANDX1 G25219 (.A1(W21754), .A2(W11898), .ZN(W37770));
  NANDX1 G25220 (.A1(W36945), .A2(W25572), .ZN(W37762));
  NANDX1 G25221 (.A1(W29242), .A2(W15754), .ZN(W37866));
  NANDX1 G25222 (.A1(W34259), .A2(W33201), .ZN(W37904));
  NANDX1 G25223 (.A1(W33174), .A2(W36161), .ZN(O9263));
  NANDX1 G25224 (.A1(W21807), .A2(I1280), .ZN(O9262));
  NANDX1 G25225 (.A1(W854), .A2(W34885), .ZN(W37896));
  NANDX1 G25226 (.A1(W21601), .A2(W15507), .ZN(O9261));
  NANDX1 G25227 (.A1(I753), .A2(W22928), .ZN(W37889));
  NANDX1 G25228 (.A1(W9796), .A2(W35934), .ZN(O9255));
  NANDX1 G25229 (.A1(W23216), .A2(W32485), .ZN(W37878));
  NANDX1 G25230 (.A1(W3756), .A2(W36813), .ZN(O9249));
  NANDX1 G25231 (.A1(W19702), .A2(W14414), .ZN(O9246));
  NANDX1 G25232 (.A1(W34073), .A2(W24786), .ZN(W37869));
  NANDX1 G25233 (.A1(W19519), .A2(W4337), .ZN(W38043));
  NANDX1 G25234 (.A1(W24335), .A2(W8712), .ZN(O9242));
  NANDX1 G25235 (.A1(W2278), .A2(W28595), .ZN(O9240));
  NANDX1 G25236 (.A1(W7853), .A2(W15199), .ZN(W37856));
  NANDX1 G25237 (.A1(W7713), .A2(W4433), .ZN(O9236));
  NANDX1 G25238 (.A1(W30538), .A2(W14672), .ZN(O9234));
  NANDX1 G25239 (.A1(W1278), .A2(W35573), .ZN(O9232));
  NANDX1 G25240 (.A1(W37404), .A2(W17836), .ZN(W37844));
  NANDX1 G25241 (.A1(W11110), .A2(W3466), .ZN(O9226));
  NANDX1 G25242 (.A1(W10539), .A2(W19504), .ZN(W37840));
  NANDX1 G25243 (.A1(I1993), .A2(W10018), .ZN(O9223));
  NANDX1 G25244 (.A1(W23688), .A2(W7326), .ZN(W37836));
  NANDX1 G25245 (.A1(W16739), .A2(W22547), .ZN(W38239));
  NANDX1 G25246 (.A1(W9768), .A2(W5482), .ZN(O9478));
  NANDX1 G25247 (.A1(W11749), .A2(W18992), .ZN(W38282));
  NANDX1 G25248 (.A1(W412), .A2(W36580), .ZN(O9477));
  NANDX1 G25249 (.A1(W6753), .A2(W30445), .ZN(O9474));
  NANDX1 G25250 (.A1(W9989), .A2(W12770), .ZN(W38276));
  NANDX1 G25251 (.A1(W13613), .A2(W13408), .ZN(W38271));
  NANDX1 G25252 (.A1(W36589), .A2(W30544), .ZN(W38264));
  NANDX1 G25253 (.A1(W2584), .A2(W296), .ZN(O9467));
  NANDX1 G25254 (.A1(W6749), .A2(W25810), .ZN(O9463));
  NANDX1 G25255 (.A1(W34100), .A2(W24469), .ZN(W38253));
  NANDX1 G25256 (.A1(W5069), .A2(W1525), .ZN(O9460));
  NANDX1 G25257 (.A1(W19892), .A2(W23849), .ZN(O9454));
  NANDX1 G25258 (.A1(W28358), .A2(W10418), .ZN(W38288));
  NANDX1 G25259 (.A1(W11928), .A2(W37139), .ZN(O9450));
  NANDX1 G25260 (.A1(I1011), .A2(W17370), .ZN(W38230));
  NANDX1 G25261 (.A1(W34165), .A2(W12968), .ZN(O9446));
  NANDX1 G25262 (.A1(W10721), .A2(W30341), .ZN(W38226));
  NANDX1 G25263 (.A1(W7254), .A2(W33774), .ZN(W38223));
  NANDX1 G25264 (.A1(W7197), .A2(W27098), .ZN(W38220));
  NANDX1 G25265 (.A1(W7414), .A2(W3071), .ZN(W38219));
  NANDX1 G25266 (.A1(W21053), .A2(W7227), .ZN(O9441));
  NANDX1 G25267 (.A1(W27801), .A2(W14109), .ZN(O9440));
  NANDX1 G25268 (.A1(W31834), .A2(W27271), .ZN(O9439));
  NANDX1 G25269 (.A1(W34580), .A2(W23110), .ZN(W38213));
  NANDX1 G25270 (.A1(W12177), .A2(W30111), .ZN(O9504));
  NANDX1 G25271 (.A1(W19832), .A2(W32933), .ZN(W38352));
  NANDX1 G25272 (.A1(W17162), .A2(W13722), .ZN(W38351));
  NANDX1 G25273 (.A1(W26469), .A2(I1677), .ZN(W38349));
  NANDX1 G25274 (.A1(W17484), .A2(W24914), .ZN(W38346));
  NANDX1 G25275 (.A1(W16148), .A2(W33715), .ZN(O9518));
  NANDX1 G25276 (.A1(W6078), .A2(W5475), .ZN(W38341));
  NANDX1 G25277 (.A1(W31383), .A2(W7764), .ZN(W38340));
  NANDX1 G25278 (.A1(W25524), .A2(W22564), .ZN(O9514));
  NANDX1 G25279 (.A1(W8742), .A2(W6866), .ZN(W38333));
  NANDX1 G25280 (.A1(W12637), .A2(W30591), .ZN(O9510));
  NANDX1 G25281 (.A1(W30132), .A2(W19802), .ZN(O9506));
  NANDX1 G25282 (.A1(W3436), .A2(W1230), .ZN(W38209));
  NANDX1 G25283 (.A1(W27730), .A2(W38305), .ZN(W38320));
  NANDX1 G25284 (.A1(W30103), .A2(W25971), .ZN(O9502));
  NANDX1 G25285 (.A1(W25949), .A2(W675), .ZN(O9501));
  NANDX1 G25286 (.A1(W25002), .A2(W25489), .ZN(O9497));
  NANDX1 G25287 (.A1(I1439), .A2(W14294), .ZN(O9492));
  NANDX1 G25288 (.A1(W3114), .A2(W6071), .ZN(O9491));
  NANDX1 G25289 (.A1(W13094), .A2(W8429), .ZN(W38298));
  NANDX1 G25290 (.A1(W29620), .A2(W25292), .ZN(W38297));
  NANDX1 G25291 (.A1(W7671), .A2(W2085), .ZN(O9488));
  NANDX1 G25292 (.A1(W33774), .A2(W13523), .ZN(O9485));
  NANDX1 G25293 (.A1(W32399), .A2(W16814), .ZN(O9484));
  NANDX1 G25294 (.A1(W31025), .A2(W34239), .ZN(O9362));
  NANDX1 G25295 (.A1(W36340), .A2(I61), .ZN(O9380));
  NANDX1 G25296 (.A1(I1654), .A2(W26077), .ZN(O9375));
  NANDX1 G25297 (.A1(W32728), .A2(W667), .ZN(W38102));
  NANDX1 G25298 (.A1(W20269), .A2(W10894), .ZN(O9374));
  NANDX1 G25299 (.A1(W10539), .A2(W32546), .ZN(O9370));
  NANDX1 G25300 (.A1(W31478), .A2(W33200), .ZN(O9368));
  NANDX1 G25301 (.A1(W18034), .A2(W36543), .ZN(W38091));
  NANDX1 G25302 (.A1(W22331), .A2(W36708), .ZN(W38089));
  NANDX1 G25303 (.A1(W30961), .A2(I1325), .ZN(W38088));
  NANDX1 G25304 (.A1(W18204), .A2(W24837), .ZN(W38087));
  NANDX1 G25305 (.A1(W2010), .A2(W29599), .ZN(W38084));
  NANDX1 G25306 (.A1(W7208), .A2(W27875), .ZN(W38082));
  NANDX1 G25307 (.A1(W24549), .A2(W1659), .ZN(O9383));
  NANDX1 G25308 (.A1(W5138), .A2(W12148), .ZN(W38078));
  NANDX1 G25309 (.A1(W19294), .A2(W27730), .ZN(O9361));
  NANDX1 G25310 (.A1(W19926), .A2(W25038), .ZN(W38075));
  NANDX1 G25311 (.A1(W7540), .A2(W6603), .ZN(O9360));
  NANDX1 G25312 (.A1(W14895), .A2(W27802), .ZN(W38067));
  NANDX1 G25313 (.A1(W15821), .A2(W13695), .ZN(O9354));
  NANDX1 G25314 (.A1(W36647), .A2(W4392), .ZN(W38061));
  NANDX1 G25315 (.A1(W19708), .A2(W35149), .ZN(O9348));
  NANDX1 G25316 (.A1(W18442), .A2(W826), .ZN(W38050));
  NANDX1 G25317 (.A1(W14888), .A2(W37823), .ZN(O9345));
  NANDX1 G25318 (.A1(W18477), .A2(W36164), .ZN(W38046));
  NANDX1 G25319 (.A1(W33884), .A2(W25289), .ZN(W38172));
  NANDX1 G25320 (.A1(W28345), .A2(W25069), .ZN(O9433));
  NANDX1 G25321 (.A1(W21785), .A2(W3737), .ZN(O9432));
  NANDX1 G25322 (.A1(W3644), .A2(W37899), .ZN(O9429));
  NANDX1 G25323 (.A1(W18483), .A2(W10118), .ZN(O9427));
  NANDX1 G25324 (.A1(W21997), .A2(W38102), .ZN(O9423));
  NANDX1 G25325 (.A1(W36208), .A2(W32487), .ZN(W38187));
  NANDX1 G25326 (.A1(W686), .A2(W14053), .ZN(W38186));
  NANDX1 G25327 (.A1(W22828), .A2(W23739), .ZN(W38185));
  NANDX1 G25328 (.A1(W17256), .A2(W19381), .ZN(W38184));
  NANDX1 G25329 (.A1(W5236), .A2(W27497), .ZN(W38181));
  NANDX1 G25330 (.A1(W14167), .A2(W28253), .ZN(O9418));
  NANDX1 G25331 (.A1(W18676), .A2(I349), .ZN(O5965));
  NANDX1 G25332 (.A1(I1881), .A2(W3132), .ZN(W38171));
  NANDX1 G25333 (.A1(W27962), .A2(W35130), .ZN(W38168));
  NANDX1 G25334 (.A1(W19124), .A2(W10712), .ZN(W38161));
  NANDX1 G25335 (.A1(I2), .A2(I3), .ZN(W1));
  NANDX1 G25336 (.A1(W36077), .A2(W16908), .ZN(O9406));
  NANDX1 G25337 (.A1(W36921), .A2(W23050), .ZN(O9402));
  NANDX1 G25338 (.A1(W20476), .A2(W35912), .ZN(W38141));
  NANDX1 G25339 (.A1(W35267), .A2(W37128), .ZN(O9393));
  NANDX1 G25340 (.A1(W21044), .A2(W23794), .ZN(O9391));
  NANDX1 G25341 (.A1(W9648), .A2(W26419), .ZN(O9388));
  NANDX1 G25342 (.A1(W7270), .A2(W7690), .ZN(O9385));
  NANDX1 G25343 (.A1(W1883), .A2(W2395), .ZN(W4512));
  NANDX1 G25344 (.A1(W1130), .A2(I870), .ZN(W4500));
  NANDX1 G25345 (.A1(W1019), .A2(W533), .ZN(W4501));
  NANDX1 G25346 (.A1(I1074), .A2(W8215), .ZN(O1668));
  NANDX1 G25347 (.A1(W1718), .A2(I1152), .ZN(W4504));
  NANDX1 G25348 (.A1(W5914), .A2(W5314), .ZN(W8145));
  NANDX1 G25349 (.A1(W2948), .A2(I1716), .ZN(W8143));
  NANDX1 G25350 (.A1(I881), .A2(W1985), .ZN(W4511));
  NANDX1 G25351 (.A1(W17975), .A2(W15672), .ZN(W18875));
  NANDX1 G25352 (.A1(I331), .A2(W1187), .ZN(W13185));
  NANDX1 G25353 (.A1(W257), .A2(W7609), .ZN(W13180));
  NANDX1 G25354 (.A1(W13491), .A2(W3321), .ZN(W18872));
  NANDX1 G25355 (.A1(W11164), .A2(W16930), .ZN(O1665));
  NANDX1 G25356 (.A1(W9876), .A2(W11238), .ZN(O1664));
  NANDX1 G25357 (.A1(I435), .A2(I1974), .ZN(W4516));
  NANDX1 G25358 (.A1(W16543), .A2(W3432), .ZN(W18865));
  NANDX1 G25359 (.A1(W4488), .A2(W1390), .ZN(O213));
  NANDX1 G25360 (.A1(W7926), .A2(W860), .ZN(W8139));
  NANDX1 G25361 (.A1(W1553), .A2(W2688), .ZN(W8137));
  NANDX1 G25362 (.A1(W6833), .A2(W6573), .ZN(W8153));
  NANDX1 G25363 (.A1(W2935), .A2(W1063), .ZN(O1674));
  NANDX1 G25364 (.A1(W539), .A2(W1791), .ZN(W4487));
  NANDX1 G25365 (.A1(W3505), .A2(W2937), .ZN(W4489));
  NANDX1 G25366 (.A1(W11490), .A2(W5510), .ZN(W13171));
  NANDX1 G25367 (.A1(W18745), .A2(W2568), .ZN(W18896));
  NANDX1 G25368 (.A1(W2332), .A2(W3952), .ZN(W4491));
  NANDX1 G25369 (.A1(W10043), .A2(I288), .ZN(W18893));
  NANDX1 G25370 (.A1(W1145), .A2(W2896), .ZN(W4493));
  NANDX1 G25371 (.A1(W845), .A2(W4012), .ZN(W4525));
  NANDX1 G25372 (.A1(W2509), .A2(I1214), .ZN(O58));
  NANDX1 G25373 (.A1(W3319), .A2(W10495), .ZN(W13173));
  NANDX1 G25374 (.A1(W2514), .A2(I744), .ZN(W4496));
  NANDX1 G25375 (.A1(W922), .A2(W8221), .ZN(W13176));
  NANDX1 G25376 (.A1(W7266), .A2(I301), .ZN(W8149));
  NANDX1 G25377 (.A1(W2607), .A2(W3962), .ZN(O1671));
  NANDX1 G25378 (.A1(W865), .A2(I144), .ZN(W8148));
  NANDX1 G25379 (.A1(W11643), .A2(W3775), .ZN(W13178));
  NANDX1 G25380 (.A1(W17526), .A2(W12643), .ZN(O1655));
  NANDX1 G25381 (.A1(W7151), .A2(W4810), .ZN(W8133));
  NANDX1 G25382 (.A1(I1603), .A2(W5038), .ZN(W18837));
  NANDX1 G25383 (.A1(W11048), .A2(W12657), .ZN(W13203));
  NANDX1 G25384 (.A1(W108), .A2(W2320), .ZN(W13205));
  NANDX1 G25385 (.A1(W16923), .A2(I1807), .ZN(O1656));
  NANDX1 G25386 (.A1(I1563), .A2(W9612), .ZN(W13208));
  NANDX1 G25387 (.A1(W11438), .A2(W5686), .ZN(W13209));
  NANDX1 G25388 (.A1(I563), .A2(W11731), .ZN(W13210));
  NANDX1 G25389 (.A1(W2323), .A2(W1158), .ZN(W4543));
  NANDX1 G25390 (.A1(W14935), .A2(W15174), .ZN(W18840));
  NANDX1 G25391 (.A1(I1232), .A2(W1300), .ZN(W4545));
  NANDX1 G25392 (.A1(W1727), .A2(W7266), .ZN(W18829));
  NANDX1 G25393 (.A1(W4947), .A2(I1403), .ZN(W18827));
  NANDX1 G25394 (.A1(W736), .A2(W4457), .ZN(W4548));
  NANDX1 G25395 (.A1(W4968), .A2(W3502), .ZN(W13217));
  NANDX1 G25396 (.A1(I1788), .A2(W349), .ZN(W18824));
  NANDX1 G25397 (.A1(W837), .A2(W18119), .ZN(W18822));
  NANDX1 G25398 (.A1(I1352), .A2(W4772), .ZN(W13219));
  NANDX1 G25399 (.A1(W2932), .A2(W2214), .ZN(W4532));
  NANDX1 G25400 (.A1(I415), .A2(W266), .ZN(W18856));
  NANDX1 G25401 (.A1(W5901), .A2(W2939), .ZN(W13192));
  NANDX1 G25402 (.A1(W7962), .A2(W5221), .ZN(W18852));
  NANDX1 G25403 (.A1(W2735), .A2(W2007), .ZN(W4529));
  NANDX1 G25404 (.A1(W3528), .A2(I117), .ZN(W13194));
  NANDX1 G25405 (.A1(W16535), .A2(W3845), .ZN(W18850));
  NANDX1 G25406 (.A1(I1588), .A2(I728), .ZN(W13195));
  NANDX1 G25407 (.A1(W10964), .A2(W3797), .ZN(W18847));
  NANDX1 G25408 (.A1(W6586), .A2(W4267), .ZN(W13168));
  NANDX1 G25409 (.A1(W2738), .A2(W12028), .ZN(W13196));
  NANDX1 G25410 (.A1(I521), .A2(W385), .ZN(W4535));
  NANDX1 G25411 (.A1(W17712), .A2(W16000), .ZN(W18844));
  NANDX1 G25412 (.A1(W18483), .A2(I609), .ZN(W18842));
  NANDX1 G25413 (.A1(W3954), .A2(W1986), .ZN(W4537));
  NANDX1 G25414 (.A1(W11297), .A2(W10551), .ZN(W13198));
  NANDX1 G25415 (.A1(W1672), .A2(I1473), .ZN(W4538));
  NANDX1 G25416 (.A1(W42), .A2(W1866), .ZN(W4539));
  NANDX1 G25417 (.A1(W2307), .A2(W12460), .ZN(W18954));
  NANDX1 G25418 (.A1(W9247), .A2(W11368), .ZN(W13148));
  NANDX1 G25419 (.A1(W10626), .A2(I1878), .ZN(W18963));
  NANDX1 G25420 (.A1(W11209), .A2(W8797), .ZN(W18962));
  NANDX1 G25421 (.A1(W7601), .A2(I1448), .ZN(W18959));
  NANDX1 G25422 (.A1(W14961), .A2(I711), .ZN(W18957));
  NANDX1 G25423 (.A1(W4559), .A2(W1108), .ZN(W8180));
  NANDX1 G25424 (.A1(I1957), .A2(W1700), .ZN(W4435));
  NANDX1 G25425 (.A1(W9675), .A2(W8813), .ZN(W18956));
  NANDX1 G25426 (.A1(I1956), .A2(W2476), .ZN(W4436));
  NANDX1 G25427 (.A1(W7071), .A2(W12810), .ZN(W13146));
  NANDX1 G25428 (.A1(I259), .A2(I686), .ZN(W4437));
  NANDX1 G25429 (.A1(W6984), .A2(W5294), .ZN(W8179));
  NANDX1 G25430 (.A1(W7254), .A2(I1732), .ZN(W18952));
  NANDX1 G25431 (.A1(W2318), .A2(W7544), .ZN(W13154));
  NANDX1 G25432 (.A1(I1296), .A2(W1149), .ZN(W4444));
  NANDX1 G25433 (.A1(W2222), .A2(W4901), .ZN(W13156));
  NANDX1 G25434 (.A1(W3149), .A2(W1946), .ZN(W4449));
  NANDX1 G25435 (.A1(W4976), .A2(W16129), .ZN(O1679));
  NANDX1 G25436 (.A1(W1374), .A2(W3706), .ZN(W4421));
  NANDX1 G25437 (.A1(W5179), .A2(W3920), .ZN(W8187));
  NANDX1 G25438 (.A1(W10333), .A2(W1531), .ZN(O1685));
  NANDX1 G25439 (.A1(W11208), .A2(W8858), .ZN(W13137));
  NANDX1 G25440 (.A1(W2868), .A2(W1495), .ZN(W13138));
  NANDX1 G25441 (.A1(W913), .A2(W6031), .ZN(W18980));
  NANDX1 G25442 (.A1(W8134), .A2(W12520), .ZN(W18979));
  NANDX1 G25443 (.A1(I1538), .A2(I548), .ZN(W8185));
  NANDX1 G25444 (.A1(W4017), .A2(W149), .ZN(W4420));
  NANDX1 G25445 (.A1(W2283), .A2(W2497), .ZN(W4450));
  NANDX1 G25446 (.A1(W3818), .A2(W1298), .ZN(W4422));
  NANDX1 G25447 (.A1(W3970), .A2(W4293), .ZN(W4424));
  NANDX1 G25448 (.A1(W1430), .A2(W6315), .ZN(W8184));
  NANDX1 G25449 (.A1(W3479), .A2(W2019), .ZN(W8183));
  NANDX1 G25450 (.A1(W4807), .A2(W15668), .ZN(O1683));
  NANDX1 G25451 (.A1(W8271), .A2(I1263), .ZN(O1682));
  NANDX1 G25452 (.A1(I964), .A2(W10624), .ZN(W13143));
  NANDX1 G25453 (.A1(W16338), .A2(W11571), .ZN(O1681));
  NANDX1 G25454 (.A1(W14210), .A2(W7348), .ZN(W18910));
  NANDX1 G25455 (.A1(W2883), .A2(I1998), .ZN(W4465));
  NANDX1 G25456 (.A1(W11675), .A2(W1453), .ZN(W18923));
  NANDX1 G25457 (.A1(W6238), .A2(W7768), .ZN(W18920));
  NANDX1 G25458 (.A1(W246), .A2(W2257), .ZN(W4467));
  NANDX1 G25459 (.A1(W7102), .A2(W7031), .ZN(W18916));
  NANDX1 G25460 (.A1(W3990), .A2(W102), .ZN(W4468));
  NANDX1 G25461 (.A1(W3250), .A2(W6996), .ZN(W8168));
  NANDX1 G25462 (.A1(W3257), .A2(W4408), .ZN(W4478));
  NANDX1 G25463 (.A1(W910), .A2(W3083), .ZN(W4462));
  NANDX1 G25464 (.A1(W6003), .A2(W1127), .ZN(W18909));
  NANDX1 G25465 (.A1(W1512), .A2(W3034), .ZN(W8160));
  NANDX1 G25466 (.A1(W10698), .A2(W12457), .ZN(W18907));
  NANDX1 G25467 (.A1(W5920), .A2(W8040), .ZN(W8158));
  NANDX1 G25468 (.A1(W1381), .A2(W9901), .ZN(W13166));
  NANDX1 G25469 (.A1(I64), .A2(W1888), .ZN(W4483));
  NANDX1 G25470 (.A1(W2547), .A2(W4197), .ZN(W4485));
  NANDX1 G25471 (.A1(I1178), .A2(W2025), .ZN(W13167));
  NANDX1 G25472 (.A1(W12987), .A2(W3819), .ZN(W18932));
  NANDX1 G25473 (.A1(W4215), .A2(W2069), .ZN(W18944));
  NANDX1 G25474 (.A1(I966), .A2(W5663), .ZN(W8176));
  NANDX1 G25475 (.A1(W10535), .A2(W1150), .ZN(W18942));
  NANDX1 G25476 (.A1(W6287), .A2(W17407), .ZN(W18941));
  NANDX1 G25477 (.A1(W878), .A2(W842), .ZN(W8171));
  NANDX1 G25478 (.A1(W16980), .A2(W2840), .ZN(W18937));
  NANDX1 G25479 (.A1(W3757), .A2(W3162), .ZN(W4456));
  NANDX1 G25480 (.A1(W3881), .A2(W5266), .ZN(W13161));
  NANDX1 G25481 (.A1(W6820), .A2(W2344), .ZN(W13220));
  NANDX1 G25482 (.A1(W5953), .A2(W830), .ZN(W18931));
  NANDX1 G25483 (.A1(W17260), .A2(I23), .ZN(W18930));
  NANDX1 G25484 (.A1(W4453), .A2(W4999), .ZN(W8170));
  NANDX1 G25485 (.A1(W1443), .A2(W4256), .ZN(W4459));
  NANDX1 G25486 (.A1(W12912), .A2(I726), .ZN(W18928));
  NANDX1 G25487 (.A1(I1028), .A2(W1364), .ZN(W18927));
  NANDX1 G25488 (.A1(I433), .A2(I1536), .ZN(W4460));
  NANDX1 G25489 (.A1(W10140), .A2(W17874), .ZN(O1678));
  NANDX1 G25490 (.A1(W2815), .A2(W592), .ZN(W13281));
  NANDX1 G25491 (.A1(W18616), .A2(W12427), .ZN(O1624));
  NANDX1 G25492 (.A1(W3262), .A2(W286), .ZN(W4633));
  NANDX1 G25493 (.A1(W3659), .A2(I117), .ZN(W18696));
  NANDX1 G25494 (.A1(W7244), .A2(W7023), .ZN(W8105));
  NANDX1 G25495 (.A1(W17246), .A2(W13125), .ZN(O1623));
  NANDX1 G25496 (.A1(W725), .A2(W2257), .ZN(W8099));
  NANDX1 G25497 (.A1(I754), .A2(W2694), .ZN(W4634));
  NANDX1 G25498 (.A1(W519), .A2(W12302), .ZN(O1622));
  NANDX1 G25499 (.A1(W2790), .A2(W3568), .ZN(W13278));
  NANDX1 G25500 (.A1(W11003), .A2(W11167), .ZN(W13273));
  NANDX1 G25501 (.A1(W10970), .A2(W4101), .ZN(W13282));
  NANDX1 G25502 (.A1(W11841), .A2(W18330), .ZN(W18686));
  NANDX1 G25503 (.A1(I895), .A2(I1439), .ZN(O212));
  NANDX1 G25504 (.A1(W8070), .A2(W12511), .ZN(O1620));
  NANDX1 G25505 (.A1(W743), .A2(W16927), .ZN(W18680));
  NANDX1 G25506 (.A1(W15739), .A2(W12087), .ZN(W18678));
  NANDX1 G25507 (.A1(W2404), .A2(W10553), .ZN(W18676));
  NANDX1 G25508 (.A1(W18303), .A2(W3942), .ZN(W18675));
  NANDX1 G25509 (.A1(W5906), .A2(W10110), .ZN(W18709));
  NANDX1 G25510 (.A1(W2533), .A2(W1701), .ZN(W18721));
  NANDX1 G25511 (.A1(I85), .A2(W1079), .ZN(W18716));
  NANDX1 G25512 (.A1(I46), .A2(W7626), .ZN(W8109));
  NANDX1 G25513 (.A1(W4740), .A2(W15522), .ZN(W18713));
  NANDX1 G25514 (.A1(I1482), .A2(W4632), .ZN(W13260));
  NANDX1 G25515 (.A1(W5325), .A2(W11985), .ZN(W13261));
  NANDX1 G25516 (.A1(W703), .A2(W2651), .ZN(W4620));
  NANDX1 G25517 (.A1(W11578), .A2(W6006), .ZN(O721));
  NANDX1 G25518 (.A1(W8214), .A2(W10141), .ZN(O1618));
  NANDX1 G25519 (.A1(W11452), .A2(W10363), .ZN(W13266));
  NANDX1 G25520 (.A1(I407), .A2(I1029), .ZN(W4627));
  NANDX1 G25521 (.A1(W2760), .A2(W5819), .ZN(W8106));
  NANDX1 G25522 (.A1(I354), .A2(I844), .ZN(W4630));
  NANDX1 G25523 (.A1(W6172), .A2(W16594), .ZN(W18703));
  NANDX1 G25524 (.A1(W6031), .A2(W12049), .ZN(W13272));
  NANDX1 G25525 (.A1(W9086), .A2(W16284), .ZN(W18702));
  NANDX1 G25526 (.A1(W15807), .A2(W9944), .ZN(W18700));
  NANDX1 G25527 (.A1(W16815), .A2(W4203), .ZN(W18640));
  NANDX1 G25528 (.A1(W3131), .A2(W8022), .ZN(W8079));
  NANDX1 G25529 (.A1(W534), .A2(W9768), .ZN(W13303));
  NANDX1 G25530 (.A1(W13180), .A2(W1968), .ZN(O725));
  NANDX1 G25531 (.A1(W17785), .A2(W17400), .ZN(O1611));
  NANDX1 G25532 (.A1(W9630), .A2(W10786), .ZN(W13308));
  NANDX1 G25533 (.A1(W1569), .A2(W14374), .ZN(O1610));
  NANDX1 G25534 (.A1(W14731), .A2(W5690), .ZN(O1609));
  NANDX1 G25535 (.A1(W1478), .A2(W16633), .ZN(O1608));
  NANDX1 G25536 (.A1(W9362), .A2(W2840), .ZN(O1613));
  NANDX1 G25537 (.A1(W2155), .A2(I977), .ZN(W4663));
  NANDX1 G25538 (.A1(W1901), .A2(W6525), .ZN(W18638));
  NANDX1 G25539 (.A1(I1498), .A2(W3924), .ZN(W8078));
  NANDX1 G25540 (.A1(W1080), .A2(W5725), .ZN(W8076));
  NANDX1 G25541 (.A1(W2411), .A2(W784), .ZN(W4668));
  NANDX1 G25542 (.A1(W1293), .A2(W8340), .ZN(W18633));
  NANDX1 G25543 (.A1(W12366), .A2(W4961), .ZN(W13310));
  NANDX1 G25544 (.A1(I238), .A2(W310), .ZN(W8074));
  NANDX1 G25545 (.A1(W2664), .A2(W3112), .ZN(W8089));
  NANDX1 G25546 (.A1(W16447), .A2(W8152), .ZN(W18673));
  NANDX1 G25547 (.A1(W4453), .A2(W3742), .ZN(W4646));
  NANDX1 G25548 (.A1(W3929), .A2(W1305), .ZN(W13289));
  NANDX1 G25549 (.A1(W12198), .A2(W4941), .ZN(W13290));
  NANDX1 G25550 (.A1(W12024), .A2(W7660), .ZN(W13292));
  NANDX1 G25551 (.A1(W3918), .A2(W2417), .ZN(W4649));
  NANDX1 G25552 (.A1(W6511), .A2(W9802), .ZN(W18669));
  NANDX1 G25553 (.A1(W11974), .A2(W17800), .ZN(W18667));
  NANDX1 G25554 (.A1(W11723), .A2(W10438), .ZN(W13259));
  NANDX1 G25555 (.A1(W12354), .A2(W890), .ZN(O1617));
  NANDX1 G25556 (.A1(W4322), .A2(W1365), .ZN(W18662));
  NANDX1 G25557 (.A1(W18447), .A2(W8646), .ZN(W18661));
  NANDX1 G25558 (.A1(W4745), .A2(I793), .ZN(W8082));
  NANDX1 G25559 (.A1(W2966), .A2(W84), .ZN(W4656));
  NANDX1 G25560 (.A1(W11180), .A2(W12928), .ZN(W18652));
  NANDX1 G25561 (.A1(I1848), .A2(W17550), .ZN(O1615));
  NANDX1 G25562 (.A1(W12449), .A2(W4796), .ZN(W18650));
  NANDX1 G25563 (.A1(W1482), .A2(W6816), .ZN(W13235));
  NANDX1 G25564 (.A1(I811), .A2(W8987), .ZN(W13228));
  NANDX1 G25565 (.A1(I1912), .A2(W11), .ZN(W8124));
  NANDX1 G25566 (.A1(W3372), .A2(I600), .ZN(O714));
  NANDX1 G25567 (.A1(W13015), .A2(W15281), .ZN(O1647));
  NANDX1 G25568 (.A1(W4477), .A2(I583), .ZN(W4574));
  NANDX1 G25569 (.A1(W17079), .A2(W4510), .ZN(O1646));
  NANDX1 G25570 (.A1(W3827), .A2(I942), .ZN(W4576));
  NANDX1 G25571 (.A1(W6359), .A2(W18492), .ZN(W18780));
  NANDX1 G25572 (.A1(W12637), .A2(W15350), .ZN(W18778));
  NANDX1 G25573 (.A1(W3294), .A2(W7697), .ZN(W18793));
  NANDX1 G25574 (.A1(W12830), .A2(W4688), .ZN(W18777));
  NANDX1 G25575 (.A1(W199), .A2(W1056), .ZN(W8120));
  NANDX1 G25576 (.A1(W4152), .A2(W2847), .ZN(W4582));
  NANDX1 G25577 (.A1(W13071), .A2(W13221), .ZN(O1643));
  NANDX1 G25578 (.A1(W10482), .A2(I1190), .ZN(W13240));
  NANDX1 G25579 (.A1(W2371), .A2(W1740), .ZN(W4584));
  NANDX1 G25580 (.A1(W3873), .A2(W5925), .ZN(W13242));
  NANDX1 G25581 (.A1(W7912), .A2(W3662), .ZN(W13245));
  NANDX1 G25582 (.A1(W15168), .A2(W12361), .ZN(O1650));
  NANDX1 G25583 (.A1(W2134), .A2(W634), .ZN(W4556));
  NANDX1 G25584 (.A1(W132), .A2(W4345), .ZN(W4558));
  NANDX1 G25585 (.A1(W2201), .A2(W154), .ZN(W18816));
  NANDX1 G25586 (.A1(W11575), .A2(W1527), .ZN(W13222));
  NANDX1 G25587 (.A1(W2446), .A2(W6459), .ZN(W13225));
  NANDX1 G25588 (.A1(W5529), .A2(I1246), .ZN(W8127));
  NANDX1 G25589 (.A1(W10442), .A2(W7638), .ZN(W18809));
  NANDX1 G25590 (.A1(W16148), .A2(W8198), .ZN(W18804));
  NANDX1 G25591 (.A1(I744), .A2(I437), .ZN(W18768));
  NANDX1 G25592 (.A1(W2247), .A2(I967), .ZN(W4562));
  NANDX1 G25593 (.A1(W4223), .A2(W2148), .ZN(O60));
  NANDX1 G25594 (.A1(I74), .A2(W17126), .ZN(W18801));
  NANDX1 G25595 (.A1(W3694), .A2(W526), .ZN(W13227));
  NANDX1 G25596 (.A1(I1194), .A2(I832), .ZN(W4567));
  NANDX1 G25597 (.A1(W540), .A2(W14803), .ZN(W18795));
  NANDX1 G25598 (.A1(W1043), .A2(W17222), .ZN(W18794));
  NANDX1 G25599 (.A1(W3794), .A2(I1247), .ZN(W8126));
  NANDX1 G25600 (.A1(W5744), .A2(W4924), .ZN(W18736));
  NANDX1 G25601 (.A1(W14410), .A2(W7118), .ZN(W18745));
  NANDX1 G25602 (.A1(W6168), .A2(W13387), .ZN(W18744));
  NANDX1 G25603 (.A1(W1042), .A2(W574), .ZN(W4598));
  NANDX1 G25604 (.A1(W840), .A2(I1409), .ZN(W8113));
  NANDX1 G25605 (.A1(W3855), .A2(W532), .ZN(W4601));
  NANDX1 G25606 (.A1(W3635), .A2(W1594), .ZN(O1632));
  NANDX1 G25607 (.A1(I1180), .A2(I1157), .ZN(W4606));
  NANDX1 G25608 (.A1(I1190), .A2(W238), .ZN(W8112));
  NANDX1 G25609 (.A1(W4341), .A2(W6860), .ZN(W8116));
  NANDX1 G25610 (.A1(W16086), .A2(W2201), .ZN(W18734));
  NANDX1 G25611 (.A1(W11426), .A2(W8391), .ZN(O1631));
  NANDX1 G25612 (.A1(I1004), .A2(W555), .ZN(W4612));
  NANDX1 G25613 (.A1(W1460), .A2(W8224), .ZN(W18729));
  NANDX1 G25614 (.A1(W9159), .A2(W7014), .ZN(W13256));
  NANDX1 G25615 (.A1(W10990), .A2(W5904), .ZN(W18725));
  NANDX1 G25616 (.A1(W2250), .A2(W5637), .ZN(W13257));
  NANDX1 G25617 (.A1(W1507), .A2(W4885), .ZN(O1630));
  NANDX1 G25618 (.A1(W5469), .A2(W8048), .ZN(O1638));
  NANDX1 G25619 (.A1(W9442), .A2(W14066), .ZN(W18767));
  NANDX1 G25620 (.A1(I629), .A2(W7657), .ZN(W8119));
  NANDX1 G25621 (.A1(W6071), .A2(W17867), .ZN(O1639));
  NANDX1 G25622 (.A1(W9797), .A2(W12910), .ZN(W18763));
  NANDX1 G25623 (.A1(I432), .A2(W3734), .ZN(W4592));
  NANDX1 G25624 (.A1(W18029), .A2(W8815), .ZN(W18760));
  NANDX1 G25625 (.A1(W8063), .A2(I1612), .ZN(W13248));
  NANDX1 G25626 (.A1(W4610), .A2(W14729), .ZN(W18759));
  NANDX1 G25627 (.A1(I1042), .A2(W7654), .ZN(W13132));
  NANDX1 G25628 (.A1(I782), .A2(W3645), .ZN(W4593));
  NANDX1 G25629 (.A1(W5173), .A2(I1852), .ZN(W13249));
  NANDX1 G25630 (.A1(I1701), .A2(W2697), .ZN(W8118));
  NANDX1 G25631 (.A1(W3044), .A2(W1618), .ZN(O1635));
  NANDX1 G25632 (.A1(W7833), .A2(W228), .ZN(W18752));
  NANDX1 G25633 (.A1(W15570), .A2(W8389), .ZN(O1634));
  NANDX1 G25634 (.A1(W11808), .A2(W17045), .ZN(W18748));
  NANDX1 G25635 (.A1(W5159), .A2(W1037), .ZN(W13251));
  NANDX1 G25636 (.A1(W3903), .A2(W1109), .ZN(W4248));
  NANDX1 G25637 (.A1(W3616), .A2(W3395), .ZN(W4244));
  NANDX1 G25638 (.A1(W1718), .A2(W10479), .ZN(W13050));
  NANDX1 G25639 (.A1(I752), .A2(W2164), .ZN(W4245));
  NANDX1 G25640 (.A1(W1948), .A2(I604), .ZN(W8252));
  NANDX1 G25641 (.A1(W3064), .A2(W5713), .ZN(W13052));
  NANDX1 G25642 (.A1(W16658), .A2(W5947), .ZN(W19213));
  NANDX1 G25643 (.A1(W328), .A2(W6769), .ZN(W13053));
  NANDX1 G25644 (.A1(W11470), .A2(W1468), .ZN(W19208));
  NANDX1 G25645 (.A1(I1981), .A2(W3879), .ZN(W4246));
  NANDX1 G25646 (.A1(W11783), .A2(W8193), .ZN(W19217));
  NANDX1 G25647 (.A1(W7312), .A2(W7203), .ZN(W13054));
  NANDX1 G25648 (.A1(W3496), .A2(W8237), .ZN(W19203));
  NANDX1 G25649 (.A1(W5605), .A2(W7847), .ZN(W19202));
  NANDX1 G25650 (.A1(W1104), .A2(W4642), .ZN(W19201));
  NANDX1 G25651 (.A1(W4516), .A2(W12015), .ZN(W19200));
  NANDX1 G25652 (.A1(W9316), .A2(W571), .ZN(W13055));
  NANDX1 G25653 (.A1(W7503), .A2(W3325), .ZN(W19198));
  NANDX1 G25654 (.A1(I8), .A2(I1679), .ZN(O218));
  NANDX1 G25655 (.A1(I1878), .A2(W1522), .ZN(O683));
  NANDX1 G25656 (.A1(W9829), .A2(W15851), .ZN(O1730));
  NANDX1 G25657 (.A1(W641), .A2(W10881), .ZN(W19235));
  NANDX1 G25658 (.A1(W3707), .A2(W5113), .ZN(W8260));
  NANDX1 G25659 (.A1(W2081), .A2(W2528), .ZN(W8258));
  NANDX1 G25660 (.A1(W8740), .A2(W2955), .ZN(W19230));
  NANDX1 G25661 (.A1(W7083), .A2(W10305), .ZN(W19227));
  NANDX1 G25662 (.A1(W18587), .A2(W4484), .ZN(W19226));
  NANDX1 G25663 (.A1(W3884), .A2(W5501), .ZN(O682));
  NANDX1 G25664 (.A1(W3767), .A2(W4270), .ZN(O687));
  NANDX1 G25665 (.A1(W12832), .A2(W10662), .ZN(W13040));
  NANDX1 G25666 (.A1(W6864), .A2(W4760), .ZN(O1728));
  NANDX1 G25667 (.A1(W7628), .A2(W2419), .ZN(O684));
  NANDX1 G25668 (.A1(W8533), .A2(W10801), .ZN(W13044));
  NANDX1 G25669 (.A1(W13248), .A2(W17952), .ZN(W19220));
  NANDX1 G25670 (.A1(W98), .A2(W948), .ZN(W4242));
  NANDX1 G25671 (.A1(W12417), .A2(W2240), .ZN(O1727));
  NANDX1 G25672 (.A1(W3934), .A2(W3703), .ZN(W13048));
  NANDX1 G25673 (.A1(W2938), .A2(W3340), .ZN(W13071));
  NANDX1 G25674 (.A1(W3880), .A2(W2065), .ZN(W8244));
  NANDX1 G25675 (.A1(W1550), .A2(W7586), .ZN(W13067));
  NANDX1 G25676 (.A1(W6855), .A2(W4841), .ZN(W19180));
  NANDX1 G25677 (.A1(W17840), .A2(W7394), .ZN(W19177));
  NANDX1 G25678 (.A1(W4537), .A2(W9418), .ZN(W19175));
  NANDX1 G25679 (.A1(W4176), .A2(W4019), .ZN(W19173));
  NANDX1 G25680 (.A1(W5454), .A2(W7690), .ZN(O689));
  NANDX1 G25681 (.A1(I339), .A2(W8025), .ZN(W13070));
  NANDX1 G25682 (.A1(I600), .A2(W1845), .ZN(W4270));
  NANDX1 G25683 (.A1(W9085), .A2(W1979), .ZN(W19170));
  NANDX1 G25684 (.A1(W8382), .A2(W18947), .ZN(O1721));
  NANDX1 G25685 (.A1(W296), .A2(W253), .ZN(W4276));
  NANDX1 G25686 (.A1(I248), .A2(W14649), .ZN(O1720));
  NANDX1 G25687 (.A1(I1341), .A2(W1584), .ZN(W4277));
  NANDX1 G25688 (.A1(W51), .A2(I1759), .ZN(W8243));
  NANDX1 G25689 (.A1(W1486), .A2(W11309), .ZN(W13074));
  NANDX1 G25690 (.A1(W11875), .A2(W3414), .ZN(O1719));
  NANDX1 G25691 (.A1(I1903), .A2(W318), .ZN(W4261));
  NANDX1 G25692 (.A1(W12056), .A2(I1826), .ZN(W19196));
  NANDX1 G25693 (.A1(I445), .A2(W2655), .ZN(W4251));
  NANDX1 G25694 (.A1(W4157), .A2(W3656), .ZN(W4252));
  NANDX1 G25695 (.A1(W8868), .A2(W10504), .ZN(W13058));
  NANDX1 G25696 (.A1(W1226), .A2(I3), .ZN(W8247));
  NANDX1 G25697 (.A1(W568), .A2(W2565), .ZN(W4256));
  NANDX1 G25698 (.A1(W4056), .A2(W2491), .ZN(W4257));
  NANDX1 G25699 (.A1(W3805), .A2(W1487), .ZN(W4258));
  NANDX1 G25700 (.A1(W6944), .A2(W10591), .ZN(W13033));
  NANDX1 G25701 (.A1(W11135), .A2(W11878), .ZN(W13059));
  NANDX1 G25702 (.A1(W12096), .A2(W13020), .ZN(W19190));
  NANDX1 G25703 (.A1(I354), .A2(I135), .ZN(W4264));
  NANDX1 G25704 (.A1(W3709), .A2(W11491), .ZN(W19187));
  NANDX1 G25705 (.A1(W17615), .A2(W12459), .ZN(W19186));
  NANDX1 G25706 (.A1(W5210), .A2(W10098), .ZN(W13064));
  NANDX1 G25707 (.A1(I659), .A2(W2526), .ZN(W4268));
  NANDX1 G25708 (.A1(W3322), .A2(W3271), .ZN(W4269));
  NANDX1 G25709 (.A1(W9585), .A2(W8915), .ZN(W12990));
  NANDX1 G25710 (.A1(W2970), .A2(W2056), .ZN(W4167));
  NANDX1 G25711 (.A1(W16573), .A2(W17031), .ZN(W19286));
  NANDX1 G25712 (.A1(W13755), .A2(W1238), .ZN(W19285));
  NANDX1 G25713 (.A1(W6112), .A2(W12448), .ZN(O1741));
  NANDX1 G25714 (.A1(W10385), .A2(W9506), .ZN(W19281));
  NANDX1 G25715 (.A1(I1936), .A2(W5572), .ZN(W12987));
  NANDX1 G25716 (.A1(W7423), .A2(W4283), .ZN(W8288));
  NANDX1 G25717 (.A1(W2279), .A2(W10454), .ZN(W19280));
  NANDX1 G25718 (.A1(W8641), .A2(W6126), .ZN(W19279));
  NANDX1 G25719 (.A1(W18594), .A2(W356), .ZN(W19288));
  NANDX1 G25720 (.A1(W2943), .A2(W95), .ZN(W4177));
  NANDX1 G25721 (.A1(W7111), .A2(W5651), .ZN(W12996));
  NANDX1 G25722 (.A1(W1973), .A2(W1468), .ZN(W4179));
  NANDX1 G25723 (.A1(I372), .A2(W11287), .ZN(W12997));
  NANDX1 G25724 (.A1(W6769), .A2(W8525), .ZN(W12998));
  NANDX1 G25725 (.A1(W1891), .A2(W1941), .ZN(W4182));
  NANDX1 G25726 (.A1(W1801), .A2(W2434), .ZN(W8285));
  NANDX1 G25727 (.A1(W2939), .A2(W6227), .ZN(O1738));
  NANDX1 G25728 (.A1(W3716), .A2(W14286), .ZN(W19301));
  NANDX1 G25729 (.A1(I370), .A2(W2956), .ZN(W8292));
  NANDX1 G25730 (.A1(W7029), .A2(W11738), .ZN(W12982));
  NANDX1 G25731 (.A1(W157), .A2(W1020), .ZN(W4156));
  NANDX1 G25732 (.A1(W1280), .A2(W282), .ZN(W4157));
  NANDX1 G25733 (.A1(W1073), .A2(W2306), .ZN(W4160));
  NANDX1 G25734 (.A1(I1552), .A2(I1102), .ZN(W4161));
  NANDX1 G25735 (.A1(W4693), .A2(I140), .ZN(W8290));
  NANDX1 G25736 (.A1(W698), .A2(W18883), .ZN(W19303));
  NANDX1 G25737 (.A1(W728), .A2(W8554), .ZN(W13000));
  NANDX1 G25738 (.A1(W19234), .A2(W16961), .ZN(W19300));
  NANDX1 G25739 (.A1(W9564), .A2(W13097), .ZN(W19294));
  NANDX1 G25740 (.A1(W6821), .A2(W11818), .ZN(W19293));
  NANDX1 G25741 (.A1(I917), .A2(I315), .ZN(W4163));
  NANDX1 G25742 (.A1(W16327), .A2(W10522), .ZN(W19291));
  NANDX1 G25743 (.A1(W3924), .A2(I1425), .ZN(W4165));
  NANDX1 G25744 (.A1(W7915), .A2(I930), .ZN(W19290));
  NANDX1 G25745 (.A1(W3395), .A2(W2265), .ZN(W8289));
  NANDX1 G25746 (.A1(I44), .A2(W385), .ZN(W19245));
  NANDX1 G25747 (.A1(W2870), .A2(I431), .ZN(W4212));
  NANDX1 G25748 (.A1(W10121), .A2(W10272), .ZN(W19248));
  NANDX1 G25749 (.A1(W10591), .A2(W9754), .ZN(W19247));
  NANDX1 G25750 (.A1(W7240), .A2(W2968), .ZN(W8267));
  NANDX1 G25751 (.A1(W994), .A2(W773), .ZN(W4218));
  NANDX1 G25752 (.A1(I1429), .A2(W1180), .ZN(W4220));
  NANDX1 G25753 (.A1(W6986), .A2(W3425), .ZN(W8263));
  NANDX1 G25754 (.A1(W1918), .A2(W3534), .ZN(W4223));
  NANDX1 G25755 (.A1(W12469), .A2(I1568), .ZN(W13021));
  NANDX1 G25756 (.A1(W1875), .A2(W6453), .ZN(W8261));
  NANDX1 G25757 (.A1(W13789), .A2(W4377), .ZN(W19243));
  NANDX1 G25758 (.A1(I1590), .A2(W10997), .ZN(W13025));
  NANDX1 G25759 (.A1(W6332), .A2(W12476), .ZN(O1732));
  NANDX1 G25760 (.A1(W10824), .A2(I1500), .ZN(W13026));
  NANDX1 G25761 (.A1(W9438), .A2(W9391), .ZN(W19240));
  NANDX1 G25762 (.A1(W8478), .A2(I1992), .ZN(W13028));
  NANDX1 G25763 (.A1(W10548), .A2(W8956), .ZN(W13032));
  NANDX1 G25764 (.A1(W5757), .A2(W8154), .ZN(W13011));
  NANDX1 G25765 (.A1(I1622), .A2(W1360), .ZN(W19269));
  NANDX1 G25766 (.A1(W6970), .A2(W5622), .ZN(W13001));
  NANDX1 G25767 (.A1(W11561), .A2(W8235), .ZN(W19265));
  NANDX1 G25768 (.A1(W1594), .A2(W1081), .ZN(W4189));
  NANDX1 G25769 (.A1(W5031), .A2(W2279), .ZN(W8281));
  NANDX1 G25770 (.A1(W12175), .A2(W16367), .ZN(W19263));
  NANDX1 G25771 (.A1(W3761), .A2(W3131), .ZN(W8279));
  NANDX1 G25772 (.A1(W2796), .A2(W1964), .ZN(W4205));
  NANDX1 G25773 (.A1(W2244), .A2(W6768), .ZN(O216));
  NANDX1 G25774 (.A1(W1207), .A2(I1168), .ZN(W4207));
  NANDX1 G25775 (.A1(W16831), .A2(W7729), .ZN(O1736));
  NANDX1 G25776 (.A1(W2682), .A2(W2848), .ZN(W4208));
  NANDX1 G25777 (.A1(W16601), .A2(W14064), .ZN(W19257));
  NANDX1 G25778 (.A1(W7364), .A2(W3903), .ZN(W8277));
  NANDX1 G25779 (.A1(W3429), .A2(W2271), .ZN(W4209));
  NANDX1 G25780 (.A1(W11889), .A2(W3060), .ZN(W13019));
  NANDX1 G25781 (.A1(W2522), .A2(I1015), .ZN(W8274));
  NANDX1 G25782 (.A1(W11), .A2(W5002), .ZN(W8200));
  NANDX1 G25783 (.A1(W6929), .A2(I1703), .ZN(W8203));
  NANDX1 G25784 (.A1(W1207), .A2(W10383), .ZN(W19049));
  NANDX1 G25785 (.A1(W15946), .A2(W12147), .ZN(W19048));
  NANDX1 G25786 (.A1(W2113), .A2(I967), .ZN(W4366));
  NANDX1 G25787 (.A1(W1286), .A2(W3217), .ZN(W4367));
  NANDX1 G25788 (.A1(W337), .A2(W3839), .ZN(W4372));
  NANDX1 G25789 (.A1(W18656), .A2(W8228), .ZN(W19043));
  NANDX1 G25790 (.A1(I1464), .A2(W2006), .ZN(W4374));
  NANDX1 G25791 (.A1(W2589), .A2(W5885), .ZN(W19041));
  NANDX1 G25792 (.A1(W1606), .A2(I198), .ZN(W4364));
  NANDX1 G25793 (.A1(W378), .A2(W2290), .ZN(W4376));
  NANDX1 G25794 (.A1(W2852), .A2(W1628), .ZN(W4380));
  NANDX1 G25795 (.A1(W1794), .A2(W1522), .ZN(W4385));
  NANDX1 G25796 (.A1(W17552), .A2(W6036), .ZN(O1693));
  NANDX1 G25797 (.A1(W2051), .A2(W923), .ZN(W4387));
  NANDX1 G25798 (.A1(W15428), .A2(W10166), .ZN(W19031));
  NANDX1 G25799 (.A1(W7556), .A2(W5837), .ZN(W19029));
  NANDX1 G25800 (.A1(W1053), .A2(W12), .ZN(O56));
  NANDX1 G25801 (.A1(W15422), .A2(W5753), .ZN(W19063));
  NANDX1 G25802 (.A1(I1597), .A2(W15978), .ZN(W19069));
  NANDX1 G25803 (.A1(W9292), .A2(W3697), .ZN(W13107));
  NANDX1 G25804 (.A1(I19), .A2(W628), .ZN(W4354));
  NANDX1 G25805 (.A1(W6144), .A2(W7686), .ZN(W8210));
  NANDX1 G25806 (.A1(W7355), .A2(W225), .ZN(W19067));
  NANDX1 G25807 (.A1(I1754), .A2(I1303), .ZN(W8208));
  NANDX1 G25808 (.A1(W7678), .A2(I725), .ZN(W8205));
  NANDX1 G25809 (.A1(W344), .A2(W4550), .ZN(W19064));
  NANDX1 G25810 (.A1(W18091), .A2(W3977), .ZN(W19027));
  NANDX1 G25811 (.A1(W11950), .A2(W7429), .ZN(O1698));
  NANDX1 G25812 (.A1(W17358), .A2(I727), .ZN(O1697));
  NANDX1 G25813 (.A1(W17217), .A2(W15358), .ZN(O1696));
  NANDX1 G25814 (.A1(W1898), .A2(W8686), .ZN(W13112));
  NANDX1 G25815 (.A1(W3146), .A2(I923), .ZN(W19057));
  NANDX1 G25816 (.A1(W941), .A2(W2146), .ZN(W4359));
  NANDX1 G25817 (.A1(I1393), .A2(W1530), .ZN(W19055));
  NANDX1 G25818 (.A1(W10791), .A2(W16939), .ZN(W19053));
  NANDX1 G25819 (.A1(I806), .A2(I1082), .ZN(W4408));
  NANDX1 G25820 (.A1(W6110), .A2(W8405), .ZN(W13124));
  NANDX1 G25821 (.A1(I1354), .A2(I1280), .ZN(W4400));
  NANDX1 G25822 (.A1(W6096), .A2(W1726), .ZN(W8192));
  NANDX1 G25823 (.A1(I928), .A2(W3578), .ZN(W4402));
  NANDX1 G25824 (.A1(W3675), .A2(W233), .ZN(W4404));
  NANDX1 G25825 (.A1(W4572), .A2(W17509), .ZN(W19003));
  NANDX1 G25826 (.A1(W12381), .A2(W4339), .ZN(W13125));
  NANDX1 G25827 (.A1(W8299), .A2(W17293), .ZN(W18996));
  NANDX1 G25828 (.A1(W2699), .A2(W7788), .ZN(W8193));
  NANDX1 G25829 (.A1(W4918), .A2(W6848), .ZN(W13128));
  NANDX1 G25830 (.A1(W18579), .A2(W13813), .ZN(W18993));
  NANDX1 G25831 (.A1(W4237), .A2(W16709), .ZN(W18989));
  NANDX1 G25832 (.A1(W7684), .A2(W3447), .ZN(W18988));
  NANDX1 G25833 (.A1(W3165), .A2(W3909), .ZN(W13129));
  NANDX1 G25834 (.A1(W3108), .A2(W6617), .ZN(W8189));
  NANDX1 G25835 (.A1(W12659), .A2(W10331), .ZN(W18986));
  NANDX1 G25836 (.A1(W6716), .A2(W3409), .ZN(O214));
  NANDX1 G25837 (.A1(W7804), .A2(W18502), .ZN(W19017));
  NANDX1 G25838 (.A1(W6401), .A2(W2629), .ZN(O698));
  NANDX1 G25839 (.A1(W2067), .A2(I1576), .ZN(W4393));
  NANDX1 G25840 (.A1(W15004), .A2(W6907), .ZN(W19026));
  NANDX1 G25841 (.A1(W1814), .A2(W4358), .ZN(W19024));
  NANDX1 G25842 (.A1(W5348), .A2(W3318), .ZN(O699));
  NANDX1 G25843 (.A1(W156), .A2(W11316), .ZN(W19022));
  NANDX1 G25844 (.A1(W5787), .A2(W2074), .ZN(W19021));
  NANDX1 G25845 (.A1(W910), .A2(I1982), .ZN(W19019));
  NANDX1 G25846 (.A1(W14157), .A2(W5910), .ZN(W19070));
  NANDX1 G25847 (.A1(W692), .A2(W6478), .ZN(W8197));
  NANDX1 G25848 (.A1(W7027), .A2(W8236), .ZN(O1692));
  NANDX1 G25849 (.A1(W2909), .A2(I32), .ZN(W4395));
  NANDX1 G25850 (.A1(W6358), .A2(W14018), .ZN(W19013));
  NANDX1 G25851 (.A1(W4988), .A2(W266), .ZN(W8195));
  NANDX1 G25852 (.A1(W14008), .A2(W3331), .ZN(W19012));
  NANDX1 G25853 (.A1(W4534), .A2(W6913), .ZN(W8194));
  NANDX1 G25854 (.A1(W1871), .A2(I1907), .ZN(W4397));
  NANDX1 G25855 (.A1(W2289), .A2(I1632), .ZN(W19119));
  NANDX1 G25856 (.A1(I1851), .A2(W10589), .ZN(W19131));
  NANDX1 G25857 (.A1(W5087), .A2(W18311), .ZN(W19129));
  NANDX1 G25858 (.A1(I5), .A2(W11327), .ZN(O692));
  NANDX1 G25859 (.A1(W3246), .A2(I1900), .ZN(W4308));
  NANDX1 G25860 (.A1(W16746), .A2(W15251), .ZN(W19124));
  NANDX1 G25861 (.A1(W2448), .A2(W3355), .ZN(W13081));
  NANDX1 G25862 (.A1(W3825), .A2(W70), .ZN(W8231));
  NANDX1 G25863 (.A1(W10447), .A2(W1461), .ZN(W13085));
  NANDX1 G25864 (.A1(W2220), .A2(W802), .ZN(W4313));
  NANDX1 G25865 (.A1(W4504), .A2(W17817), .ZN(O1712));
  NANDX1 G25866 (.A1(I1312), .A2(W3117), .ZN(W4316));
  NANDX1 G25867 (.A1(W14913), .A2(W1684), .ZN(O1709));
  NANDX1 G25868 (.A1(W7209), .A2(I1844), .ZN(W8229));
  NANDX1 G25869 (.A1(W5815), .A2(W11398), .ZN(W19117));
  NANDX1 G25870 (.A1(W7553), .A2(W7827), .ZN(W8227));
  NANDX1 G25871 (.A1(W11997), .A2(W8405), .ZN(W19113));
  NANDX1 G25872 (.A1(W1077), .A2(I1763), .ZN(W4319));
  NANDX1 G25873 (.A1(I1287), .A2(W4170), .ZN(W8226));
  NANDX1 G25874 (.A1(W168), .A2(I1284), .ZN(W19152));
  NANDX1 G25875 (.A1(I694), .A2(W586), .ZN(W4280));
  NANDX1 G25876 (.A1(I1353), .A2(I640), .ZN(W4281));
  NANDX1 G25877 (.A1(W1609), .A2(I654), .ZN(W4283));
  NANDX1 G25878 (.A1(I1441), .A2(W1614), .ZN(W4285));
  NANDX1 G25879 (.A1(W3513), .A2(W515), .ZN(W4287));
  NANDX1 G25880 (.A1(W3969), .A2(W7174), .ZN(W19157));
  NANDX1 G25881 (.A1(W15634), .A2(W8381), .ZN(W19156));
  NANDX1 G25882 (.A1(I175), .A2(W4167), .ZN(W4293));
  NANDX1 G25883 (.A1(W6423), .A2(W9400), .ZN(W19109));
  NANDX1 G25884 (.A1(W4085), .A2(W3252), .ZN(W19150));
  NANDX1 G25885 (.A1(W4843), .A2(W8893), .ZN(W19146));
  NANDX1 G25886 (.A1(W6028), .A2(W14696), .ZN(W19144));
  NANDX1 G25887 (.A1(W5177), .A2(W2397), .ZN(W8237));
  NANDX1 G25888 (.A1(W1308), .A2(W7109), .ZN(W13076));
  NANDX1 G25889 (.A1(W6134), .A2(W5749), .ZN(W13077));
  NANDX1 G25890 (.A1(W5183), .A2(W593), .ZN(W8236));
  NANDX1 G25891 (.A1(W12630), .A2(W8733), .ZN(W19134));
  NANDX1 G25892 (.A1(W2626), .A2(W1300), .ZN(W4342));
  NANDX1 G25893 (.A1(W670), .A2(W15018), .ZN(O1705));
  NANDX1 G25894 (.A1(W7306), .A2(W9982), .ZN(O1704));
  NANDX1 G25895 (.A1(W6879), .A2(W572), .ZN(W13100));
  NANDX1 G25896 (.A1(W579), .A2(W1825), .ZN(W4337));
  NANDX1 G25897 (.A1(I1370), .A2(W3574), .ZN(W4338));
  NANDX1 G25898 (.A1(W13893), .A2(I896), .ZN(W19080));
  NANDX1 G25899 (.A1(W5070), .A2(W7825), .ZN(W13102));
  NANDX1 G25900 (.A1(W2602), .A2(W5782), .ZN(W8216));
  NANDX1 G25901 (.A1(W4763), .A2(W3512), .ZN(W19089));
  NANDX1 G25902 (.A1(W12403), .A2(W1790), .ZN(W19076));
  NANDX1 G25903 (.A1(W1607), .A2(W431), .ZN(O1700));
  NANDX1 G25904 (.A1(W1989), .A2(W3575), .ZN(W4345));
  NANDX1 G25905 (.A1(W627), .A2(W1371), .ZN(W4346));
  NANDX1 G25906 (.A1(W10141), .A2(W4401), .ZN(W13104));
  NANDX1 G25907 (.A1(W10308), .A2(W14268), .ZN(W19072));
  NANDX1 G25908 (.A1(W6340), .A2(W7604), .ZN(W8214));
  NANDX1 G25909 (.A1(I568), .A2(I1577), .ZN(W4350));
  NANDX1 G25910 (.A1(W3546), .A2(W888), .ZN(W4326));
  NANDX1 G25911 (.A1(W10122), .A2(W5659), .ZN(W19108));
  NANDX1 G25912 (.A1(W3133), .A2(W1874), .ZN(W4321));
  NANDX1 G25913 (.A1(W1171), .A2(W3271), .ZN(W4323));
  NANDX1 G25914 (.A1(I538), .A2(W419), .ZN(W4324));
  NANDX1 G25915 (.A1(W8466), .A2(W2738), .ZN(W19098));
  NANDX1 G25916 (.A1(W7246), .A2(W12000), .ZN(O694));
  NANDX1 G25917 (.A1(W11795), .A2(W6969), .ZN(W13092));
  NANDX1 G25918 (.A1(W4527), .A2(W6100), .ZN(W8223));
  NANDX1 G25919 (.A1(W2955), .A2(W4309), .ZN(W4670));
  NANDX1 G25920 (.A1(W6398), .A2(W1512), .ZN(W8221));
  NANDX1 G25921 (.A1(W2316), .A2(W946), .ZN(W4328));
  NANDX1 G25922 (.A1(W4304), .A2(W1356), .ZN(W19096));
  NANDX1 G25923 (.A1(W6096), .A2(W7966), .ZN(W8219));
  NANDX1 G25924 (.A1(I235), .A2(W3867), .ZN(W4335));
  NANDX1 G25925 (.A1(I216), .A2(W12181), .ZN(W19094));
  NANDX1 G25926 (.A1(W7155), .A2(W5930), .ZN(W13095));
  NANDX1 G25927 (.A1(W16754), .A2(W14438), .ZN(W19090));
  NANDX1 G25928 (.A1(W6444), .A2(W12837), .ZN(W13545));
  NANDX1 G25929 (.A1(W7504), .A2(W8860), .ZN(W13540));
  NANDX1 G25930 (.A1(W9744), .A2(W7725), .ZN(W13541));
  NANDX1 G25931 (.A1(W3356), .A2(W294), .ZN(O68));
  NANDX1 G25932 (.A1(W3049), .A2(W841), .ZN(W4954));
  NANDX1 G25933 (.A1(W3095), .A2(W2427), .ZN(W4956));
  NANDX1 G25934 (.A1(I1086), .A2(W2156), .ZN(W13543));
  NANDX1 G25935 (.A1(W11518), .A2(W12662), .ZN(W13544));
  NANDX1 G25936 (.A1(W5400), .A2(I895), .ZN(W18147));
  NANDX1 G25937 (.A1(W4755), .A2(W3480), .ZN(W4957));
  NANDX1 G25938 (.A1(W9312), .A2(W8793), .ZN(W18162));
  NANDX1 G25939 (.A1(W5999), .A2(W16429), .ZN(W18145));
  NANDX1 G25940 (.A1(I1603), .A2(W3080), .ZN(W4958));
  NANDX1 G25941 (.A1(W13683), .A2(W10967), .ZN(W18138));
  NANDX1 G25942 (.A1(W3508), .A2(W1476), .ZN(W4959));
  NANDX1 G25943 (.A1(I1193), .A2(W4346), .ZN(W4960));
  NANDX1 G25944 (.A1(W16517), .A2(W1786), .ZN(W18137));
  NANDX1 G25945 (.A1(I434), .A2(W3756), .ZN(W4961));
  NANDX1 G25946 (.A1(W12488), .A2(W5671), .ZN(W13549));
  NANDX1 G25947 (.A1(I412), .A2(W1249), .ZN(W4939));
  NANDX1 G25948 (.A1(W194), .A2(I55), .ZN(W4925));
  NANDX1 G25949 (.A1(W1184), .A2(I1888), .ZN(W4927));
  NANDX1 G25950 (.A1(I1874), .A2(W5167), .ZN(W13529));
  NANDX1 G25951 (.A1(I1808), .A2(I1714), .ZN(W18182));
  NANDX1 G25952 (.A1(I634), .A2(W3586), .ZN(W4931));
  NANDX1 G25953 (.A1(W9139), .A2(W7028), .ZN(W13531));
  NANDX1 G25954 (.A1(W5784), .A2(W111), .ZN(W13532));
  NANDX1 G25955 (.A1(W1636), .A2(W4296), .ZN(W7935));
  NANDX1 G25956 (.A1(W2083), .A2(W4490), .ZN(W4965));
  NANDX1 G25957 (.A1(W12024), .A2(W1471), .ZN(O753));
  NANDX1 G25958 (.A1(W1900), .A2(W10861), .ZN(W18177));
  NANDX1 G25959 (.A1(I337), .A2(W3204), .ZN(O67));
  NANDX1 G25960 (.A1(W4468), .A2(W4651), .ZN(W4943));
  NANDX1 G25961 (.A1(W2875), .A2(W1119), .ZN(W4945));
  NANDX1 G25962 (.A1(W1142), .A2(W1491), .ZN(W4947));
  NANDX1 G25963 (.A1(W10226), .A2(I1982), .ZN(W18164));
  NANDX1 G25964 (.A1(W6118), .A2(W5396), .ZN(W7932));
  NANDX1 G25965 (.A1(W3886), .A2(W10754), .ZN(W13575));
  NANDX1 G25966 (.A1(W3355), .A2(W4453), .ZN(W4976));
  NANDX1 G25967 (.A1(I346), .A2(I1602), .ZN(O1503));
  NANDX1 G25968 (.A1(W4096), .A2(W1193), .ZN(W4978));
  NANDX1 G25969 (.A1(W4468), .A2(I376), .ZN(W4979));
  NANDX1 G25970 (.A1(I1722), .A2(W12368), .ZN(W18112));
  NANDX1 G25971 (.A1(W50), .A2(W3306), .ZN(W4981));
  NANDX1 G25972 (.A1(W1572), .A2(W8227), .ZN(W18110));
  NANDX1 G25973 (.A1(I1447), .A2(W15), .ZN(W4983));
  NANDX1 G25974 (.A1(W13287), .A2(W8740), .ZN(O1504));
  NANDX1 G25975 (.A1(W5648), .A2(W6554), .ZN(W7911));
  NANDX1 G25976 (.A1(W7320), .A2(I996), .ZN(W7910));
  NANDX1 G25977 (.A1(W2712), .A2(W1659), .ZN(W4985));
  NANDX1 G25978 (.A1(W5639), .A2(I718), .ZN(W7909));
  NANDX1 G25979 (.A1(W1288), .A2(W10362), .ZN(W18105));
  NANDX1 G25980 (.A1(W516), .A2(W13135), .ZN(W13579));
  NANDX1 G25981 (.A1(W1511), .A2(W2554), .ZN(W4993));
  NANDX1 G25982 (.A1(W1087), .A2(I1912), .ZN(W4994));
  NANDX1 G25983 (.A1(W2504), .A2(W6369), .ZN(W13561));
  NANDX1 G25984 (.A1(W13092), .A2(W9922), .ZN(W13555));
  NANDX1 G25985 (.A1(W8334), .A2(W8991), .ZN(W13557));
  NANDX1 G25986 (.A1(W13134), .A2(I32), .ZN(W18124));
  NANDX1 G25987 (.A1(I636), .A2(W6194), .ZN(O758));
  NANDX1 G25988 (.A1(W1814), .A2(W4225), .ZN(W4966));
  NANDX1 G25989 (.A1(W3573), .A2(W3024), .ZN(W4968));
  NANDX1 G25990 (.A1(I1072), .A2(W1432), .ZN(W4969));
  NANDX1 G25991 (.A1(W1759), .A2(W9873), .ZN(O1505));
  NANDX1 G25992 (.A1(W2487), .A2(W14252), .ZN(W18185));
  NANDX1 G25993 (.A1(W8575), .A2(W10396), .ZN(W18116));
  NANDX1 G25994 (.A1(W11273), .A2(W481), .ZN(W13563));
  NANDX1 G25995 (.A1(W312), .A2(I457), .ZN(W4970));
  NANDX1 G25996 (.A1(W1858), .A2(W4832), .ZN(W4972));
  NANDX1 G25997 (.A1(W7197), .A2(W6025), .ZN(W7915));
  NANDX1 G25998 (.A1(W7719), .A2(W4405), .ZN(W13571));
  NANDX1 G25999 (.A1(I922), .A2(I404), .ZN(W7913));
  NANDX1 G26000 (.A1(W4688), .A2(W1912), .ZN(W4975));
  NANDX1 G26001 (.A1(W5956), .A2(W1290), .ZN(W7964));
  NANDX1 G26002 (.A1(W7612), .A2(W4045), .ZN(W13494));
  NANDX1 G26003 (.A1(W8323), .A2(W2170), .ZN(W18257));
  NANDX1 G26004 (.A1(I715), .A2(I280), .ZN(W4891));
  NANDX1 G26005 (.A1(W11706), .A2(W8240), .ZN(W18254));
  NANDX1 G26006 (.A1(W6668), .A2(W17257), .ZN(O1526));
  NANDX1 G26007 (.A1(W11009), .A2(W17604), .ZN(W18249));
  NANDX1 G26008 (.A1(I241), .A2(W3773), .ZN(O66));
  NANDX1 G26009 (.A1(W10485), .A2(W5704), .ZN(W13499));
  NANDX1 G26010 (.A1(W5494), .A2(W14794), .ZN(W18248));
  NANDX1 G26011 (.A1(W13247), .A2(W13768), .ZN(W18260));
  NANDX1 G26012 (.A1(I1778), .A2(W5317), .ZN(W7963));
  NANDX1 G26013 (.A1(W535), .A2(W2049), .ZN(W4900));
  NANDX1 G26014 (.A1(W14771), .A2(W7935), .ZN(W18241));
  NANDX1 G26015 (.A1(W10823), .A2(W2255), .ZN(O1523));
  NANDX1 G26016 (.A1(W4885), .A2(W4867), .ZN(W18235));
  NANDX1 G26017 (.A1(W16951), .A2(W5794), .ZN(W18234));
  NANDX1 G26018 (.A1(W4993), .A2(W13711), .ZN(W18233));
  NANDX1 G26019 (.A1(W9941), .A2(W12271), .ZN(O1522));
  NANDX1 G26020 (.A1(W2788), .A2(W671), .ZN(W7969));
  NANDX1 G26021 (.A1(W6002), .A2(W269), .ZN(W7970));
  NANDX1 G26022 (.A1(W4155), .A2(W1205), .ZN(W18275));
  NANDX1 G26023 (.A1(W10611), .A2(W1796), .ZN(W18274));
  NANDX1 G26024 (.A1(W6007), .A2(W8474), .ZN(W13487));
  NANDX1 G26025 (.A1(I80), .A2(W14987), .ZN(W18270));
  NANDX1 G26026 (.A1(W3684), .A2(W2367), .ZN(W13488));
  NANDX1 G26027 (.A1(W8917), .A2(W5424), .ZN(W18268));
  NANDX1 G26028 (.A1(W4055), .A2(I1444), .ZN(W4884));
  NANDX1 G26029 (.A1(I1880), .A2(W1686), .ZN(W4901));
  NANDX1 G26030 (.A1(W545), .A2(W2122), .ZN(W4885));
  NANDX1 G26031 (.A1(I956), .A2(W1722), .ZN(W4886));
  NANDX1 G26032 (.A1(W3033), .A2(W8578), .ZN(W13489));
  NANDX1 G26033 (.A1(W761), .A2(I64), .ZN(W4888));
  NANDX1 G26034 (.A1(W3357), .A2(W5464), .ZN(W7968));
  NANDX1 G26035 (.A1(W1282), .A2(W8033), .ZN(O1531));
  NANDX1 G26036 (.A1(I394), .A2(W8411), .ZN(O1529));
  NANDX1 G26037 (.A1(W2230), .A2(W1327), .ZN(W7966));
  NANDX1 G26038 (.A1(W9765), .A2(W3220), .ZN(W18199));
  NANDX1 G26039 (.A1(W3802), .A2(W3728), .ZN(W4918));
  NANDX1 G26040 (.A1(W11540), .A2(W5544), .ZN(O1519));
  NANDX1 G26041 (.A1(W12674), .A2(W17727), .ZN(W18205));
  NANDX1 G26042 (.A1(W7612), .A2(W898), .ZN(W7946));
  NANDX1 G26043 (.A1(W381), .A2(I439), .ZN(W13517));
  NANDX1 G26044 (.A1(I1179), .A2(W2549), .ZN(W4920));
  NANDX1 G26045 (.A1(W3636), .A2(W16197), .ZN(W18203));
  NANDX1 G26046 (.A1(W583), .A2(W13242), .ZN(W13520));
  NANDX1 G26047 (.A1(W4800), .A2(W4019), .ZN(W7952));
  NANDX1 G26048 (.A1(W1381), .A2(W16170), .ZN(W18197));
  NANDX1 G26049 (.A1(W15667), .A2(W2830), .ZN(W18196));
  NANDX1 G26050 (.A1(W9358), .A2(I1348), .ZN(O1518));
  NANDX1 G26051 (.A1(W3173), .A2(W6079), .ZN(W13524));
  NANDX1 G26052 (.A1(W11099), .A2(W8825), .ZN(W13525));
  NANDX1 G26053 (.A1(W350), .A2(W6676), .ZN(W7937));
  NANDX1 G26054 (.A1(W8874), .A2(W1063), .ZN(W18187));
  NANDX1 G26055 (.A1(W6804), .A2(W856), .ZN(W13527));
  NANDX1 G26056 (.A1(W2142), .A2(I1880), .ZN(W4908));
  NANDX1 G26057 (.A1(W2138), .A2(W3069), .ZN(W4902));
  NANDX1 G26058 (.A1(W2254), .A2(W4803), .ZN(W4903));
  NANDX1 G26059 (.A1(W10323), .A2(W16683), .ZN(W18226));
  NANDX1 G26060 (.A1(I1988), .A2(W3875), .ZN(W7957));
  NANDX1 G26061 (.A1(W515), .A2(W4545), .ZN(W7956));
  NANDX1 G26062 (.A1(W8497), .A2(W6708), .ZN(W13504));
  NANDX1 G26063 (.A1(W2219), .A2(W3151), .ZN(W13505));
  NANDX1 G26064 (.A1(W7638), .A2(I1726), .ZN(W7955));
  NANDX1 G26065 (.A1(W7067), .A2(W6906), .ZN(W18101));
  NANDX1 G26066 (.A1(I1819), .A2(W2453), .ZN(W4909));
  NANDX1 G26067 (.A1(W12676), .A2(W9028), .ZN(W18216));
  NANDX1 G26068 (.A1(I1445), .A2(W4053), .ZN(W4912));
  NANDX1 G26069 (.A1(W4153), .A2(W2699), .ZN(O751));
  NANDX1 G26070 (.A1(W2980), .A2(W3090), .ZN(W4915));
  NANDX1 G26071 (.A1(W2705), .A2(W1335), .ZN(W7953));
  NANDX1 G26072 (.A1(W2878), .A2(W693), .ZN(W4916));
  NANDX1 G26073 (.A1(W1516), .A2(W6010), .ZN(W13516));
  NANDX1 G26074 (.A1(W938), .A2(I1255), .ZN(W5059));
  NANDX1 G26075 (.A1(W3540), .A2(W7701), .ZN(W17997));
  NANDX1 G26076 (.A1(W3427), .A2(W4771), .ZN(W5048));
  NANDX1 G26077 (.A1(I370), .A2(W10185), .ZN(W17995));
  NANDX1 G26078 (.A1(W2722), .A2(W927), .ZN(W13629));
  NANDX1 G26079 (.A1(I981), .A2(W2146), .ZN(W5054));
  NANDX1 G26080 (.A1(W2916), .A2(W5847), .ZN(W17988));
  NANDX1 G26081 (.A1(W15336), .A2(W3031), .ZN(W17987));
  NANDX1 G26082 (.A1(I1323), .A2(W6518), .ZN(W7870));
  NANDX1 G26083 (.A1(I501), .A2(W12019), .ZN(W13632));
  NANDX1 G26084 (.A1(W227), .A2(W17222), .ZN(W18000));
  NANDX1 G26085 (.A1(W114), .A2(W12052), .ZN(W17982));
  NANDX1 G26086 (.A1(W4814), .A2(W0), .ZN(W7864));
  NANDX1 G26087 (.A1(W813), .A2(W6296), .ZN(W17976));
  NANDX1 G26088 (.A1(W4477), .A2(W4609), .ZN(W13634));
  NANDX1 G26089 (.A1(W4290), .A2(W3659), .ZN(W5066));
  NANDX1 G26090 (.A1(W4498), .A2(W4150), .ZN(W5067));
  NANDX1 G26091 (.A1(W2104), .A2(W4469), .ZN(W5069));
  NANDX1 G26092 (.A1(W9474), .A2(W1998), .ZN(W17969));
  NANDX1 G26093 (.A1(W17946), .A2(W11127), .ZN(O1484));
  NANDX1 G26094 (.A1(W11788), .A2(W10388), .ZN(W18020));
  NANDX1 G26095 (.A1(I1301), .A2(W1882), .ZN(W13621));
  NANDX1 G26096 (.A1(W6406), .A2(W13533), .ZN(W18018));
  NANDX1 G26097 (.A1(W1868), .A2(I1277), .ZN(W5039));
  NANDX1 G26098 (.A1(W2823), .A2(I1547), .ZN(W5040));
  NANDX1 G26099 (.A1(W10567), .A2(W9336), .ZN(W18015));
  NANDX1 G26100 (.A1(W14138), .A2(W445), .ZN(W18014));
  NANDX1 G26101 (.A1(W13872), .A2(W14897), .ZN(W18013));
  NANDX1 G26102 (.A1(W8320), .A2(W2617), .ZN(W17967));
  NANDX1 G26103 (.A1(W2001), .A2(W1981), .ZN(W18010));
  NANDX1 G26104 (.A1(I1969), .A2(W3417), .ZN(W5042));
  NANDX1 G26105 (.A1(W639), .A2(I1302), .ZN(W13628));
  NANDX1 G26106 (.A1(W3614), .A2(W6515), .ZN(W18007));
  NANDX1 G26107 (.A1(W14110), .A2(W11953), .ZN(W18005));
  NANDX1 G26108 (.A1(W9981), .A2(W1695), .ZN(W18004));
  NANDX1 G26109 (.A1(W6948), .A2(W10327), .ZN(O1481));
  NANDX1 G26110 (.A1(W3029), .A2(W4517), .ZN(W7873));
  NANDX1 G26111 (.A1(W2113), .A2(W11316), .ZN(W13656));
  NANDX1 G26112 (.A1(W2284), .A2(W3444), .ZN(W5086));
  NANDX1 G26113 (.A1(W1213), .A2(W492), .ZN(O203));
  NANDX1 G26114 (.A1(W2430), .A2(W6568), .ZN(W17937));
  NANDX1 G26115 (.A1(W4609), .A2(W3223), .ZN(W5089));
  NANDX1 G26116 (.A1(W1813), .A2(W10880), .ZN(O768));
  NANDX1 G26117 (.A1(I503), .A2(W12799), .ZN(W17933));
  NANDX1 G26118 (.A1(W769), .A2(W3692), .ZN(W7846));
  NANDX1 G26119 (.A1(W6725), .A2(W12598), .ZN(W13655));
  NANDX1 G26120 (.A1(W3151), .A2(W8548), .ZN(W13647));
  NANDX1 G26121 (.A1(W6247), .A2(W2272), .ZN(W7845));
  NANDX1 G26122 (.A1(W1823), .A2(W4224), .ZN(W5092));
  NANDX1 G26123 (.A1(W9259), .A2(W9535), .ZN(O770));
  NANDX1 G26124 (.A1(I1220), .A2(W8971), .ZN(O1469));
  NANDX1 G26125 (.A1(W3831), .A2(W5754), .ZN(O1468));
  NANDX1 G26126 (.A1(W447), .A2(I1930), .ZN(W5100));
  NANDX1 G26127 (.A1(W15735), .A2(W15224), .ZN(W17922));
  NANDX1 G26128 (.A1(W1876), .A2(W4114), .ZN(W17921));
  NANDX1 G26129 (.A1(W10336), .A2(W15627), .ZN(W17950));
  NANDX1 G26130 (.A1(W2828), .A2(W584), .ZN(W13635));
  NANDX1 G26131 (.A1(W10187), .A2(W3555), .ZN(O1477));
  NANDX1 G26132 (.A1(I191), .A2(I950), .ZN(W5073));
  NANDX1 G26133 (.A1(W11460), .A2(W9306), .ZN(W17960));
  NANDX1 G26134 (.A1(I1582), .A2(W16421), .ZN(W17959));
  NANDX1 G26135 (.A1(W1418), .A2(W8283), .ZN(O1476));
  NANDX1 G26136 (.A1(W6610), .A2(W7), .ZN(W7858));
  NANDX1 G26137 (.A1(W16035), .A2(I1638), .ZN(W17953));
  NANDX1 G26138 (.A1(W3881), .A2(I1850), .ZN(W7876));
  NANDX1 G26139 (.A1(W4760), .A2(I393), .ZN(W5076));
  NANDX1 G26140 (.A1(W6969), .A2(W7881), .ZN(O1474));
  NANDX1 G26141 (.A1(W12082), .A2(W13059), .ZN(W13638));
  NANDX1 G26142 (.A1(W1634), .A2(I1862), .ZN(W7851));
  NANDX1 G26143 (.A1(W1992), .A2(W7733), .ZN(W13643));
  NANDX1 G26144 (.A1(W1303), .A2(W4003), .ZN(W7850));
  NANDX1 G26145 (.A1(W13130), .A2(W8619), .ZN(W13644));
  NANDX1 G26146 (.A1(W4166), .A2(W298), .ZN(W5084));
  NANDX1 G26147 (.A1(W12762), .A2(W3815), .ZN(W13598));
  NANDX1 G26148 (.A1(W1033), .A2(W13778), .ZN(W18074));
  NANDX1 G26149 (.A1(W4057), .A2(W9814), .ZN(O764));
  NANDX1 G26150 (.A1(W860), .A2(W7111), .ZN(O1497));
  NANDX1 G26151 (.A1(W707), .A2(I1962), .ZN(W5009));
  NANDX1 G26152 (.A1(W3834), .A2(I967), .ZN(W5011));
  NANDX1 G26153 (.A1(W9433), .A2(W1579), .ZN(O1496));
  NANDX1 G26154 (.A1(W6762), .A2(W2211), .ZN(W18070));
  NANDX1 G26155 (.A1(I82), .A2(W7819), .ZN(W18069));
  NANDX1 G26156 (.A1(W226), .A2(W619), .ZN(W13597));
  NANDX1 G26157 (.A1(W3765), .A2(W4791), .ZN(O70));
  NANDX1 G26158 (.A1(W479), .A2(W1010), .ZN(O71));
  NANDX1 G26159 (.A1(W3171), .A2(W6370), .ZN(W7898));
  NANDX1 G26160 (.A1(W12616), .A2(W7993), .ZN(W13600));
  NANDX1 G26161 (.A1(W11129), .A2(W8111), .ZN(W18062));
  NANDX1 G26162 (.A1(W1804), .A2(W1964), .ZN(W5015));
  NANDX1 G26163 (.A1(W3669), .A2(W4720), .ZN(W13601));
  NANDX1 G26164 (.A1(W2848), .A2(W4790), .ZN(W5018));
  NANDX1 G26165 (.A1(W911), .A2(W13647), .ZN(W18057));
  NANDX1 G26166 (.A1(W8364), .A2(W8584), .ZN(O1500));
  NANDX1 G26167 (.A1(W17962), .A2(W11993), .ZN(W18099));
  NANDX1 G26168 (.A1(W3242), .A2(W6794), .ZN(W13583));
  NANDX1 G26169 (.A1(W4383), .A2(W8371), .ZN(W13584));
  NANDX1 G26170 (.A1(W4095), .A2(W3118), .ZN(W13585));
  NANDX1 G26171 (.A1(W10235), .A2(W10480), .ZN(W13586));
  NANDX1 G26172 (.A1(W2403), .A2(I1557), .ZN(W5002));
  NANDX1 G26173 (.A1(W3775), .A2(W10114), .ZN(W18091));
  NANDX1 G26174 (.A1(W4897), .A2(W15486), .ZN(W18090));
  NANDX1 G26175 (.A1(I1378), .A2(W697), .ZN(W13602));
  NANDX1 G26176 (.A1(W2511), .A2(W10549), .ZN(W18087));
  NANDX1 G26177 (.A1(W10386), .A2(W12539), .ZN(W13588));
  NANDX1 G26178 (.A1(W7303), .A2(W12314), .ZN(W18085));
  NANDX1 G26179 (.A1(W4438), .A2(W16098), .ZN(W18084));
  NANDX1 G26180 (.A1(W4088), .A2(W2478), .ZN(W7904));
  NANDX1 G26181 (.A1(W7737), .A2(W8453), .ZN(O1498));
  NANDX1 G26182 (.A1(I290), .A2(W7979), .ZN(W18079));
  NANDX1 G26183 (.A1(W11800), .A2(I1364), .ZN(W13595));
  NANDX1 G26184 (.A1(W4274), .A2(W13255), .ZN(W13614));
  NANDX1 G26185 (.A1(I489), .A2(W14610), .ZN(W18042));
  NANDX1 G26186 (.A1(W15209), .A2(W1901), .ZN(W18039));
  NANDX1 G26187 (.A1(W2500), .A2(I1072), .ZN(W5028));
  NANDX1 G26188 (.A1(W2577), .A2(I1245), .ZN(W7884));
  NANDX1 G26189 (.A1(W6299), .A2(W3088), .ZN(W13612));
  NANDX1 G26190 (.A1(W13498), .A2(W11513), .ZN(O1488));
  NANDX1 G26191 (.A1(I1547), .A2(W4679), .ZN(W18031));
  NANDX1 G26192 (.A1(W1435), .A2(W11320), .ZN(W13613));
  NANDX1 G26193 (.A1(W17037), .A2(W12398), .ZN(W18043));
  NANDX1 G26194 (.A1(W3349), .A2(W1849), .ZN(W7881));
  NANDX1 G26195 (.A1(W12137), .A2(W4541), .ZN(W13615));
  NANDX1 G26196 (.A1(W6662), .A2(W2920), .ZN(W7880));
  NANDX1 G26197 (.A1(W8346), .A2(W9302), .ZN(O1487));
  NANDX1 G26198 (.A1(I895), .A2(W348), .ZN(W7879));
  NANDX1 G26199 (.A1(I18), .A2(W10583), .ZN(O766));
  NANDX1 G26200 (.A1(W3851), .A2(W260), .ZN(W5034));
  NANDX1 G26201 (.A1(W4795), .A2(I873), .ZN(W7878));
  NANDX1 G26202 (.A1(W1954), .A2(W570), .ZN(W5022));
  NANDX1 G26203 (.A1(W16192), .A2(W8436), .ZN(W18055));
  NANDX1 G26204 (.A1(I519), .A2(W2544), .ZN(W5019));
  NANDX1 G26205 (.A1(W1157), .A2(I895), .ZN(W7896));
  NANDX1 G26206 (.A1(W7767), .A2(W5380), .ZN(W7894));
  NANDX1 G26207 (.A1(W5223), .A2(W16403), .ZN(W18051));
  NANDX1 G26208 (.A1(W2720), .A2(W1329), .ZN(W7892));
  NANDX1 G26209 (.A1(W5008), .A2(W4033), .ZN(W18049));
  NANDX1 G26210 (.A1(W2593), .A2(W4866), .ZN(W5021));
  NANDX1 G26211 (.A1(W85), .A2(W4190), .ZN(W7972));
  NANDX1 G26212 (.A1(W3684), .A2(W4933), .ZN(W5024));
  NANDX1 G26213 (.A1(W10842), .A2(W4804), .ZN(W18048));
  NANDX1 G26214 (.A1(W4965), .A2(I1634), .ZN(W7888));
  NANDX1 G26215 (.A1(W4687), .A2(W2228), .ZN(W5026));
  NANDX1 G26216 (.A1(W12439), .A2(W7995), .ZN(W18047));
  NANDX1 G26217 (.A1(W12506), .A2(W12151), .ZN(W18046));
  NANDX1 G26218 (.A1(W13545), .A2(W4482), .ZN(O1489));
  NANDX1 G26219 (.A1(W2264), .A2(I1060), .ZN(W5027));
  NANDX1 G26220 (.A1(W11752), .A2(W17050), .ZN(W18494));
  NANDX1 G26221 (.A1(W16282), .A2(W5636), .ZN(W18504));
  NANDX1 G26222 (.A1(W592), .A2(W8566), .ZN(W13359));
  NANDX1 G26223 (.A1(W8706), .A2(W8943), .ZN(W13361));
  NANDX1 G26224 (.A1(W3997), .A2(I1262), .ZN(W4740));
  NANDX1 G26225 (.A1(W4262), .A2(W4819), .ZN(W18502));
  NANDX1 G26226 (.A1(W1143), .A2(W4009), .ZN(W4741));
  NANDX1 G26227 (.A1(W2555), .A2(W7865), .ZN(W18499));
  NANDX1 G26228 (.A1(W13029), .A2(W8790), .ZN(W18498));
  NANDX1 G26229 (.A1(W7615), .A2(W10400), .ZN(O1574));
  NANDX1 G26230 (.A1(W5154), .A2(W6336), .ZN(O735));
  NANDX1 G26231 (.A1(I1497), .A2(W11149), .ZN(W13365));
  NANDX1 G26232 (.A1(W12783), .A2(I1132), .ZN(W13368));
  NANDX1 G26233 (.A1(W16338), .A2(W15385), .ZN(O1573));
  NANDX1 G26234 (.A1(W12732), .A2(W998), .ZN(W18489));
  NANDX1 G26235 (.A1(W10857), .A2(W11731), .ZN(W13369));
  NANDX1 G26236 (.A1(W148), .A2(W3166), .ZN(W8037));
  NANDX1 G26237 (.A1(I186), .A2(W16781), .ZN(W18486));
  NANDX1 G26238 (.A1(W10799), .A2(W12384), .ZN(W13374));
  NANDX1 G26239 (.A1(W3255), .A2(W3694), .ZN(W8046));
  NANDX1 G26240 (.A1(W728), .A2(W1069), .ZN(W4725));
  NANDX1 G26241 (.A1(W1713), .A2(W12362), .ZN(W18530));
  NANDX1 G26242 (.A1(W16409), .A2(I1709), .ZN(O1582));
  NANDX1 G26243 (.A1(W871), .A2(W17530), .ZN(O1581));
  NANDX1 G26244 (.A1(I1863), .A2(W3250), .ZN(W18527));
  NANDX1 G26245 (.A1(W6969), .A2(I378), .ZN(W8053));
  NANDX1 G26246 (.A1(W662), .A2(W3952), .ZN(W8052));
  NANDX1 G26247 (.A1(W1823), .A2(W7711), .ZN(W8049));
  NANDX1 G26248 (.A1(W7993), .A2(W638), .ZN(W18484));
  NANDX1 G26249 (.A1(W15911), .A2(W14115), .ZN(W18515));
  NANDX1 G26250 (.A1(W2442), .A2(W923), .ZN(W4731));
  NANDX1 G26251 (.A1(W2587), .A2(W2894), .ZN(W18512));
  NANDX1 G26252 (.A1(W4533), .A2(I1570), .ZN(W18511));
  NANDX1 G26253 (.A1(W12311), .A2(W16923), .ZN(W18510));
  NANDX1 G26254 (.A1(W8253), .A2(W15548), .ZN(W18509));
  NANDX1 G26255 (.A1(W1558), .A2(W3983), .ZN(W13357));
  NANDX1 G26256 (.A1(W17264), .A2(I708), .ZN(W18508));
  NANDX1 G26257 (.A1(W12840), .A2(W12341), .ZN(W13394));
  NANDX1 G26258 (.A1(W6320), .A2(I1932), .ZN(W8028));
  NANDX1 G26259 (.A1(W8910), .A2(W13246), .ZN(W13391));
  NANDX1 G26260 (.A1(W3661), .A2(W6432), .ZN(W8027));
  NANDX1 G26261 (.A1(W1076), .A2(W11211), .ZN(W18463));
  NANDX1 G26262 (.A1(W7743), .A2(W8536), .ZN(W13393));
  NANDX1 G26263 (.A1(W5158), .A2(W2642), .ZN(W18461));
  NANDX1 G26264 (.A1(W3707), .A2(W232), .ZN(W4777));
  NANDX1 G26265 (.A1(W6792), .A2(W8925), .ZN(O1571));
  NANDX1 G26266 (.A1(W1158), .A2(W2921), .ZN(W4768));
  NANDX1 G26267 (.A1(W484), .A2(W1686), .ZN(W18457));
  NANDX1 G26268 (.A1(W4385), .A2(I668), .ZN(W4778));
  NANDX1 G26269 (.A1(I912), .A2(W4748), .ZN(W4779));
  NANDX1 G26270 (.A1(W335), .A2(W1839), .ZN(O737));
  NANDX1 G26271 (.A1(W3455), .A2(W2073), .ZN(W4781));
  NANDX1 G26272 (.A1(W4229), .A2(W5324), .ZN(W13398));
  NANDX1 G26273 (.A1(W4997), .A2(W6383), .ZN(W18453));
  NANDX1 G26274 (.A1(W14646), .A2(W12058), .ZN(O1570));
  NANDX1 G26275 (.A1(I223), .A2(W4083), .ZN(W8031));
  NANDX1 G26276 (.A1(W4418), .A2(W10180), .ZN(W18483));
  NANDX1 G26277 (.A1(W815), .A2(W1382), .ZN(W4750));
  NANDX1 G26278 (.A1(W11905), .A2(W2986), .ZN(W18482));
  NANDX1 G26279 (.A1(W1569), .A2(W9689), .ZN(W13377));
  NANDX1 G26280 (.A1(W9056), .A2(W635), .ZN(W13381));
  NANDX1 G26281 (.A1(W455), .A2(W64), .ZN(W4754));
  NANDX1 G26282 (.A1(I11), .A2(W1103), .ZN(W4756));
  NANDX1 G26283 (.A1(I1300), .A2(W2138), .ZN(W4757));
  NANDX1 G26284 (.A1(W9727), .A2(W18330), .ZN(W18535));
  NANDX1 G26285 (.A1(W6750), .A2(W5570), .ZN(W18475));
  NANDX1 G26286 (.A1(W8760), .A2(W11651), .ZN(W18474));
  NANDX1 G26287 (.A1(W12860), .A2(W12797), .ZN(W13386));
  NANDX1 G26288 (.A1(W1903), .A2(W2431), .ZN(W4763));
  NANDX1 G26289 (.A1(W12616), .A2(W4577), .ZN(W18469));
  NANDX1 G26290 (.A1(W8017), .A2(W7461), .ZN(W13388));
  NANDX1 G26291 (.A1(I1177), .A2(W928), .ZN(W4766));
  NANDX1 G26292 (.A1(W1494), .A2(W3386), .ZN(W4767));
  NANDX1 G26293 (.A1(I1079), .A2(W18013), .ZN(W18596));
  NANDX1 G26294 (.A1(W9691), .A2(W8394), .ZN(W13323));
  NANDX1 G26295 (.A1(W13171), .A2(W5376), .ZN(W18605));
  NANDX1 G26296 (.A1(W10103), .A2(W5829), .ZN(W18604));
  NANDX1 G26297 (.A1(W1139), .A2(W5779), .ZN(W8069));
  NANDX1 G26298 (.A1(W2665), .A2(W1625), .ZN(W4691));
  NANDX1 G26299 (.A1(W6069), .A2(W16545), .ZN(W18602));
  NANDX1 G26300 (.A1(W18435), .A2(W16001), .ZN(W18601));
  NANDX1 G26301 (.A1(W5703), .A2(I16), .ZN(W8066));
  NANDX1 G26302 (.A1(W14759), .A2(W2528), .ZN(W18597));
  NANDX1 G26303 (.A1(I1403), .A2(W4636), .ZN(W4687));
  NANDX1 G26304 (.A1(W10297), .A2(W9822), .ZN(W13327));
  NANDX1 G26305 (.A1(W12305), .A2(W10158), .ZN(W18594));
  NANDX1 G26306 (.A1(W1118), .A2(W1168), .ZN(W4695));
  NANDX1 G26307 (.A1(W1656), .A2(I1751), .ZN(W4696));
  NANDX1 G26308 (.A1(W11003), .A2(W10133), .ZN(W13329));
  NANDX1 G26309 (.A1(I1042), .A2(W2867), .ZN(W18590));
  NANDX1 G26310 (.A1(W9722), .A2(W1191), .ZN(W18589));
  NANDX1 G26311 (.A1(W12700), .A2(W8255), .ZN(O1595));
  NANDX1 G26312 (.A1(I1553), .A2(W6655), .ZN(W18620));
  NANDX1 G26313 (.A1(W1845), .A2(W2614), .ZN(W4673));
  NANDX1 G26314 (.A1(W5683), .A2(W10291), .ZN(W13311));
  NANDX1 G26315 (.A1(I713), .A2(W15502), .ZN(W18629));
  NANDX1 G26316 (.A1(W205), .A2(W4898), .ZN(W8073));
  NANDX1 G26317 (.A1(I877), .A2(W2396), .ZN(W4678));
  NANDX1 G26318 (.A1(W8304), .A2(W9412), .ZN(W13312));
  NANDX1 G26319 (.A1(I1854), .A2(W1256), .ZN(W4682));
  NANDX1 G26320 (.A1(W11925), .A2(W7893), .ZN(O726));
  NANDX1 G26321 (.A1(W2729), .A2(W2939), .ZN(O730));
  NANDX1 G26322 (.A1(I1403), .A2(W2079), .ZN(W8071));
  NANDX1 G26323 (.A1(W3473), .A2(I672), .ZN(W4683));
  NANDX1 G26324 (.A1(W8178), .A2(W2030), .ZN(W13320));
  NANDX1 G26325 (.A1(W2852), .A2(I1804), .ZN(W8070));
  NANDX1 G26326 (.A1(W18257), .A2(W7619), .ZN(O1603));
  NANDX1 G26327 (.A1(W2298), .A2(W8099), .ZN(W13321));
  NANDX1 G26328 (.A1(W147), .A2(I1577), .ZN(W4686));
  NANDX1 G26329 (.A1(W7220), .A2(W6753), .ZN(O1601));
  NANDX1 G26330 (.A1(W257), .A2(I656), .ZN(W18548));
  NANDX1 G26331 (.A1(W5126), .A2(W7304), .ZN(W13344));
  NANDX1 G26332 (.A1(I298), .A2(W14679), .ZN(W18556));
  NANDX1 G26333 (.A1(I831), .A2(W5319), .ZN(W18555));
  NANDX1 G26334 (.A1(W2231), .A2(W11889), .ZN(W18554));
  NANDX1 G26335 (.A1(W4551), .A2(W4681), .ZN(W4717));
  NANDX1 G26336 (.A1(W1820), .A2(I456), .ZN(W13348));
  NANDX1 G26337 (.A1(W4119), .A2(W18461), .ZN(W18550));
  NANDX1 G26338 (.A1(W582), .A2(W4420), .ZN(W4718));
  NANDX1 G26339 (.A1(W11426), .A2(W3964), .ZN(W18557));
  NANDX1 G26340 (.A1(W3114), .A2(W4404), .ZN(W18546));
  NANDX1 G26341 (.A1(W4656), .A2(W2199), .ZN(W4719));
  NANDX1 G26342 (.A1(W2967), .A2(W2168), .ZN(W4722));
  NANDX1 G26343 (.A1(W483), .A2(W3824), .ZN(W4723));
  NANDX1 G26344 (.A1(W130), .A2(I567), .ZN(W18541));
  NANDX1 G26345 (.A1(W8762), .A2(W16142), .ZN(W18539));
  NANDX1 G26346 (.A1(W3702), .A2(W7405), .ZN(W18536));
  NANDX1 G26347 (.A1(W3855), .A2(W4200), .ZN(W4724));
  NANDX1 G26348 (.A1(W3806), .A2(W719), .ZN(W8059));
  NANDX1 G26349 (.A1(W4554), .A2(W397), .ZN(W4705));
  NANDX1 G26350 (.A1(W5389), .A2(W191), .ZN(W8064));
  NANDX1 G26351 (.A1(W197), .A2(W3320), .ZN(W4706));
  NANDX1 G26352 (.A1(W18452), .A2(W18168), .ZN(O1591));
  NANDX1 G26353 (.A1(W7894), .A2(W9163), .ZN(W13332));
  NANDX1 G26354 (.A1(W110), .A2(W4649), .ZN(W8063));
  NANDX1 G26355 (.A1(W2230), .A2(W3773), .ZN(W13336));
  NANDX1 G26356 (.A1(W7422), .A2(W14895), .ZN(W18572));
  NANDX1 G26357 (.A1(I735), .A2(W11963), .ZN(W18450));
  NANDX1 G26358 (.A1(I1004), .A2(W89), .ZN(W4712));
  NANDX1 G26359 (.A1(I90), .A2(W7010), .ZN(O210));
  NANDX1 G26360 (.A1(W4792), .A2(W4907), .ZN(W8057));
  NANDX1 G26361 (.A1(W15072), .A2(W2567), .ZN(W18565));
  NANDX1 G26362 (.A1(W3336), .A2(W7248), .ZN(W8056));
  NANDX1 G26363 (.A1(W253), .A2(W3), .ZN(O1586));
  NANDX1 G26364 (.A1(W99), .A2(I137), .ZN(W13341));
  NANDX1 G26365 (.A1(W3786), .A2(W7113), .ZN(W8055));
  NANDX1 G26366 (.A1(W7679), .A2(W14267), .ZN(O1548));
  NANDX1 G26367 (.A1(I1326), .A2(W4314), .ZN(W4840));
  NANDX1 G26368 (.A1(W2021), .A2(I1692), .ZN(O1551));
  NANDX1 G26369 (.A1(I50), .A2(W3253), .ZN(W4842));
  NANDX1 G26370 (.A1(I547), .A2(W1809), .ZN(W4843));
  NANDX1 G26371 (.A1(W3395), .A2(W6267), .ZN(W7987));
  NANDX1 G26372 (.A1(W2190), .A2(W2383), .ZN(O1550));
  NANDX1 G26373 (.A1(W11313), .A2(W5707), .ZN(W18337));
  NANDX1 G26374 (.A1(I194), .A2(W1568), .ZN(W7984));
  NANDX1 G26375 (.A1(I640), .A2(I1763), .ZN(W4845));
  NANDX1 G26376 (.A1(I879), .A2(W6861), .ZN(W18343));
  NANDX1 G26377 (.A1(W9241), .A2(I1215), .ZN(W13465));
  NANDX1 G26378 (.A1(W4898), .A2(W4938), .ZN(W7983));
  NANDX1 G26379 (.A1(W9510), .A2(W4404), .ZN(W18327));
  NANDX1 G26380 (.A1(W7013), .A2(W340), .ZN(W7981));
  NANDX1 G26381 (.A1(W4348), .A2(W2143), .ZN(W18323));
  NANDX1 G26382 (.A1(W2482), .A2(W9586), .ZN(O1545));
  NANDX1 G26383 (.A1(W2570), .A2(I1542), .ZN(W13467));
  NANDX1 G26384 (.A1(I618), .A2(W223), .ZN(W4851));
  NANDX1 G26385 (.A1(W8353), .A2(W7747), .ZN(W18352));
  NANDX1 G26386 (.A1(W2177), .A2(W7406), .ZN(W13452));
  NANDX1 G26387 (.A1(W1255), .A2(W7340), .ZN(W13453));
  NANDX1 G26388 (.A1(W6602), .A2(W4955), .ZN(W18361));
  NANDX1 G26389 (.A1(W585), .A2(W1022), .ZN(W4833));
  NANDX1 G26390 (.A1(W1385), .A2(I181), .ZN(W7991));
  NANDX1 G26391 (.A1(W8949), .A2(W15443), .ZN(W18355));
  NANDX1 G26392 (.A1(W6746), .A2(W3106), .ZN(W13457));
  NANDX1 G26393 (.A1(W6742), .A2(I1937), .ZN(W18354));
  NANDX1 G26394 (.A1(W4808), .A2(W3369), .ZN(W7980));
  NANDX1 G26395 (.A1(W15480), .A2(W2214), .ZN(O1555));
  NANDX1 G26396 (.A1(W18145), .A2(W14327), .ZN(O1554));
  NANDX1 G26397 (.A1(W7413), .A2(W5213), .ZN(W7990));
  NANDX1 G26398 (.A1(W1578), .A2(W3226), .ZN(W4837));
  NANDX1 G26399 (.A1(W1672), .A2(W4342), .ZN(O744));
  NANDX1 G26400 (.A1(W3486), .A2(W3822), .ZN(O1552));
  NANDX1 G26401 (.A1(W4109), .A2(W6261), .ZN(W7989));
  NANDX1 G26402 (.A1(W14981), .A2(W4066), .ZN(W18344));
  NANDX1 G26403 (.A1(W13487), .A2(W6793), .ZN(W18286));
  NANDX1 G26404 (.A1(W4665), .A2(W563), .ZN(W4866));
  NANDX1 G26405 (.A1(W12303), .A2(W3357), .ZN(W18297));
  NANDX1 G26406 (.A1(W2145), .A2(W8801), .ZN(W18294));
  NANDX1 G26407 (.A1(W14726), .A2(W9375), .ZN(W18293));
  NANDX1 G26408 (.A1(W2758), .A2(W3021), .ZN(W4869));
  NANDX1 G26409 (.A1(W3155), .A2(W2819), .ZN(O65));
  NANDX1 G26410 (.A1(I263), .A2(W12726), .ZN(W18288));
  NANDX1 G26411 (.A1(W2745), .A2(W4541), .ZN(W4875));
  NANDX1 G26412 (.A1(I1482), .A2(W3650), .ZN(W18301));
  NANDX1 G26413 (.A1(W10319), .A2(W10933), .ZN(O1537));
  NANDX1 G26414 (.A1(W17566), .A2(W576), .ZN(O1536));
  NANDX1 G26415 (.A1(W17785), .A2(W5180), .ZN(W18282));
  NANDX1 G26416 (.A1(W4797), .A2(W12362), .ZN(W18280));
  NANDX1 G26417 (.A1(W7957), .A2(W16264), .ZN(W18279));
  NANDX1 G26418 (.A1(W4497), .A2(W1252), .ZN(W7973));
  NANDX1 G26419 (.A1(I1358), .A2(W13137), .ZN(W18277));
  NANDX1 G26420 (.A1(W12455), .A2(W9338), .ZN(W13484));
  NANDX1 G26421 (.A1(W6365), .A2(W12374), .ZN(W13474));
  NANDX1 G26422 (.A1(W3699), .A2(W1695), .ZN(W18318));
  NANDX1 G26423 (.A1(I126), .A2(W1400), .ZN(W18317));
  NANDX1 G26424 (.A1(W6075), .A2(W9087), .ZN(W13470));
  NANDX1 G26425 (.A1(W5262), .A2(W2864), .ZN(O1543));
  NANDX1 G26426 (.A1(I514), .A2(W3252), .ZN(O1542));
  NANDX1 G26427 (.A1(W2013), .A2(W4430), .ZN(W4855));
  NANDX1 G26428 (.A1(W5214), .A2(W9411), .ZN(W13473));
  NANDX1 G26429 (.A1(W16369), .A2(W5977), .ZN(W18310));
  NANDX1 G26430 (.A1(W14061), .A2(W1449), .ZN(W18365));
  NANDX1 G26431 (.A1(W11129), .A2(W9361), .ZN(W18308));
  NANDX1 G26432 (.A1(W7417), .A2(W10535), .ZN(W18307));
  NANDX1 G26433 (.A1(W249), .A2(W8977), .ZN(W13475));
  NANDX1 G26434 (.A1(W5536), .A2(W8656), .ZN(O747));
  NANDX1 G26435 (.A1(W2886), .A2(I590), .ZN(W7978));
  NANDX1 G26436 (.A1(W12539), .A2(W1989), .ZN(W13478));
  NANDX1 G26437 (.A1(I1851), .A2(I1564), .ZN(W4864));
  NANDX1 G26438 (.A1(W4514), .A2(W1967), .ZN(W4865));
  NANDX1 G26439 (.A1(I1266), .A2(I4), .ZN(W13418));
  NANDX1 G26440 (.A1(W5341), .A2(W1903), .ZN(O1565));
  NANDX1 G26441 (.A1(W1249), .A2(I388), .ZN(W4798));
  NANDX1 G26442 (.A1(W263), .A2(W1937), .ZN(W18425));
  NANDX1 G26443 (.A1(W675), .A2(I21), .ZN(W4799));
  NANDX1 G26444 (.A1(I771), .A2(W5294), .ZN(W13412));
  NANDX1 G26445 (.A1(W5837), .A2(W8986), .ZN(W13413));
  NANDX1 G26446 (.A1(I413), .A2(W1817), .ZN(W4802));
  NANDX1 G26447 (.A1(W381), .A2(W3395), .ZN(O739));
  NANDX1 G26448 (.A1(W7427), .A2(W8974), .ZN(W13417));
  NANDX1 G26449 (.A1(W4921), .A2(W14019), .ZN(W18428));
  NANDX1 G26450 (.A1(W465), .A2(W314), .ZN(W4804));
  NANDX1 G26451 (.A1(W6129), .A2(W7140), .ZN(W8010));
  NANDX1 G26452 (.A1(I1983), .A2(W2295), .ZN(W13424));
  NANDX1 G26453 (.A1(W860), .A2(W7272), .ZN(W13425));
  NANDX1 G26454 (.A1(W10784), .A2(W17886), .ZN(W18414));
  NANDX1 G26455 (.A1(I649), .A2(W2350), .ZN(W4811));
  NANDX1 G26456 (.A1(W7397), .A2(W8654), .ZN(W13427));
  NANDX1 G26457 (.A1(W1574), .A2(W3803), .ZN(O64));
  NANDX1 G26458 (.A1(W17135), .A2(W9288), .ZN(W18438));
  NANDX1 G26459 (.A1(W8495), .A2(I572), .ZN(W18447));
  NANDX1 G26460 (.A1(W4136), .A2(W5907), .ZN(W13408));
  NANDX1 G26461 (.A1(W3890), .A2(I792), .ZN(W4791));
  NANDX1 G26462 (.A1(W590), .A2(W477), .ZN(W4793));
  NANDX1 G26463 (.A1(W3547), .A2(W3784), .ZN(W4795));
  NANDX1 G26464 (.A1(W11878), .A2(W16620), .ZN(W18442));
  NANDX1 G26465 (.A1(W8347), .A2(W10819), .ZN(W18440));
  NANDX1 G26466 (.A1(W1432), .A2(W2647), .ZN(W4797));
  NANDX1 G26467 (.A1(W14831), .A2(W13320), .ZN(W18410));
  NANDX1 G26468 (.A1(I1079), .A2(W5772), .ZN(W13409));
  NANDX1 G26469 (.A1(W13176), .A2(W3121), .ZN(W18437));
  NANDX1 G26470 (.A1(W12239), .A2(W11158), .ZN(W18436));
  NANDX1 G26471 (.A1(W17773), .A2(W17962), .ZN(W18435));
  NANDX1 G26472 (.A1(W17445), .A2(W1789), .ZN(O1568));
  NANDX1 G26473 (.A1(W2868), .A2(W14487), .ZN(W18433));
  NANDX1 G26474 (.A1(W3298), .A2(I1253), .ZN(O208));
  NANDX1 G26475 (.A1(W9332), .A2(W12820), .ZN(W13410));
  NANDX1 G26476 (.A1(W23), .A2(W6695), .ZN(W7998));
  NANDX1 G26477 (.A1(W7756), .A2(W17180), .ZN(W18384));
  NANDX1 G26478 (.A1(W2268), .A2(W4389), .ZN(W4824));
  NANDX1 G26479 (.A1(I57), .A2(W5045), .ZN(W18381));
  NANDX1 G26480 (.A1(W3072), .A2(I854), .ZN(W13436));
  NANDX1 G26481 (.A1(W9323), .A2(W15037), .ZN(W18380));
  NANDX1 G26482 (.A1(W7833), .A2(W624), .ZN(W7999));
  NANDX1 G26483 (.A1(W2092), .A2(W11846), .ZN(O742));
  NANDX1 G26484 (.A1(I579), .A2(W2630), .ZN(W4827));
  NANDX1 G26485 (.A1(I455), .A2(I126), .ZN(W13435));
  NANDX1 G26486 (.A1(W3528), .A2(I1294), .ZN(W13442));
  NANDX1 G26487 (.A1(W4987), .A2(W4241), .ZN(W13443));
  NANDX1 G26488 (.A1(I240), .A2(I1763), .ZN(W13444));
  NANDX1 G26489 (.A1(W4465), .A2(W3517), .ZN(W4828));
  NANDX1 G26490 (.A1(W5583), .A2(W8237), .ZN(W13445));
  NANDX1 G26491 (.A1(W6989), .A2(W7833), .ZN(W13446));
  NANDX1 G26492 (.A1(W165), .A2(W7137), .ZN(W7997));
  NANDX1 G26493 (.A1(W4195), .A2(W3186), .ZN(W13451));
  NANDX1 G26494 (.A1(W62), .A2(I1110), .ZN(W4818));
  NANDX1 G26495 (.A1(W3689), .A2(I956), .ZN(W4814));
  NANDX1 G26496 (.A1(W6334), .A2(W7336), .ZN(W8006));
  NANDX1 G26497 (.A1(W14472), .A2(W13680), .ZN(O1559));
  NANDX1 G26498 (.A1(W4172), .A2(W4182), .ZN(W8005));
  NANDX1 G26499 (.A1(W12290), .A2(W4838), .ZN(W13430));
  NANDX1 G26500 (.A1(W1977), .A2(W1780), .ZN(W4816));
  NANDX1 G26501 (.A1(W3922), .A2(W4119), .ZN(W8004));
  NANDX1 G26502 (.A1(W7281), .A2(W17391), .ZN(W18398));
  NANDX1 G26503 (.A1(W8958), .A2(W13144), .ZN(O1747));
  NANDX1 G26504 (.A1(W11419), .A2(W2434), .ZN(W18395));
  NANDX1 G26505 (.A1(I1992), .A2(W2435), .ZN(W4820));
  NANDX1 G26506 (.A1(W8337), .A2(W3037), .ZN(W18394));
  NANDX1 G26507 (.A1(W2534), .A2(W6702), .ZN(W8003));
  NANDX1 G26508 (.A1(W1852), .A2(W10114), .ZN(W13433));
  NANDX1 G26509 (.A1(W9956), .A2(W2731), .ZN(W18388));
  NANDX1 G26510 (.A1(W9068), .A2(W12046), .ZN(W18387));
  NANDX1 G26511 (.A1(W14195), .A2(W7899), .ZN(W18385));
  NANDX1 G26512 (.A1(I1440), .A2(W3412), .ZN(W3469));
  NANDX1 G26513 (.A1(W3223), .A2(W2320), .ZN(W3461));
  NANDX1 G26514 (.A1(W12654), .A2(W1366), .ZN(O1967));
  NANDX1 G26515 (.A1(W2289), .A2(I1200), .ZN(W3462));
  NANDX1 G26516 (.A1(W8254), .A2(W5758), .ZN(W20275));
  NANDX1 G26517 (.A1(W6481), .A2(W643), .ZN(W12503));
  NANDX1 G26518 (.A1(W7074), .A2(W1020), .ZN(W12504));
  NANDX1 G26519 (.A1(I1256), .A2(W3053), .ZN(W3467));
  NANDX1 G26520 (.A1(W9136), .A2(W7040), .ZN(W12505));
  NANDX1 G26521 (.A1(W9999), .A2(W8094), .ZN(W12506));
  NANDX1 G26522 (.A1(W828), .A2(W3144), .ZN(W3460));
  NANDX1 G26523 (.A1(I488), .A2(W2579), .ZN(W3470));
  NANDX1 G26524 (.A1(W5366), .A2(W6072), .ZN(W8598));
  NANDX1 G26525 (.A1(W4511), .A2(W7466), .ZN(W8595));
  NANDX1 G26526 (.A1(I1843), .A2(W2448), .ZN(W3471));
  NANDX1 G26527 (.A1(W3306), .A2(I1698), .ZN(W3473));
  NANDX1 G26528 (.A1(W37), .A2(W2188), .ZN(W8594));
  NANDX1 G26529 (.A1(I96), .A2(I1326), .ZN(W3474));
  NANDX1 G26530 (.A1(W1270), .A2(I1872), .ZN(W3475));
  NANDX1 G26531 (.A1(I430), .A2(I368), .ZN(W3451));
  NANDX1 G26532 (.A1(W15428), .A2(W6624), .ZN(W20294));
  NANDX1 G26533 (.A1(W11178), .A2(W3180), .ZN(W20293));
  NANDX1 G26534 (.A1(W11799), .A2(W20228), .ZN(W20292));
  NANDX1 G26535 (.A1(I1940), .A2(W1516), .ZN(W3447));
  NANDX1 G26536 (.A1(W11189), .A2(W12288), .ZN(W12497));
  NANDX1 G26537 (.A1(W8602), .A2(W1942), .ZN(W20291));
  NANDX1 G26538 (.A1(W2289), .A2(W2597), .ZN(W3449));
  NANDX1 G26539 (.A1(W329), .A2(W7403), .ZN(W20289));
  NANDX1 G26540 (.A1(W12006), .A2(I1940), .ZN(W20263));
  NANDX1 G26541 (.A1(I114), .A2(W9358), .ZN(W12498));
  NANDX1 G26542 (.A1(I1147), .A2(W483), .ZN(W3453));
  NANDX1 G26543 (.A1(W10673), .A2(W3693), .ZN(O1969));
  NANDX1 G26544 (.A1(W1607), .A2(W268), .ZN(W3454));
  NANDX1 G26545 (.A1(W19025), .A2(W13011), .ZN(W20281));
  NANDX1 G26546 (.A1(I38), .A2(W2270), .ZN(W3457));
  NANDX1 G26547 (.A1(W2179), .A2(W11396), .ZN(W12502));
  NANDX1 G26548 (.A1(W4256), .A2(W2027), .ZN(W20279));
  NANDX1 G26549 (.A1(W2522), .A2(W2766), .ZN(W8586));
  NANDX1 G26550 (.A1(W16927), .A2(W7232), .ZN(W20240));
  NANDX1 G26551 (.A1(I1888), .A2(W8331), .ZN(O1958));
  NANDX1 G26552 (.A1(W5877), .A2(W2928), .ZN(W8588));
  NANDX1 G26553 (.A1(W6586), .A2(W12652), .ZN(W20238));
  NANDX1 G26554 (.A1(W1697), .A2(W20138), .ZN(W20237));
  NANDX1 G26555 (.A1(I1134), .A2(W1837), .ZN(W12522));
  NANDX1 G26556 (.A1(W15169), .A2(W8580), .ZN(W20233));
  NANDX1 G26557 (.A1(W8976), .A2(W17892), .ZN(W20232));
  NANDX1 G26558 (.A1(W6051), .A2(W339), .ZN(W12526));
  NANDX1 G26559 (.A1(W2324), .A2(W10627), .ZN(W12520));
  NANDX1 G26560 (.A1(W3238), .A2(I1029), .ZN(W3499));
  NANDX1 G26561 (.A1(W848), .A2(W3371), .ZN(W8584));
  NANDX1 G26562 (.A1(W433), .A2(W8376), .ZN(W8578));
  NANDX1 G26563 (.A1(I1477), .A2(W775), .ZN(W12528));
  NANDX1 G26564 (.A1(W2125), .A2(W78), .ZN(W3503));
  NANDX1 G26565 (.A1(W459), .A2(W769), .ZN(W12532));
  NANDX1 G26566 (.A1(W4983), .A2(W6352), .ZN(W12533));
  NANDX1 G26567 (.A1(W10919), .A2(W9675), .ZN(W20222));
  NANDX1 G26568 (.A1(W1113), .A2(W1869), .ZN(W3482));
  NANDX1 G26569 (.A1(I371), .A2(W2456), .ZN(W20261));
  NANDX1 G26570 (.A1(W20068), .A2(W13311), .ZN(W20260));
  NANDX1 G26571 (.A1(W4540), .A2(W8211), .ZN(W12508));
  NANDX1 G26572 (.A1(I1518), .A2(W1348), .ZN(W3479));
  NANDX1 G26573 (.A1(W5552), .A2(W1646), .ZN(W12509));
  NANDX1 G26574 (.A1(W43), .A2(W4986), .ZN(W12510));
  NANDX1 G26575 (.A1(I1749), .A2(W10450), .ZN(W12511));
  NANDX1 G26576 (.A1(W5696), .A2(W5272), .ZN(W12512));
  NANDX1 G26577 (.A1(W12773), .A2(W15188), .ZN(O1970));
  NANDX1 G26578 (.A1(W5740), .A2(W6295), .ZN(O1963));
  NANDX1 G26579 (.A1(W8268), .A2(I1066), .ZN(O605));
  NANDX1 G26580 (.A1(W9029), .A2(W2220), .ZN(W12519));
  NANDX1 G26581 (.A1(W5406), .A2(W3750), .ZN(W8591));
  NANDX1 G26582 (.A1(I630), .A2(W291), .ZN(W3484));
  NANDX1 G26583 (.A1(I124), .A2(W2648), .ZN(W3487));
  NANDX1 G26584 (.A1(I161), .A2(W10560), .ZN(W20247));
  NANDX1 G26585 (.A1(W4056), .A2(W18489), .ZN(O1959));
  NANDX1 G26586 (.A1(I1172), .A2(W1455), .ZN(W3404));
  NANDX1 G26587 (.A1(W11870), .A2(W8399), .ZN(W12467));
  NANDX1 G26588 (.A1(I351), .A2(W2677), .ZN(W3399));
  NANDX1 G26589 (.A1(W3312), .A2(W19894), .ZN(W20358));
  NANDX1 G26590 (.A1(W18005), .A2(W13417), .ZN(W20357));
  NANDX1 G26591 (.A1(W7453), .A2(W8379), .ZN(W8621));
  NANDX1 G26592 (.A1(W4948), .A2(W1389), .ZN(O1985));
  NANDX1 G26593 (.A1(W2793), .A2(I194), .ZN(W3401));
  NANDX1 G26594 (.A1(I1267), .A2(W6592), .ZN(W12470));
  NANDX1 G26595 (.A1(W6304), .A2(W3752), .ZN(O1980));
  NANDX1 G26596 (.A1(W10352), .A2(W8776), .ZN(W20364));
  NANDX1 G26597 (.A1(W19026), .A2(W15015), .ZN(W20341));
  NANDX1 G26598 (.A1(W7624), .A2(W1185), .ZN(W8619));
  NANDX1 G26599 (.A1(W4735), .A2(W7771), .ZN(W8617));
  NANDX1 G26600 (.A1(W6317), .A2(W6084), .ZN(W12475));
  NANDX1 G26601 (.A1(W17501), .A2(W3703), .ZN(O1977));
  NANDX1 G26602 (.A1(W3010), .A2(I1332), .ZN(W3411));
  NANDX1 G26603 (.A1(W59), .A2(I259), .ZN(W3412));
  NANDX1 G26604 (.A1(W7835), .A2(W2090), .ZN(W8616));
  NANDX1 G26605 (.A1(W1136), .A2(W1134), .ZN(W8632));
  NANDX1 G26606 (.A1(W1813), .A2(W8185), .ZN(W12456));
  NANDX1 G26607 (.A1(W3478), .A2(W5575), .ZN(W12457));
  NANDX1 G26608 (.A1(I1052), .A2(W1718), .ZN(W3377));
  NANDX1 G26609 (.A1(W2271), .A2(W1508), .ZN(W3378));
  NANDX1 G26610 (.A1(W2742), .A2(W8393), .ZN(W12459));
  NANDX1 G26611 (.A1(W19666), .A2(W5294), .ZN(W20383));
  NANDX1 G26612 (.A1(W1485), .A2(W1765), .ZN(W3382));
  NANDX1 G26613 (.A1(I574), .A2(W2676), .ZN(W3384));
  NANDX1 G26614 (.A1(I527), .A2(I259), .ZN(W12476));
  NANDX1 G26615 (.A1(I243), .A2(W1014), .ZN(W3386));
  NANDX1 G26616 (.A1(W8124), .A2(W4353), .ZN(W8629));
  NANDX1 G26617 (.A1(W6020), .A2(W8258), .ZN(W8627));
  NANDX1 G26618 (.A1(W18245), .A2(W4101), .ZN(W20376));
  NANDX1 G26619 (.A1(W4371), .A2(W3100), .ZN(W8622));
  NANDX1 G26620 (.A1(W3015), .A2(I1136), .ZN(W3394));
  NANDX1 G26621 (.A1(W1783), .A2(W2565), .ZN(W3395));
  NANDX1 G26622 (.A1(W18535), .A2(W3592), .ZN(W20365));
  NANDX1 G26623 (.A1(W7031), .A2(W12424), .ZN(W20305));
  NANDX1 G26624 (.A1(I600), .A2(W3471), .ZN(W20313));
  NANDX1 G26625 (.A1(W6319), .A2(W7119), .ZN(W8608));
  NANDX1 G26626 (.A1(I1233), .A2(W2227), .ZN(W3436));
  NANDX1 G26627 (.A1(W1638), .A2(W2852), .ZN(W3437));
  NANDX1 G26628 (.A1(W11731), .A2(W10597), .ZN(W12489));
  NANDX1 G26629 (.A1(W13063), .A2(W17538), .ZN(W20307));
  NANDX1 G26630 (.A1(W5246), .A2(W5573), .ZN(W8605));
  NANDX1 G26631 (.A1(W1514), .A2(W1702), .ZN(W3440));
  NANDX1 G26632 (.A1(I800), .A2(W3047), .ZN(W3433));
  NANDX1 G26633 (.A1(W13771), .A2(W3348), .ZN(W20303));
  NANDX1 G26634 (.A1(W12692), .A2(W7823), .ZN(W20301));
  NANDX1 G26635 (.A1(W3265), .A2(I1148), .ZN(W3444));
  NANDX1 G26636 (.A1(W18074), .A2(W5943), .ZN(W20300));
  NANDX1 G26637 (.A1(W12127), .A2(W11963), .ZN(W20298));
  NANDX1 G26638 (.A1(W9058), .A2(W11936), .ZN(W12493));
  NANDX1 G26639 (.A1(W1259), .A2(W2380), .ZN(W3445));
  NANDX1 G26640 (.A1(I1654), .A2(W1247), .ZN(W12496));
  NANDX1 G26641 (.A1(W17651), .A2(W7024), .ZN(W20322));
  NANDX1 G26642 (.A1(W7590), .A2(W1372), .ZN(W12477));
  NANDX1 G26643 (.A1(W1874), .A2(W7052), .ZN(W20330));
  NANDX1 G26644 (.A1(W1648), .A2(W1264), .ZN(W3417));
  NANDX1 G26645 (.A1(W4293), .A2(W12730), .ZN(W20328));
  NANDX1 G26646 (.A1(I792), .A2(W7139), .ZN(W12478));
  NANDX1 G26647 (.A1(I1444), .A2(W2636), .ZN(W8614));
  NANDX1 G26648 (.A1(W14901), .A2(W3357), .ZN(W20326));
  NANDX1 G26649 (.A1(W11836), .A2(W17903), .ZN(W20324));
  NANDX1 G26650 (.A1(W7495), .A2(I1535), .ZN(W8575));
  NANDX1 G26651 (.A1(W10059), .A2(W1427), .ZN(W12480));
  NANDX1 G26652 (.A1(W295), .A2(W3208), .ZN(W3420));
  NANDX1 G26653 (.A1(W17802), .A2(W7860), .ZN(W20321));
  NANDX1 G26654 (.A1(I1193), .A2(W2448), .ZN(W3424));
  NANDX1 G26655 (.A1(W15681), .A2(W3663), .ZN(O1975));
  NANDX1 G26656 (.A1(I567), .A2(W644), .ZN(W12482));
  NANDX1 G26657 (.A1(W8426), .A2(W6440), .ZN(W8610));
  NANDX1 G26658 (.A1(W80), .A2(I820), .ZN(W3428));
  NANDX1 G26659 (.A1(W15059), .A2(W113), .ZN(W20099));
  NANDX1 G26660 (.A1(W1976), .A2(W266), .ZN(W12582));
  NANDX1 G26661 (.A1(W11760), .A2(W421), .ZN(W20105));
  NANDX1 G26662 (.A1(W1558), .A2(I237), .ZN(W3594));
  NANDX1 G26663 (.A1(W2592), .A2(W7811), .ZN(W8541));
  NANDX1 G26664 (.A1(W11249), .A2(W2304), .ZN(W20104));
  NANDX1 G26665 (.A1(W6), .A2(W2044), .ZN(W3595));
  NANDX1 G26666 (.A1(I18), .A2(W4580), .ZN(W12586));
  NANDX1 G26667 (.A1(W355), .A2(W9091), .ZN(W12588));
  NANDX1 G26668 (.A1(W1700), .A2(I1015), .ZN(W12590));
  NANDX1 G26669 (.A1(W7048), .A2(W6987), .ZN(W20111));
  NANDX1 G26670 (.A1(W284), .A2(W2986), .ZN(W3602));
  NANDX1 G26671 (.A1(W2347), .A2(W5795), .ZN(O235));
  NANDX1 G26672 (.A1(W16501), .A2(W11369), .ZN(O1926));
  NANDX1 G26673 (.A1(W2307), .A2(W3169), .ZN(W3604));
  NANDX1 G26674 (.A1(W6250), .A2(W17701), .ZN(W20095));
  NANDX1 G26675 (.A1(W1880), .A2(W135), .ZN(W3607));
  NANDX1 G26676 (.A1(W11210), .A2(W6383), .ZN(W20091));
  NANDX1 G26677 (.A1(W6237), .A2(W9593), .ZN(W12595));
  NANDX1 G26678 (.A1(W2620), .A2(I888), .ZN(O39));
  NANDX1 G26679 (.A1(W14352), .A2(I1033), .ZN(O1934));
  NANDX1 G26680 (.A1(W15523), .A2(W19673), .ZN(W20126));
  NANDX1 G26681 (.A1(W19023), .A2(W19813), .ZN(W20125));
  NANDX1 G26682 (.A1(W2778), .A2(W314), .ZN(W3577));
  NANDX1 G26683 (.A1(W4089), .A2(W20075), .ZN(O1932));
  NANDX1 G26684 (.A1(W16647), .A2(W8934), .ZN(W20118));
  NANDX1 G26685 (.A1(W9811), .A2(W4521), .ZN(W12574));
  NANDX1 G26686 (.A1(W2872), .A2(I180), .ZN(W3583));
  NANDX1 G26687 (.A1(W2592), .A2(W7916), .ZN(W12596));
  NANDX1 G26688 (.A1(W2240), .A2(W6397), .ZN(O616));
  NANDX1 G26689 (.A1(W2549), .A2(W7890), .ZN(W8548));
  NANDX1 G26690 (.A1(I1224), .A2(W1756), .ZN(W12577));
  NANDX1 G26691 (.A1(W4752), .A2(W2136), .ZN(O618));
  NANDX1 G26692 (.A1(W2324), .A2(W3054), .ZN(W8543));
  NANDX1 G26693 (.A1(W1403), .A2(W3583), .ZN(W3587));
  NANDX1 G26694 (.A1(W2627), .A2(I1703), .ZN(W3591));
  NANDX1 G26695 (.A1(W7535), .A2(W1492), .ZN(W12580));
  NANDX1 G26696 (.A1(W10607), .A2(W2382), .ZN(W20058));
  NANDX1 G26697 (.A1(W5236), .A2(W11139), .ZN(W12611));
  NANDX1 G26698 (.A1(W9229), .A2(W597), .ZN(W12612));
  NANDX1 G26699 (.A1(W4483), .A2(W3301), .ZN(W8528));
  NANDX1 G26700 (.A1(I953), .A2(W42), .ZN(W3629));
  NANDX1 G26701 (.A1(W11571), .A2(W4991), .ZN(W12616));
  NANDX1 G26702 (.A1(I1564), .A2(W2850), .ZN(W3636));
  NANDX1 G26703 (.A1(W11374), .A2(W271), .ZN(W20062));
  NANDX1 G26704 (.A1(W13411), .A2(W17291), .ZN(W20059));
  NANDX1 G26705 (.A1(W8508), .A2(W1953), .ZN(W12609));
  NANDX1 G26706 (.A1(W16450), .A2(W15071), .ZN(O1918));
  NANDX1 G26707 (.A1(W233), .A2(W105), .ZN(W8526));
  NANDX1 G26708 (.A1(I1842), .A2(W3427), .ZN(W20054));
  NANDX1 G26709 (.A1(W6686), .A2(W8113), .ZN(W8520));
  NANDX1 G26710 (.A1(W17121), .A2(W7926), .ZN(O1917));
  NANDX1 G26711 (.A1(I235), .A2(I154), .ZN(W3642));
  NANDX1 G26712 (.A1(W13078), .A2(W4410), .ZN(W20050));
  NANDX1 G26713 (.A1(W2170), .A2(W536), .ZN(W3645));
  NANDX1 G26714 (.A1(W9081), .A2(W8759), .ZN(W12603));
  NANDX1 G26715 (.A1(W11088), .A2(W2985), .ZN(W12599));
  NANDX1 G26716 (.A1(W3406), .A2(W6799), .ZN(O621));
  NANDX1 G26717 (.A1(W3813), .A2(W6033), .ZN(W12601));
  NANDX1 G26718 (.A1(W3102), .A2(I1281), .ZN(W3613));
  NANDX1 G26719 (.A1(W13916), .A2(W9346), .ZN(W20086));
  NANDX1 G26720 (.A1(W551), .A2(W4120), .ZN(W8532));
  NANDX1 G26721 (.A1(W2143), .A2(W817), .ZN(W3614));
  NANDX1 G26722 (.A1(W9214), .A2(W8427), .ZN(W20084));
  NANDX1 G26723 (.A1(W17417), .A2(W2645), .ZN(W20129));
  NANDX1 G26724 (.A1(W3625), .A2(W10135), .ZN(W12605));
  NANDX1 G26725 (.A1(W2421), .A2(W1197), .ZN(W3619));
  NANDX1 G26726 (.A1(W7798), .A2(W11653), .ZN(O622));
  NANDX1 G26727 (.A1(I349), .A2(W3059), .ZN(W3622));
  NANDX1 G26728 (.A1(W735), .A2(W9489), .ZN(W20078));
  NANDX1 G26729 (.A1(W4909), .A2(W14536), .ZN(W20076));
  NANDX1 G26730 (.A1(W1430), .A2(W13801), .ZN(W20074));
  NANDX1 G26731 (.A1(I1212), .A2(W7540), .ZN(W8530));
  NANDX1 G26732 (.A1(W4913), .A2(W8095), .ZN(W8570));
  NANDX1 G26733 (.A1(W951), .A2(I1518), .ZN(W3520));
  NANDX1 G26734 (.A1(I816), .A2(I1509), .ZN(W3524));
  NANDX1 G26735 (.A1(W2956), .A2(I182), .ZN(W3527));
  NANDX1 G26736 (.A1(W19776), .A2(W15120), .ZN(W20194));
  NANDX1 G26737 (.A1(W11997), .A2(W2560), .ZN(O1949));
  NANDX1 G26738 (.A1(W2046), .A2(W2828), .ZN(W3528));
  NANDX1 G26739 (.A1(W1705), .A2(W3980), .ZN(W20190));
  NANDX1 G26740 (.A1(W138), .A2(I344), .ZN(W8572));
  NANDX1 G26741 (.A1(W1840), .A2(W406), .ZN(W3531));
  NANDX1 G26742 (.A1(W3358), .A2(I1876), .ZN(O1951));
  NANDX1 G26743 (.A1(W11051), .A2(W9308), .ZN(W12543));
  NANDX1 G26744 (.A1(W279), .A2(W82), .ZN(W3535));
  NANDX1 G26745 (.A1(W2964), .A2(W1806), .ZN(W3537));
  NANDX1 G26746 (.A1(W3826), .A2(I659), .ZN(W20182));
  NANDX1 G26747 (.A1(I198), .A2(W1217), .ZN(W3538));
  NANDX1 G26748 (.A1(W1532), .A2(I1887), .ZN(W3539));
  NANDX1 G26749 (.A1(W7570), .A2(I1831), .ZN(W8569));
  NANDX1 G26750 (.A1(W15851), .A2(I301), .ZN(O1948));
  NANDX1 G26751 (.A1(I846), .A2(W1085), .ZN(W3512));
  NANDX1 G26752 (.A1(W15000), .A2(W15730), .ZN(W20217));
  NANDX1 G26753 (.A1(W463), .A2(I777), .ZN(W3507));
  NANDX1 G26754 (.A1(W4381), .A2(W8035), .ZN(W20214));
  NANDX1 G26755 (.A1(W7555), .A2(W8724), .ZN(W20213));
  NANDX1 G26756 (.A1(W1260), .A2(W5323), .ZN(W12535));
  NANDX1 G26757 (.A1(W11392), .A2(W529), .ZN(W20210));
  NANDX1 G26758 (.A1(W2734), .A2(W2135), .ZN(W3509));
  NANDX1 G26759 (.A1(W1879), .A2(W2409), .ZN(W3510));
  NANDX1 G26760 (.A1(W12605), .A2(W11162), .ZN(W20177));
  NANDX1 G26761 (.A1(W16408), .A2(W2783), .ZN(W20206));
  NANDX1 G26762 (.A1(W19209), .A2(W15148), .ZN(W20204));
  NANDX1 G26763 (.A1(W8029), .A2(W7155), .ZN(W8574));
  NANDX1 G26764 (.A1(W7366), .A2(W3790), .ZN(W12538));
  NANDX1 G26765 (.A1(W12969), .A2(W1341), .ZN(O1952));
  NANDX1 G26766 (.A1(W17425), .A2(W6416), .ZN(W20200));
  NANDX1 G26767 (.A1(W2863), .A2(W1883), .ZN(W3517));
  NANDX1 G26768 (.A1(W1843), .A2(W1654), .ZN(W3518));
  NANDX1 G26769 (.A1(W8651), .A2(W9824), .ZN(O1940));
  NANDX1 G26770 (.A1(W2667), .A2(W4661), .ZN(O612));
  NANDX1 G26771 (.A1(I1202), .A2(W5845), .ZN(W12560));
  NANDX1 G26772 (.A1(W3631), .A2(W10900), .ZN(W20152));
  NANDX1 G26773 (.A1(W194), .A2(W12389), .ZN(W12561));
  NANDX1 G26774 (.A1(W17899), .A2(W11521), .ZN(W20151));
  NANDX1 G26775 (.A1(W609), .A2(W836), .ZN(W3566));
  NANDX1 G26776 (.A1(W2640), .A2(W819), .ZN(W3567));
  NANDX1 G26777 (.A1(W10200), .A2(W8840), .ZN(W12564));
  NANDX1 G26778 (.A1(W7411), .A2(W8969), .ZN(W12556));
  NANDX1 G26779 (.A1(W12021), .A2(W5598), .ZN(W20146));
  NANDX1 G26780 (.A1(W1653), .A2(W422), .ZN(W3571));
  NANDX1 G26781 (.A1(W14650), .A2(W13905), .ZN(W20142));
  NANDX1 G26782 (.A1(W4667), .A2(W2514), .ZN(W8561));
  NANDX1 G26783 (.A1(I948), .A2(W2656), .ZN(W8559));
  NANDX1 G26784 (.A1(I1604), .A2(W13996), .ZN(W20137));
  NANDX1 G26785 (.A1(W231), .A2(W5354), .ZN(W12569));
  NANDX1 G26786 (.A1(W5333), .A2(W455), .ZN(W8557));
  NANDX1 G26787 (.A1(I1025), .A2(I870), .ZN(W3555));
  NANDX1 G26788 (.A1(W5478), .A2(W5283), .ZN(W8564));
  NANDX1 G26789 (.A1(W9404), .A2(W8752), .ZN(W20176));
  NANDX1 G26790 (.A1(W8362), .A2(W2721), .ZN(W12549));
  NANDX1 G26791 (.A1(I1562), .A2(W6832), .ZN(O1946));
  NANDX1 G26792 (.A1(W8992), .A2(W3066), .ZN(W12550));
  NANDX1 G26793 (.A1(I138), .A2(I1915), .ZN(W3553));
  NANDX1 G26794 (.A1(W15535), .A2(I224), .ZN(W20167));
  NANDX1 G26795 (.A1(W459), .A2(I840), .ZN(O610));
  NANDX1 G26796 (.A1(W4105), .A2(W5842), .ZN(W12454));
  NANDX1 G26797 (.A1(W11215), .A2(W2096), .ZN(W12552));
  NANDX1 G26798 (.A1(W3921), .A2(W16559), .ZN(W20163));
  NANDX1 G26799 (.A1(W2297), .A2(W876), .ZN(W3559));
  NANDX1 G26800 (.A1(W1929), .A2(W1405), .ZN(W3560));
  NANDX1 G26801 (.A1(W9840), .A2(W2404), .ZN(W12553));
  NANDX1 G26802 (.A1(W10913), .A2(W9087), .ZN(W12554));
  NANDX1 G26803 (.A1(W8422), .A2(W1672), .ZN(O1942));
  NANDX1 G26804 (.A1(W3772), .A2(W12613), .ZN(W20156));
  NANDX1 G26805 (.A1(W18197), .A2(I1165), .ZN(W20625));
  NANDX1 G26806 (.A1(W13464), .A2(W10946), .ZN(W20636));
  NANDX1 G26807 (.A1(W9743), .A2(W4263), .ZN(W20634));
  NANDX1 G26808 (.A1(W15778), .A2(W6831), .ZN(W20631));
  NANDX1 G26809 (.A1(W19378), .A2(W14027), .ZN(W20630));
  NANDX1 G26810 (.A1(I1005), .A2(W1286), .ZN(W8729));
  NANDX1 G26811 (.A1(W3634), .A2(W2352), .ZN(W8727));
  NANDX1 G26812 (.A1(I1465), .A2(I741), .ZN(W3205));
  NANDX1 G26813 (.A1(I1988), .A2(W3065), .ZN(W3206));
  NANDX1 G26814 (.A1(W615), .A2(W1366), .ZN(W12360));
  NANDX1 G26815 (.A1(W6706), .A2(W165), .ZN(W8732));
  NANDX1 G26816 (.A1(W2182), .A2(I344), .ZN(W3207));
  NANDX1 G26817 (.A1(W603), .A2(W236), .ZN(W3208));
  NANDX1 G26818 (.A1(W9707), .A2(W9370), .ZN(W20623));
  NANDX1 G26819 (.A1(W3008), .A2(W2609), .ZN(W3211));
  NANDX1 G26820 (.A1(W19208), .A2(W10085), .ZN(W20619));
  NANDX1 G26821 (.A1(W19930), .A2(W3246), .ZN(W20618));
  NANDX1 G26822 (.A1(W660), .A2(W1236), .ZN(W3212));
  NANDX1 G26823 (.A1(I672), .A2(W3198), .ZN(W3214));
  NANDX1 G26824 (.A1(I498), .A2(I352), .ZN(W3193));
  NANDX1 G26825 (.A1(W14192), .A2(W18966), .ZN(W20661));
  NANDX1 G26826 (.A1(W996), .A2(W951), .ZN(W3187));
  NANDX1 G26827 (.A1(W890), .A2(I898), .ZN(O30));
  NANDX1 G26828 (.A1(W14057), .A2(W6093), .ZN(W20655));
  NANDX1 G26829 (.A1(W12035), .A2(W11373), .ZN(W20653));
  NANDX1 G26830 (.A1(W2674), .A2(W2107), .ZN(W3191));
  NANDX1 G26831 (.A1(W11770), .A2(W19466), .ZN(W20652));
  NANDX1 G26832 (.A1(W2133), .A2(W401), .ZN(W3192));
  NANDX1 G26833 (.A1(W20530), .A2(W20226), .ZN(W20614));
  NANDX1 G26834 (.A1(W11465), .A2(W5876), .ZN(W12355));
  NANDX1 G26835 (.A1(W9535), .A2(W7831), .ZN(W20648));
  NANDX1 G26836 (.A1(W5445), .A2(W5970), .ZN(W20646));
  NANDX1 G26837 (.A1(W1409), .A2(I332), .ZN(W3195));
  NANDX1 G26838 (.A1(W5394), .A2(I630), .ZN(W20643));
  NANDX1 G26839 (.A1(I440), .A2(W3011), .ZN(W3196));
  NANDX1 G26840 (.A1(I1760), .A2(W6816), .ZN(W8738));
  NANDX1 G26841 (.A1(W1745), .A2(W3589), .ZN(W8735));
  NANDX1 G26842 (.A1(W5256), .A2(W6936), .ZN(W8704));
  NANDX1 G26843 (.A1(W9891), .A2(W7936), .ZN(W20595));
  NANDX1 G26844 (.A1(I796), .A2(W13547), .ZN(W20592));
  NANDX1 G26845 (.A1(W17988), .A2(W6395), .ZN(O2040));
  NANDX1 G26846 (.A1(W5370), .A2(W13192), .ZN(W20590));
  NANDX1 G26847 (.A1(W2846), .A2(W17934), .ZN(W20589));
  NANDX1 G26848 (.A1(I1360), .A2(W1324), .ZN(W3233));
  NANDX1 G26849 (.A1(W7011), .A2(W8905), .ZN(W20581));
  NANDX1 G26850 (.A1(W2254), .A2(W1335), .ZN(O596));
  NANDX1 G26851 (.A1(W5445), .A2(W11882), .ZN(W12370));
  NANDX1 G26852 (.A1(W14340), .A2(W3156), .ZN(W20574));
  NANDX1 G26853 (.A1(W7648), .A2(W5940), .ZN(W8703));
  NANDX1 G26854 (.A1(W15127), .A2(W218), .ZN(O2035));
  NANDX1 G26855 (.A1(W3095), .A2(W2052), .ZN(W3241));
  NANDX1 G26856 (.A1(W14372), .A2(W18168), .ZN(W20570));
  NANDX1 G26857 (.A1(W18280), .A2(W3613), .ZN(W20569));
  NANDX1 G26858 (.A1(W2288), .A2(W2935), .ZN(W12382));
  NANDX1 G26859 (.A1(I1716), .A2(W1997), .ZN(W8700));
  NANDX1 G26860 (.A1(I694), .A2(W739), .ZN(W3221));
  NANDX1 G26861 (.A1(W666), .A2(W2335), .ZN(W12367));
  NANDX1 G26862 (.A1(I896), .A2(W1811), .ZN(W3215));
  NANDX1 G26863 (.A1(W12108), .A2(W2402), .ZN(W20609));
  NANDX1 G26864 (.A1(W4750), .A2(W1785), .ZN(W8720));
  NANDX1 G26865 (.A1(W2726), .A2(W2960), .ZN(W3216));
  NANDX1 G26866 (.A1(W10109), .A2(I1630), .ZN(W20607));
  NANDX1 G26867 (.A1(W2350), .A2(W2095), .ZN(W3220));
  NANDX1 G26868 (.A1(W16334), .A2(W3003), .ZN(W20606));
  NANDX1 G26869 (.A1(W4364), .A2(W8000), .ZN(W12352));
  NANDX1 G26870 (.A1(I860), .A2(W2522), .ZN(W3222));
  NANDX1 G26871 (.A1(I791), .A2(W2723), .ZN(W3224));
  NANDX1 G26872 (.A1(W11964), .A2(W17114), .ZN(W20601));
  NANDX1 G26873 (.A1(W20398), .A2(W13665), .ZN(W20600));
  NANDX1 G26874 (.A1(W4412), .A2(W8094), .ZN(W8712));
  NANDX1 G26875 (.A1(W5193), .A2(W5907), .ZN(W20598));
  NANDX1 G26876 (.A1(W16914), .A2(W9779), .ZN(W20597));
  NANDX1 G26877 (.A1(W2451), .A2(W590), .ZN(W3230));
  NANDX1 G26878 (.A1(W2008), .A2(W18859), .ZN(O2065));
  NANDX1 G26879 (.A1(W6799), .A2(W85), .ZN(W8774));
  NANDX1 G26880 (.A1(W3435), .A2(W8818), .ZN(W20728));
  NANDX1 G26881 (.A1(W11597), .A2(W8274), .ZN(W20725));
  NANDX1 G26882 (.A1(W7809), .A2(W4035), .ZN(W12311));
  NANDX1 G26883 (.A1(W406), .A2(W1352), .ZN(W3142));
  NANDX1 G26884 (.A1(W827), .A2(W983), .ZN(W3146));
  NANDX1 G26885 (.A1(W2123), .A2(W7078), .ZN(W12312));
  NANDX1 G26886 (.A1(I320), .A2(I55), .ZN(W3148));
  NANDX1 G26887 (.A1(W19104), .A2(W11484), .ZN(W20719));
  NANDX1 G26888 (.A1(W8837), .A2(W6579), .ZN(W20730));
  NANDX1 G26889 (.A1(W7713), .A2(W4221), .ZN(W8772));
  NANDX1 G26890 (.A1(W1455), .A2(W7433), .ZN(W8768));
  NANDX1 G26891 (.A1(W13838), .A2(W2809), .ZN(W20713));
  NANDX1 G26892 (.A1(W479), .A2(I1110), .ZN(W3155));
  NANDX1 G26893 (.A1(W3842), .A2(W3650), .ZN(W20710));
  NANDX1 G26894 (.A1(I947), .A2(W3097), .ZN(W8764));
  NANDX1 G26895 (.A1(W13471), .A2(W519), .ZN(W20709));
  NANDX1 G26896 (.A1(W6091), .A2(W16412), .ZN(O2062));
  NANDX1 G26897 (.A1(W19463), .A2(W5195), .ZN(O2070));
  NANDX1 G26898 (.A1(W2564), .A2(W1827), .ZN(W12298));
  NANDX1 G26899 (.A1(W348), .A2(W236), .ZN(W3129));
  NANDX1 G26900 (.A1(W2815), .A2(I1225), .ZN(O2072));
  NANDX1 G26901 (.A1(W9903), .A2(W8849), .ZN(W20749));
  NANDX1 G26902 (.A1(W8217), .A2(W3172), .ZN(W8781));
  NANDX1 G26903 (.A1(W17896), .A2(W5769), .ZN(W20747));
  NANDX1 G26904 (.A1(W8013), .A2(W10243), .ZN(O2071));
  NANDX1 G26905 (.A1(W5184), .A2(W11207), .ZN(W12300));
  NANDX1 G26906 (.A1(W1469), .A2(W1326), .ZN(W3160));
  NANDX1 G26907 (.A1(W4238), .A2(W8265), .ZN(W8780));
  NANDX1 G26908 (.A1(W4404), .A2(W8550), .ZN(W20739));
  NANDX1 G26909 (.A1(W4901), .A2(W16876), .ZN(W20736));
  NANDX1 G26910 (.A1(W5097), .A2(W19327), .ZN(W20735));
  NANDX1 G26911 (.A1(W16375), .A2(W5204), .ZN(W20734));
  NANDX1 G26912 (.A1(W1508), .A2(I975), .ZN(W3140));
  NANDX1 G26913 (.A1(W3965), .A2(W9487), .ZN(W20733));
  NANDX1 G26914 (.A1(I588), .A2(W8668), .ZN(W20732));
  NANDX1 G26915 (.A1(W10747), .A2(W10426), .ZN(W12346));
  NANDX1 G26916 (.A1(W2708), .A2(I846), .ZN(W12333));
  NANDX1 G26917 (.A1(W9842), .A2(W4213), .ZN(W12337));
  NANDX1 G26918 (.A1(I1650), .A2(W2383), .ZN(W8749));
  NANDX1 G26919 (.A1(W14514), .A2(W9908), .ZN(W20681));
  NANDX1 G26920 (.A1(W5116), .A2(I326), .ZN(W8748));
  NANDX1 G26921 (.A1(W13078), .A2(W16704), .ZN(W20680));
  NANDX1 G26922 (.A1(W20110), .A2(W5240), .ZN(W20679));
  NANDX1 G26923 (.A1(I1471), .A2(I863), .ZN(W3177));
  NANDX1 G26924 (.A1(W16773), .A2(W4399), .ZN(W20683));
  NANDX1 G26925 (.A1(W14887), .A2(W20623), .ZN(W20674));
  NANDX1 G26926 (.A1(W6332), .A2(W6063), .ZN(W8743));
  NANDX1 G26927 (.A1(W10725), .A2(W1684), .ZN(W12349));
  NANDX1 G26928 (.A1(I1640), .A2(I766), .ZN(W3179));
  NANDX1 G26929 (.A1(W9868), .A2(W3806), .ZN(W20666));
  NANDX1 G26930 (.A1(W5672), .A2(I396), .ZN(W20665));
  NANDX1 G26931 (.A1(W541), .A2(W1887), .ZN(W3181));
  NANDX1 G26932 (.A1(W1405), .A2(W555), .ZN(W3182));
  NANDX1 G26933 (.A1(W18517), .A2(I1361), .ZN(W20695));
  NANDX1 G26934 (.A1(W14549), .A2(W2897), .ZN(O2061));
  NANDX1 G26935 (.A1(I1399), .A2(W1211), .ZN(W3161));
  NANDX1 G26936 (.A1(W2033), .A2(I136), .ZN(W12317));
  NANDX1 G26937 (.A1(I1719), .A2(W5870), .ZN(O592));
  NANDX1 G26938 (.A1(W3978), .A2(W16023), .ZN(O2060));
  NANDX1 G26939 (.A1(W947), .A2(W2277), .ZN(W8757));
  NANDX1 G26940 (.A1(W6928), .A2(W2722), .ZN(W20697));
  NANDX1 G26941 (.A1(I902), .A2(I1471), .ZN(W3162));
  NANDX1 G26942 (.A1(W231), .A2(W2917), .ZN(W3245));
  NANDX1 G26943 (.A1(W15339), .A2(W5348), .ZN(W20694));
  NANDX1 G26944 (.A1(W1275), .A2(I1429), .ZN(W3165));
  NANDX1 G26945 (.A1(W7862), .A2(W3309), .ZN(O244));
  NANDX1 G26946 (.A1(W3339), .A2(W3047), .ZN(W12328));
  NANDX1 G26947 (.A1(W8494), .A2(W19447), .ZN(W20691));
  NANDX1 G26948 (.A1(W6305), .A2(W14774), .ZN(W20687));
  NANDX1 G26949 (.A1(W9030), .A2(W14463), .ZN(O2057));
  NANDX1 G26950 (.A1(W1527), .A2(I216), .ZN(W3172));
  NANDX1 G26951 (.A1(W3966), .A2(W875), .ZN(O2011));
  NANDX1 G26952 (.A1(W2355), .A2(W1123), .ZN(W3326));
  NANDX1 G26953 (.A1(W10128), .A2(I1621), .ZN(O601));
  NANDX1 G26954 (.A1(W13988), .A2(W8191), .ZN(W20459));
  NANDX1 G26955 (.A1(W9871), .A2(W15093), .ZN(O2013));
  NANDX1 G26956 (.A1(I354), .A2(W1677), .ZN(W3330));
  NANDX1 G26957 (.A1(W2083), .A2(I1149), .ZN(W3331));
  NANDX1 G26958 (.A1(W5300), .A2(W5292), .ZN(W8659));
  NANDX1 G26959 (.A1(W6496), .A2(W10132), .ZN(W12434));
  NANDX1 G26960 (.A1(W5353), .A2(W1418), .ZN(W20451));
  NANDX1 G26961 (.A1(W15801), .A2(W2486), .ZN(W20462));
  NANDX1 G26962 (.A1(W539), .A2(I1864), .ZN(W3337));
  NANDX1 G26963 (.A1(W2325), .A2(W4689), .ZN(W8657));
  NANDX1 G26964 (.A1(W2516), .A2(W1568), .ZN(W3341));
  NANDX1 G26965 (.A1(W6470), .A2(W7797), .ZN(W20442));
  NANDX1 G26966 (.A1(W485), .A2(W1011), .ZN(W3343));
  NANDX1 G26967 (.A1(W8212), .A2(W7964), .ZN(W8656));
  NANDX1 G26968 (.A1(W16160), .A2(W7272), .ZN(W20433));
  NANDX1 G26969 (.A1(W10147), .A2(W4581), .ZN(W20432));
  NANDX1 G26970 (.A1(I1423), .A2(W2494), .ZN(W3320));
  NANDX1 G26971 (.A1(W15689), .A2(W10782), .ZN(W20482));
  NANDX1 G26972 (.A1(W14248), .A2(W10332), .ZN(W20481));
  NANDX1 G26973 (.A1(I921), .A2(I1755), .ZN(W20480));
  NANDX1 G26974 (.A1(I1844), .A2(W9511), .ZN(W12427));
  NANDX1 G26975 (.A1(W7422), .A2(W7100), .ZN(W20474));
  NANDX1 G26976 (.A1(W18375), .A2(W4923), .ZN(W20472));
  NANDX1 G26977 (.A1(W82), .A2(W13824), .ZN(W20471));
  NANDX1 G26978 (.A1(W2998), .A2(W12357), .ZN(W20470));
  NANDX1 G26979 (.A1(W11903), .A2(W19985), .ZN(W20431));
  NANDX1 G26980 (.A1(W11367), .A2(W17222), .ZN(W20468));
  NANDX1 G26981 (.A1(W8476), .A2(I1983), .ZN(W20467));
  NANDX1 G26982 (.A1(W970), .A2(W2034), .ZN(W3321));
  NANDX1 G26983 (.A1(W868), .A2(I500), .ZN(W3322));
  NANDX1 G26984 (.A1(W13353), .A2(W10937), .ZN(W20465));
  NANDX1 G26985 (.A1(W130), .A2(W1435), .ZN(W3324));
  NANDX1 G26986 (.A1(W19601), .A2(W20305), .ZN(W20464));
  NANDX1 G26987 (.A1(W958), .A2(W2751), .ZN(W3325));
  NANDX1 G26988 (.A1(W2116), .A2(W2364), .ZN(W3370));
  NANDX1 G26989 (.A1(W18827), .A2(W673), .ZN(O2003));
  NANDX1 G26990 (.A1(W248), .A2(W1786), .ZN(W3361));
  NANDX1 G26991 (.A1(I422), .A2(W3299), .ZN(W3362));
  NANDX1 G26992 (.A1(W7706), .A2(W3600), .ZN(O2001));
  NANDX1 G26993 (.A1(W5632), .A2(W1262), .ZN(W20403));
  NANDX1 G26994 (.A1(W346), .A2(I1027), .ZN(W3363));
  NANDX1 G26995 (.A1(W123), .A2(I976), .ZN(W12451));
  NANDX1 G26996 (.A1(W681), .A2(W817), .ZN(W3369));
  NANDX1 G26997 (.A1(W1662), .A2(W5670), .ZN(W8639));
  NANDX1 G26998 (.A1(W7830), .A2(W6147), .ZN(W20398));
  NANDX1 G26999 (.A1(W8581), .A2(W14991), .ZN(W20395));
  NANDX1 G27000 (.A1(W421), .A2(W254), .ZN(W3371));
  NANDX1 G27001 (.A1(W9212), .A2(W11568), .ZN(O1998));
  NANDX1 G27002 (.A1(W2034), .A2(W4054), .ZN(W8635));
  NANDX1 G27003 (.A1(W19845), .A2(W17072), .ZN(O1997));
  NANDX1 G27004 (.A1(I1716), .A2(I1602), .ZN(W20389));
  NANDX1 G27005 (.A1(W5997), .A2(W2071), .ZN(W8633));
  NANDX1 G27006 (.A1(W8189), .A2(W2965), .ZN(W8647));
  NANDX1 G27007 (.A1(W10610), .A2(W11742), .ZN(W20429));
  NANDX1 G27008 (.A1(W11216), .A2(W4077), .ZN(W20428));
  NANDX1 G27009 (.A1(W1409), .A2(W2531), .ZN(W3345));
  NANDX1 G27010 (.A1(W5461), .A2(I1886), .ZN(W8650));
  NANDX1 G27011 (.A1(W11566), .A2(W186), .ZN(W12437));
  NANDX1 G27012 (.A1(W3126), .A2(W7595), .ZN(W8649));
  NANDX1 G27013 (.A1(W7467), .A2(W2412), .ZN(W8648));
  NANDX1 G27014 (.A1(W3278), .A2(W10179), .ZN(W12441));
  NANDX1 G27015 (.A1(W11087), .A2(W18708), .ZN(W20483));
  NANDX1 G27016 (.A1(W52), .A2(W20114), .ZN(W20416));
  NANDX1 G27017 (.A1(W1260), .A2(W1004), .ZN(W3355));
  NANDX1 G27018 (.A1(W16682), .A2(W8417), .ZN(W20415));
  NANDX1 G27019 (.A1(W8448), .A2(W8328), .ZN(W8646));
  NANDX1 G27020 (.A1(I224), .A2(W5532), .ZN(W12447));
  NANDX1 G27021 (.A1(W1611), .A2(W6969), .ZN(W8643));
  NANDX1 G27022 (.A1(W16043), .A2(I918), .ZN(W20409));
  NANDX1 G27023 (.A1(W2672), .A2(I774), .ZN(W8641));
  NANDX1 G27024 (.A1(W653), .A2(W3682), .ZN(W8684));
  NANDX1 G27025 (.A1(W2829), .A2(I915), .ZN(W8694));
  NANDX1 G27026 (.A1(W15607), .A2(W6806), .ZN(W20541));
  NANDX1 G27027 (.A1(W20495), .A2(W2371), .ZN(W20540));
  NANDX1 G27028 (.A1(W825), .A2(W2983), .ZN(W3269));
  NANDX1 G27029 (.A1(W165), .A2(I1619), .ZN(W3272));
  NANDX1 G27030 (.A1(W1800), .A2(I1153), .ZN(W3273));
  NANDX1 G27031 (.A1(I1553), .A2(W299), .ZN(W3275));
  NANDX1 G27032 (.A1(W11666), .A2(W12657), .ZN(O2024));
  NANDX1 G27033 (.A1(W2794), .A2(W11831), .ZN(W12396));
  NANDX1 G27034 (.A1(W3098), .A2(I1768), .ZN(W3264));
  NANDX1 G27035 (.A1(W4101), .A2(W13593), .ZN(W20532));
  NANDX1 G27036 (.A1(I1935), .A2(W5700), .ZN(W20529));
  NANDX1 G27037 (.A1(W9818), .A2(I836), .ZN(W20528));
  NANDX1 G27038 (.A1(W1730), .A2(W752), .ZN(W3280));
  NANDX1 G27039 (.A1(W2387), .A2(W15366), .ZN(W20525));
  NANDX1 G27040 (.A1(W12297), .A2(W4147), .ZN(W12399));
  NANDX1 G27041 (.A1(W18799), .A2(I1152), .ZN(W20518));
  NANDX1 G27042 (.A1(W3169), .A2(W9488), .ZN(W12401));
  NANDX1 G27043 (.A1(I1596), .A2(W2946), .ZN(W3258));
  NANDX1 G27044 (.A1(W2182), .A2(I1568), .ZN(W3253));
  NANDX1 G27045 (.A1(W17921), .A2(W7401), .ZN(W20564));
  NANDX1 G27046 (.A1(W11590), .A2(W4185), .ZN(W20561));
  NANDX1 G27047 (.A1(W4025), .A2(W1463), .ZN(W20560));
  NANDX1 G27048 (.A1(W8566), .A2(W14301), .ZN(O2031));
  NANDX1 G27049 (.A1(I1815), .A2(I1398), .ZN(W3254));
  NANDX1 G27050 (.A1(W2992), .A2(I716), .ZN(W12387));
  NANDX1 G27051 (.A1(W854), .A2(I1330), .ZN(W3255));
  NANDX1 G27052 (.A1(W1285), .A2(W1835), .ZN(W3281));
  NANDX1 G27053 (.A1(W11538), .A2(W20331), .ZN(W20553));
  NANDX1 G27054 (.A1(W14862), .A2(W564), .ZN(W20551));
  NANDX1 G27055 (.A1(W4238), .A2(W7982), .ZN(W12388));
  NANDX1 G27056 (.A1(W9264), .A2(W6317), .ZN(W12389));
  NANDX1 G27057 (.A1(W3025), .A2(I965), .ZN(W3260));
  NANDX1 G27058 (.A1(W6798), .A2(I451), .ZN(W20545));
  NANDX1 G27059 (.A1(W2683), .A2(W270), .ZN(W3262));
  NANDX1 G27060 (.A1(W7204), .A2(W2855), .ZN(W8695));
  NANDX1 G27061 (.A1(W2082), .A2(W15786), .ZN(W20490));
  NANDX1 G27062 (.A1(I696), .A2(W14468), .ZN(W20498));
  NANDX1 G27063 (.A1(W4834), .A2(W5024), .ZN(W20497));
  NANDX1 G27064 (.A1(W2112), .A2(I1225), .ZN(W3298));
  NANDX1 G27065 (.A1(I1421), .A2(W4622), .ZN(W8673));
  NANDX1 G27066 (.A1(W7887), .A2(W16391), .ZN(W20493));
  NANDX1 G27067 (.A1(W418), .A2(W7653), .ZN(O600));
  NANDX1 G27068 (.A1(W3210), .A2(I652), .ZN(W3305));
  NANDX1 G27069 (.A1(W15195), .A2(W6726), .ZN(O2017));
  NANDX1 G27070 (.A1(I349), .A2(W15597), .ZN(W20499));
  NANDX1 G27071 (.A1(W4826), .A2(W6534), .ZN(W8671));
  NANDX1 G27072 (.A1(I1894), .A2(W905), .ZN(W3309));
  NANDX1 G27073 (.A1(W8783), .A2(W367), .ZN(W20486));
  NANDX1 G27074 (.A1(W9440), .A2(W10500), .ZN(W12424));
  NANDX1 G27075 (.A1(I911), .A2(W2706), .ZN(W3312));
  NANDX1 G27076 (.A1(W639), .A2(I1813), .ZN(W3313));
  NANDX1 G27077 (.A1(W3049), .A2(W7083), .ZN(W8667));
  NANDX1 G27078 (.A1(W5092), .A2(W2332), .ZN(W8666));
  NANDX1 G27079 (.A1(W16929), .A2(I442), .ZN(O2020));
  NANDX1 G27080 (.A1(W7330), .A2(W7068), .ZN(W12404));
  NANDX1 G27081 (.A1(W17379), .A2(W11223), .ZN(W20514));
  NANDX1 G27082 (.A1(W16413), .A2(W4255), .ZN(W20513));
  NANDX1 G27083 (.A1(W11875), .A2(W1838), .ZN(W20512));
  NANDX1 G27084 (.A1(W5125), .A2(I576), .ZN(W8680));
  NANDX1 G27085 (.A1(W232), .A2(W11764), .ZN(W12405));
  NANDX1 G27086 (.A1(W2743), .A2(W120), .ZN(W3286));
  NANDX1 G27087 (.A1(W4883), .A2(W3196), .ZN(W12406));
  NANDX1 G27088 (.A1(W2569), .A2(W2673), .ZN(W8517));
  NANDX1 G27089 (.A1(W1675), .A2(W6531), .ZN(W8679));
  NANDX1 G27090 (.A1(W13134), .A2(W8287), .ZN(W20507));
  NANDX1 G27091 (.A1(W8302), .A2(W6072), .ZN(W8677));
  NANDX1 G27092 (.A1(W7604), .A2(W13389), .ZN(W20506));
  NANDX1 G27093 (.A1(W1690), .A2(W2734), .ZN(W12412));
  NANDX1 G27094 (.A1(W2439), .A2(W1117), .ZN(W3294));
  NANDX1 G27095 (.A1(W19096), .A2(W13129), .ZN(W20503));
  NANDX1 G27096 (.A1(I249), .A2(W13329), .ZN(O2018));
  NANDX1 G27097 (.A1(I288), .A2(W11338), .ZN(W19572));
  NANDX1 G27098 (.A1(W3036), .A2(W2089), .ZN(W3974));
  NANDX1 G27099 (.A1(I1108), .A2(W845), .ZN(W3975));
  NANDX1 G27100 (.A1(W2030), .A2(I1593), .ZN(W3976));
  NANDX1 G27101 (.A1(W4759), .A2(W1601), .ZN(W8374));
  NANDX1 G27102 (.A1(W17982), .A2(W1275), .ZN(W19580));
  NANDX1 G27103 (.A1(I151), .A2(W1174), .ZN(W8373));
  NANDX1 G27104 (.A1(I670), .A2(W1649), .ZN(W3978));
  NANDX1 G27105 (.A1(W1466), .A2(W2787), .ZN(W3979));
  NANDX1 G27106 (.A1(W8875), .A2(W4327), .ZN(W12860));
  NANDX1 G27107 (.A1(W6312), .A2(W5784), .ZN(W8376));
  NANDX1 G27108 (.A1(W4651), .A2(W3401), .ZN(W12862));
  NANDX1 G27109 (.A1(W19290), .A2(W14895), .ZN(W19567));
  NANDX1 G27110 (.A1(W10743), .A2(W8013), .ZN(W12863));
  NANDX1 G27111 (.A1(W4432), .A2(I460), .ZN(W8370));
  NANDX1 G27112 (.A1(W3165), .A2(W2229), .ZN(W3984));
  NANDX1 G27113 (.A1(W12553), .A2(W12430), .ZN(W19562));
  NANDX1 G27114 (.A1(W3320), .A2(W4076), .ZN(W12867));
  NANDX1 G27115 (.A1(W15165), .A2(W15438), .ZN(O1797));
  NANDX1 G27116 (.A1(W7873), .A2(I670), .ZN(O1805));
  NANDX1 G27117 (.A1(W11587), .A2(W3300), .ZN(O1807));
  NANDX1 G27118 (.A1(W1360), .A2(W9450), .ZN(W12845));
  NANDX1 G27119 (.A1(W5052), .A2(W1237), .ZN(W8382));
  NANDX1 G27120 (.A1(W2355), .A2(I1136), .ZN(W3962));
  NANDX1 G27121 (.A1(I817), .A2(W8937), .ZN(W12851));
  NANDX1 G27122 (.A1(W683), .A2(W665), .ZN(W3964));
  NANDX1 G27123 (.A1(I179), .A2(W1067), .ZN(W19595));
  NANDX1 G27124 (.A1(W3775), .A2(W8642), .ZN(W19593));
  NANDX1 G27125 (.A1(W10347), .A2(W15717), .ZN(W19555));
  NANDX1 G27126 (.A1(I254), .A2(W4611), .ZN(W8380));
  NANDX1 G27127 (.A1(W12761), .A2(W18109), .ZN(W19591));
  NANDX1 G27128 (.A1(W1898), .A2(I389), .ZN(W8377));
  NANDX1 G27129 (.A1(W13260), .A2(W17946), .ZN(W19590));
  NANDX1 G27130 (.A1(W13034), .A2(I1266), .ZN(O1804));
  NANDX1 G27131 (.A1(W17858), .A2(W8678), .ZN(W19588));
  NANDX1 G27132 (.A1(W9868), .A2(W4382), .ZN(W12854));
  NANDX1 G27133 (.A1(W2450), .A2(W3309), .ZN(W3972));
  NANDX1 G27134 (.A1(I552), .A2(W3661), .ZN(W4007));
  NANDX1 G27135 (.A1(W3318), .A2(W1316), .ZN(W19530));
  NANDX1 G27136 (.A1(I1180), .A2(W1397), .ZN(W8360));
  NANDX1 G27137 (.A1(W3023), .A2(W3043), .ZN(W19527));
  NANDX1 G27138 (.A1(I1337), .A2(W2771), .ZN(W8359));
  NANDX1 G27139 (.A1(I1090), .A2(W3581), .ZN(W19525));
  NANDX1 G27140 (.A1(W7846), .A2(W5156), .ZN(W12891));
  NANDX1 G27141 (.A1(W16753), .A2(W4629), .ZN(W19523));
  NANDX1 G27142 (.A1(W7548), .A2(W4827), .ZN(W12892));
  NANDX1 G27143 (.A1(W9771), .A2(W10207), .ZN(W12884));
  NANDX1 G27144 (.A1(W17246), .A2(W15156), .ZN(W19520));
  NANDX1 G27145 (.A1(W256), .A2(W6026), .ZN(W12894));
  NANDX1 G27146 (.A1(W7442), .A2(W8113), .ZN(W12896));
  NANDX1 G27147 (.A1(W4177), .A2(W7872), .ZN(W8352));
  NANDX1 G27148 (.A1(I871), .A2(W2936), .ZN(W4012));
  NANDX1 G27149 (.A1(W16894), .A2(W15657), .ZN(O1788));
  NANDX1 G27150 (.A1(W1440), .A2(W2197), .ZN(W4013));
  NANDX1 G27151 (.A1(I576), .A2(W2113), .ZN(W8349));
  NANDX1 G27152 (.A1(W17227), .A2(W7773), .ZN(O1793));
  NANDX1 G27153 (.A1(W16376), .A2(W8551), .ZN(O1796));
  NANDX1 G27154 (.A1(W6196), .A2(W15500), .ZN(O1795));
  NANDX1 G27155 (.A1(W3201), .A2(W11641), .ZN(W12873));
  NANDX1 G27156 (.A1(W11574), .A2(W816), .ZN(W12876));
  NANDX1 G27157 (.A1(I1892), .A2(W7201), .ZN(W12877));
  NANDX1 G27158 (.A1(W2596), .A2(W3645), .ZN(W3995));
  NANDX1 G27159 (.A1(W12372), .A2(W10691), .ZN(W19547));
  NANDX1 G27160 (.A1(W9830), .A2(W3187), .ZN(W12878));
  NANDX1 G27161 (.A1(I220), .A2(I1883), .ZN(W8389));
  NANDX1 G27162 (.A1(W9684), .A2(W1094), .ZN(O1792));
  NANDX1 G27163 (.A1(W82), .A2(W13730), .ZN(O1791));
  NANDX1 G27164 (.A1(W6471), .A2(W8189), .ZN(W8366));
  NANDX1 G27165 (.A1(W2655), .A2(W5054), .ZN(W8365));
  NANDX1 G27166 (.A1(W5197), .A2(W15472), .ZN(W19539));
  NANDX1 G27167 (.A1(W4551), .A2(W6740), .ZN(W12879));
  NANDX1 G27168 (.A1(W5238), .A2(I448), .ZN(W8364));
  NANDX1 G27169 (.A1(W8552), .A2(W7888), .ZN(W12882));
  NANDX1 G27170 (.A1(W1638), .A2(W1283), .ZN(W3906));
  NANDX1 G27171 (.A1(W19244), .A2(W11430), .ZN(W19678));
  NANDX1 G27172 (.A1(I198), .A2(W2347), .ZN(O48));
  NANDX1 G27173 (.A1(W654), .A2(I1939), .ZN(W3902));
  NANDX1 G27174 (.A1(W1596), .A2(I913), .ZN(W3903));
  NANDX1 G27175 (.A1(I1848), .A2(W460), .ZN(W3904));
  NANDX1 G27176 (.A1(W8845), .A2(I1293), .ZN(O1821));
  NANDX1 G27177 (.A1(W9827), .A2(W7918), .ZN(W19671));
  NANDX1 G27178 (.A1(W629), .A2(W5484), .ZN(O655));
  NANDX1 G27179 (.A1(W9913), .A2(W1085), .ZN(W19667));
  NANDX1 G27180 (.A1(W1565), .A2(W2073), .ZN(W8400));
  NANDX1 G27181 (.A1(W11), .A2(W7970), .ZN(W19666));
  NANDX1 G27182 (.A1(W19180), .A2(W11654), .ZN(W19664));
  NANDX1 G27183 (.A1(I720), .A2(W2293), .ZN(W3909));
  NANDX1 G27184 (.A1(W6794), .A2(I1801), .ZN(W8395));
  NANDX1 G27185 (.A1(W924), .A2(W323), .ZN(W3911));
  NANDX1 G27186 (.A1(W3091), .A2(W3906), .ZN(W12818));
  NANDX1 G27187 (.A1(W311), .A2(W10703), .ZN(W12819));
  NANDX1 G27188 (.A1(I1271), .A2(W11505), .ZN(W12821));
  NANDX1 G27189 (.A1(W12090), .A2(W19561), .ZN(O1823));
  NANDX1 G27190 (.A1(W16854), .A2(I1762), .ZN(W19700));
  NANDX1 G27191 (.A1(I371), .A2(W18960), .ZN(W19698));
  NANDX1 G27192 (.A1(W4104), .A2(W4474), .ZN(W12797));
  NANDX1 G27193 (.A1(W1812), .A2(I1480), .ZN(W8410));
  NANDX1 G27194 (.A1(W6182), .A2(I1096), .ZN(W12799));
  NANDX1 G27195 (.A1(W7185), .A2(W2787), .ZN(O652));
  NANDX1 G27196 (.A1(W5738), .A2(W5990), .ZN(W8408));
  NANDX1 G27197 (.A1(I463), .A2(W3875), .ZN(W3894));
  NANDX1 G27198 (.A1(W8664), .A2(I1098), .ZN(W19649));
  NANDX1 G27199 (.A1(W1833), .A2(W3405), .ZN(W3897));
  NANDX1 G27200 (.A1(W1620), .A2(W4846), .ZN(W8404));
  NANDX1 G27201 (.A1(W7321), .A2(W6988), .ZN(W19683));
  NANDX1 G27202 (.A1(W11639), .A2(W3074), .ZN(W19682));
  NANDX1 G27203 (.A1(W7577), .A2(W3181), .ZN(W8401));
  NANDX1 G27204 (.A1(W4265), .A2(W15136), .ZN(W19681));
  NANDX1 G27205 (.A1(W10456), .A2(W10049), .ZN(W19680));
  NANDX1 G27206 (.A1(W4525), .A2(W1570), .ZN(W12810));
  NANDX1 G27207 (.A1(W9556), .A2(I1930), .ZN(W12836));
  NANDX1 G27208 (.A1(W3617), .A2(W693), .ZN(W3941));
  NANDX1 G27209 (.A1(W4210), .A2(W1252), .ZN(W19623));
  NANDX1 G27210 (.A1(W11467), .A2(W3216), .ZN(O1809));
  NANDX1 G27211 (.A1(W1838), .A2(W2737), .ZN(W3942));
  NANDX1 G27212 (.A1(W969), .A2(I488), .ZN(W3943));
  NANDX1 G27213 (.A1(W7402), .A2(W6930), .ZN(W8391));
  NANDX1 G27214 (.A1(W960), .A2(I983), .ZN(W3947));
  NANDX1 G27215 (.A1(W15391), .A2(W18712), .ZN(W19613));
  NANDX1 G27216 (.A1(I1722), .A2(W4933), .ZN(W19628));
  NANDX1 G27217 (.A1(W248), .A2(W255), .ZN(W3950));
  NANDX1 G27218 (.A1(W9834), .A2(W536), .ZN(W19612));
  NANDX1 G27219 (.A1(W3935), .A2(W1545), .ZN(W3952));
  NANDX1 G27220 (.A1(W2875), .A2(I1866), .ZN(W3953));
  NANDX1 G27221 (.A1(W2038), .A2(I640), .ZN(O49));
  NANDX1 G27222 (.A1(W69), .A2(W110), .ZN(W3956));
  NANDX1 G27223 (.A1(W12118), .A2(W2143), .ZN(W19609));
  NANDX1 G27224 (.A1(W12566), .A2(W13853), .ZN(W19608));
  NANDX1 G27225 (.A1(W1715), .A2(W462), .ZN(W3923));
  NANDX1 G27226 (.A1(W8399), .A2(I718), .ZN(W19648));
  NANDX1 G27227 (.A1(W8703), .A2(W11485), .ZN(W19646));
  NANDX1 G27228 (.A1(I798), .A2(I1107), .ZN(W3915));
  NANDX1 G27229 (.A1(I562), .A2(W881), .ZN(W3916));
  NANDX1 G27230 (.A1(W10381), .A2(W10247), .ZN(W12823));
  NANDX1 G27231 (.A1(W3057), .A2(W1528), .ZN(W3921));
  NANDX1 G27232 (.A1(W16507), .A2(W11500), .ZN(O1814));
  NANDX1 G27233 (.A1(W5086), .A2(W6881), .ZN(O226));
  NANDX1 G27234 (.A1(W14410), .A2(I491), .ZN(W19511));
  NANDX1 G27235 (.A1(W7808), .A2(W3149), .ZN(W19631));
  NANDX1 G27236 (.A1(I1590), .A2(I1305), .ZN(W3929));
  NANDX1 G27237 (.A1(W4623), .A2(I1514), .ZN(W12826));
  NANDX1 G27238 (.A1(W7097), .A2(W10919), .ZN(O657));
  NANDX1 G27239 (.A1(W1048), .A2(W11364), .ZN(W12829));
  NANDX1 G27240 (.A1(W2067), .A2(W5036), .ZN(W12831));
  NANDX1 G27241 (.A1(W2802), .A2(I234), .ZN(W3938));
  NANDX1 G27242 (.A1(W7205), .A2(W911), .ZN(W19629));
  NANDX1 G27243 (.A1(W458), .A2(W5131), .ZN(O667));
  NANDX1 G27244 (.A1(W14344), .A2(W1537), .ZN(W19397));
  NANDX1 G27245 (.A1(I1015), .A2(I1490), .ZN(W8314));
  NANDX1 G27246 (.A1(I192), .A2(W612), .ZN(W4098));
  NANDX1 G27247 (.A1(W3342), .A2(W3885), .ZN(W4100));
  NANDX1 G27248 (.A1(W221), .A2(W400), .ZN(W4101));
  NANDX1 G27249 (.A1(W13963), .A2(W11885), .ZN(W19391));
  NANDX1 G27250 (.A1(W5568), .A2(W5770), .ZN(W12936));
  NANDX1 G27251 (.A1(I1932), .A2(W2367), .ZN(W4104));
  NANDX1 G27252 (.A1(I723), .A2(I1504), .ZN(W4105));
  NANDX1 G27253 (.A1(W3519), .A2(W3435), .ZN(W4095));
  NANDX1 G27254 (.A1(W6455), .A2(I1610), .ZN(W8310));
  NANDX1 G27255 (.A1(I636), .A2(W4122), .ZN(W8308));
  NANDX1 G27256 (.A1(W2131), .A2(W7632), .ZN(W8307));
  NANDX1 G27257 (.A1(W14244), .A2(W12473), .ZN(W19377));
  NANDX1 G27258 (.A1(W2594), .A2(W598), .ZN(W4111));
  NANDX1 G27259 (.A1(W12702), .A2(I1450), .ZN(O669));
  NANDX1 G27260 (.A1(I1367), .A2(W11396), .ZN(W19374));
  NANDX1 G27261 (.A1(W4513), .A2(W3132), .ZN(W8305));
  NANDX1 G27262 (.A1(W5590), .A2(W487), .ZN(W12929));
  NANDX1 G27263 (.A1(I1762), .A2(I318), .ZN(W4078));
  NANDX1 G27264 (.A1(W8785), .A2(W4184), .ZN(W12922));
  NANDX1 G27265 (.A1(I877), .A2(W5080), .ZN(W12925));
  NANDX1 G27266 (.A1(W8228), .A2(W6374), .ZN(W19415));
  NANDX1 G27267 (.A1(W19120), .A2(W8830), .ZN(W19414));
  NANDX1 G27268 (.A1(W6768), .A2(W5453), .ZN(W8322));
  NANDX1 G27269 (.A1(W8039), .A2(W5058), .ZN(W8320));
  NANDX1 G27270 (.A1(W18986), .A2(W12871), .ZN(W19413));
  NANDX1 G27271 (.A1(W6822), .A2(I1991), .ZN(O1757));
  NANDX1 G27272 (.A1(W8586), .A2(I1463), .ZN(W12930));
  NANDX1 G27273 (.A1(W2727), .A2(W1344), .ZN(W4084));
  NANDX1 G27274 (.A1(W3863), .A2(W13008), .ZN(W19407));
  NANDX1 G27275 (.A1(W2444), .A2(I672), .ZN(W8318));
  NANDX1 G27276 (.A1(W3482), .A2(W579), .ZN(W4090));
  NANDX1 G27277 (.A1(W9554), .A2(W2823), .ZN(W19403));
  NANDX1 G27278 (.A1(W13346), .A2(W7741), .ZN(O1765));
  NANDX1 G27279 (.A1(W11447), .A2(W2037), .ZN(W19399));
  NANDX1 G27280 (.A1(W5990), .A2(W5919), .ZN(W8295));
  NANDX1 G27281 (.A1(W878), .A2(W1540), .ZN(W4130));
  NANDX1 G27282 (.A1(W196), .A2(I1004), .ZN(O1750));
  NANDX1 G27283 (.A1(W3256), .A2(W1815), .ZN(W4133));
  NANDX1 G27284 (.A1(W473), .A2(I1273), .ZN(W19331));
  NANDX1 G27285 (.A1(I1651), .A2(W967), .ZN(W4134));
  NANDX1 G27286 (.A1(W10231), .A2(W3), .ZN(W19330));
  NANDX1 G27287 (.A1(I1535), .A2(W2482), .ZN(W4135));
  NANDX1 G27288 (.A1(W700), .A2(W2015), .ZN(W4138));
  NANDX1 G27289 (.A1(W668), .A2(W3891), .ZN(W4127));
  NANDX1 G27290 (.A1(W19067), .A2(W12857), .ZN(O1749));
  NANDX1 G27291 (.A1(I1883), .A2(W7703), .ZN(W8294));
  NANDX1 G27292 (.A1(W1667), .A2(W3426), .ZN(W4140));
  NANDX1 G27293 (.A1(W12299), .A2(W13073), .ZN(O1748));
  NANDX1 G27294 (.A1(W5102), .A2(W11692), .ZN(W19323));
  NANDX1 G27295 (.A1(W7345), .A2(I30), .ZN(W8293));
  NANDX1 G27296 (.A1(W2391), .A2(I973), .ZN(W4145));
  NANDX1 G27297 (.A1(W3097), .A2(W2620), .ZN(O674));
  NANDX1 G27298 (.A1(W4881), .A2(I637), .ZN(W19356));
  NANDX1 G27299 (.A1(W6053), .A2(W1465), .ZN(W19367));
  NANDX1 G27300 (.A1(W7013), .A2(I206), .ZN(O1755));
  NANDX1 G27301 (.A1(W13830), .A2(W15693), .ZN(O1754));
  NANDX1 G27302 (.A1(W5191), .A2(W10691), .ZN(W19364));
  NANDX1 G27303 (.A1(W3466), .A2(W5136), .ZN(O671));
  NANDX1 G27304 (.A1(W1412), .A2(W749), .ZN(W8304));
  NANDX1 G27305 (.A1(W18713), .A2(W8670), .ZN(W19358));
  NANDX1 G27306 (.A1(W3880), .A2(W4826), .ZN(W8301));
  NANDX1 G27307 (.A1(I146), .A2(W865), .ZN(W8327));
  NANDX1 G27308 (.A1(I1503), .A2(W7965), .ZN(W12952));
  NANDX1 G27309 (.A1(W7510), .A2(W8077), .ZN(W12962));
  NANDX1 G27310 (.A1(W2173), .A2(W6983), .ZN(W19351));
  NANDX1 G27311 (.A1(W2166), .A2(W3359), .ZN(W4119));
  NANDX1 G27312 (.A1(W5510), .A2(W1375), .ZN(W19343));
  NANDX1 G27313 (.A1(W2522), .A2(W7602), .ZN(W8300));
  NANDX1 G27314 (.A1(I557), .A2(W1126), .ZN(W4120));
  NANDX1 G27315 (.A1(W5082), .A2(W6518), .ZN(W12968));
  NANDX1 G27316 (.A1(W16857), .A2(W4709), .ZN(W19476));
  NANDX1 G27317 (.A1(W2299), .A2(W14406), .ZN(W19485));
  NANDX1 G27318 (.A1(I820), .A2(W3677), .ZN(W4029));
  NANDX1 G27319 (.A1(W12214), .A2(W2040), .ZN(W12903));
  NANDX1 G27320 (.A1(W3708), .A2(W331), .ZN(W4032));
  NANDX1 G27321 (.A1(W3913), .A2(W3175), .ZN(W4033));
  NANDX1 G27322 (.A1(W513), .A2(W3159), .ZN(W4036));
  NANDX1 G27323 (.A1(I665), .A2(W7319), .ZN(W12904));
  NANDX1 G27324 (.A1(W3627), .A2(W2016), .ZN(W4037));
  NANDX1 G27325 (.A1(W10727), .A2(W17810), .ZN(W19477));
  NANDX1 G27326 (.A1(W2307), .A2(W2951), .ZN(W4028));
  NANDX1 G27327 (.A1(W14591), .A2(W7576), .ZN(W19474));
  NANDX1 G27328 (.A1(I674), .A2(W244), .ZN(W4038));
  NANDX1 G27329 (.A1(W435), .A2(W17022), .ZN(W19473));
  NANDX1 G27330 (.A1(W8855), .A2(W17893), .ZN(O1779));
  NANDX1 G27331 (.A1(W1059), .A2(I1841), .ZN(O222));
  NANDX1 G27332 (.A1(W1717), .A2(W2198), .ZN(W8332));
  NANDX1 G27333 (.A1(W3303), .A2(W1033), .ZN(W4046));
  NANDX1 G27334 (.A1(W16603), .A2(W16173), .ZN(W19467));
  NANDX1 G27335 (.A1(I1021), .A2(W12729), .ZN(W19496));
  NANDX1 G27336 (.A1(W13088), .A2(W13210), .ZN(W19508));
  NANDX1 G27337 (.A1(I1720), .A2(W10997), .ZN(W12899));
  NANDX1 G27338 (.A1(W8541), .A2(W8610), .ZN(O1786));
  NANDX1 G27339 (.A1(I1119), .A2(W4044), .ZN(W8348));
  NANDX1 G27340 (.A1(W2426), .A2(I1907), .ZN(W4021));
  NANDX1 G27341 (.A1(W4123), .A2(W1523), .ZN(W8346));
  NANDX1 G27342 (.A1(W4428), .A2(I925), .ZN(W19502));
  NANDX1 G27343 (.A1(W11351), .A2(W1104), .ZN(W19501));
  NANDX1 G27344 (.A1(W145), .A2(W2342), .ZN(W4047));
  NANDX1 G27345 (.A1(W17402), .A2(W8999), .ZN(W19494));
  NANDX1 G27346 (.A1(I1073), .A2(I1090), .ZN(W4026));
  NANDX1 G27347 (.A1(W6625), .A2(W9252), .ZN(W12902));
  NANDX1 G27348 (.A1(W16322), .A2(W19420), .ZN(O1782));
  NANDX1 G27349 (.A1(W937), .A2(W294), .ZN(W8344));
  NANDX1 G27350 (.A1(W2336), .A2(W698), .ZN(W4027));
  NANDX1 G27351 (.A1(W6902), .A2(W17584), .ZN(W19488));
  NANDX1 G27352 (.A1(W18274), .A2(W18660), .ZN(W19487));
  NANDX1 G27353 (.A1(W10172), .A2(W3684), .ZN(W12916));
  NANDX1 G27354 (.A1(W1671), .A2(W3495), .ZN(W19437));
  NANDX1 G27355 (.A1(W1212), .A2(W1383), .ZN(W4062));
  NANDX1 G27356 (.A1(W5952), .A2(W10984), .ZN(W19433));
  NANDX1 G27357 (.A1(W2061), .A2(W771), .ZN(W4066));
  NANDX1 G27358 (.A1(W3644), .A2(W3599), .ZN(W4067));
  NANDX1 G27359 (.A1(I806), .A2(I509), .ZN(W4069));
  NANDX1 G27360 (.A1(W12075), .A2(W2838), .ZN(W19428));
  NANDX1 G27361 (.A1(W72), .A2(I662), .ZN(W4072));
  NANDX1 G27362 (.A1(W7884), .A2(W6966), .ZN(O1775));
  NANDX1 G27363 (.A1(W9299), .A2(W2304), .ZN(O664));
  NANDX1 G27364 (.A1(W4954), .A2(W8544), .ZN(O1771));
  NANDX1 G27365 (.A1(W3351), .A2(W10310), .ZN(W19421));
  NANDX1 G27366 (.A1(W3646), .A2(I1733), .ZN(W19420));
  NANDX1 G27367 (.A1(W17639), .A2(W18736), .ZN(W19419));
  NANDX1 G27368 (.A1(I20), .A2(W1318), .ZN(W4076));
  NANDX1 G27369 (.A1(W8145), .A2(W4398), .ZN(W8328));
  NANDX1 G27370 (.A1(W802), .A2(I1378), .ZN(W4077));
  NANDX1 G27371 (.A1(I1557), .A2(W9980), .ZN(W19456));
  NANDX1 G27372 (.A1(I1740), .A2(I1978), .ZN(W8331));
  NANDX1 G27373 (.A1(I1824), .A2(W1448), .ZN(W4050));
  NANDX1 G27374 (.A1(W5619), .A2(W12365), .ZN(W19460));
  NANDX1 G27375 (.A1(I673), .A2(W4729), .ZN(W19459));
  NANDX1 G27376 (.A1(W6680), .A2(W5855), .ZN(W12909));
  NANDX1 G27377 (.A1(W1381), .A2(W9889), .ZN(W19457));
  NANDX1 G27378 (.A1(W7605), .A2(W10411), .ZN(W12910));
  NANDX1 G27379 (.A1(W3891), .A2(W673), .ZN(W4054));
  NANDX1 G27380 (.A1(W8705), .A2(W8223), .ZN(W12795));
  NANDX1 G27381 (.A1(W2088), .A2(I310), .ZN(W4058));
  NANDX1 G27382 (.A1(W13780), .A2(W11220), .ZN(W19452));
  NANDX1 G27383 (.A1(W5658), .A2(I1920), .ZN(W19451));
  NANDX1 G27384 (.A1(I1340), .A2(W1088), .ZN(W12912));
  NANDX1 G27385 (.A1(W18618), .A2(W11635), .ZN(W19447));
  NANDX1 G27386 (.A1(W19022), .A2(W10435), .ZN(W19446));
  NANDX1 G27387 (.A1(W3206), .A2(W2751), .ZN(W4059));
  NANDX1 G27388 (.A1(W15992), .A2(I503), .ZN(W19441));
  NANDX1 G27389 (.A1(W7539), .A2(W2169), .ZN(W8466));
  NANDX1 G27390 (.A1(I924), .A2(W418), .ZN(W3718));
  NANDX1 G27391 (.A1(I1658), .A2(W59), .ZN(W19940));
  NANDX1 G27392 (.A1(I1259), .A2(W5958), .ZN(O1889));
  NANDX1 G27393 (.A1(W1366), .A2(W1705), .ZN(W3722));
  NANDX1 G27394 (.A1(W1343), .A2(W2765), .ZN(W3723));
  NANDX1 G27395 (.A1(W315), .A2(I1248), .ZN(W19934));
  NANDX1 G27396 (.A1(W5056), .A2(I193), .ZN(W19930));
  NANDX1 G27397 (.A1(W429), .A2(I65), .ZN(W8467));
  NANDX1 G27398 (.A1(W17191), .A2(W3069), .ZN(O1885));
  NANDX1 G27399 (.A1(W14333), .A2(I436), .ZN(W19942));
  NANDX1 G27400 (.A1(W7912), .A2(W18042), .ZN(W19923));
  NANDX1 G27401 (.A1(W6234), .A2(W8108), .ZN(W12682));
  NANDX1 G27402 (.A1(W16897), .A2(W18734), .ZN(W19922));
  NANDX1 G27403 (.A1(I1935), .A2(W762), .ZN(W3728));
  NANDX1 G27404 (.A1(W13011), .A2(W3454), .ZN(O1883));
  NANDX1 G27405 (.A1(W2496), .A2(W7956), .ZN(W12684));
  NANDX1 G27406 (.A1(W10652), .A2(W14110), .ZN(W19916));
  NANDX1 G27407 (.A1(W392), .A2(W19773), .ZN(W19915));
  NANDX1 G27408 (.A1(W8298), .A2(W5040), .ZN(W19954));
  NANDX1 G27409 (.A1(W16469), .A2(W668), .ZN(W19966));
  NANDX1 G27410 (.A1(W6592), .A2(W3982), .ZN(W19964));
  NANDX1 G27411 (.A1(W12228), .A2(W17736), .ZN(W19962));
  NANDX1 G27412 (.A1(W2502), .A2(W5505), .ZN(W8484));
  NANDX1 G27413 (.A1(W7968), .A2(W2759), .ZN(O1896));
  NANDX1 G27414 (.A1(I844), .A2(W127), .ZN(W3703));
  NANDX1 G27415 (.A1(W7599), .A2(W5167), .ZN(W8482));
  NANDX1 G27416 (.A1(W1585), .A2(W7216), .ZN(W19956));
  NANDX1 G27417 (.A1(I1610), .A2(W6122), .ZN(O231));
  NANDX1 G27418 (.A1(W2442), .A2(W9139), .ZN(W12676));
  NANDX1 G27419 (.A1(W2829), .A2(W2794), .ZN(W19949));
  NANDX1 G27420 (.A1(W2768), .A2(W3350), .ZN(W3711));
  NANDX1 G27421 (.A1(W731), .A2(I157), .ZN(W19948));
  NANDX1 G27422 (.A1(W16043), .A2(W2318), .ZN(O1893));
  NANDX1 G27423 (.A1(W9247), .A2(I1870), .ZN(W19946));
  NANDX1 G27424 (.A1(W1600), .A2(I1883), .ZN(W3714));
  NANDX1 G27425 (.A1(W15377), .A2(I583), .ZN(W19944));
  NANDX1 G27426 (.A1(I1477), .A2(W7098), .ZN(W19889));
  NANDX1 G27427 (.A1(W12736), .A2(W19245), .ZN(W19897));
  NANDX1 G27428 (.A1(I1920), .A2(I753), .ZN(O42));
  NANDX1 G27429 (.A1(I220), .A2(W1494), .ZN(O43));
  NANDX1 G27430 (.A1(W3384), .A2(W1063), .ZN(W8457));
  NANDX1 G27431 (.A1(W2608), .A2(W17023), .ZN(W19895));
  NANDX1 G27432 (.A1(W1219), .A2(W4912), .ZN(W12689));
  NANDX1 G27433 (.A1(W2812), .A2(I1314), .ZN(W3753));
  NANDX1 G27434 (.A1(W1772), .A2(W15626), .ZN(W19890));
  NANDX1 G27435 (.A1(W133), .A2(I1422), .ZN(W3747));
  NANDX1 G27436 (.A1(W2248), .A2(W12456), .ZN(W12691));
  NANDX1 G27437 (.A1(W11960), .A2(W4302), .ZN(W12693));
  NANDX1 G27438 (.A1(W3693), .A2(W3451), .ZN(W3755));
  NANDX1 G27439 (.A1(W5120), .A2(W15652), .ZN(O1877));
  NANDX1 G27440 (.A1(W10161), .A2(W7592), .ZN(O635));
  NANDX1 G27441 (.A1(W6952), .A2(W16666), .ZN(W19880));
  NANDX1 G27442 (.A1(W14057), .A2(I1666), .ZN(O1876));
  NANDX1 G27443 (.A1(W991), .A2(W516), .ZN(W19876));
  NANDX1 G27444 (.A1(W5510), .A2(W12745), .ZN(W19908));
  NANDX1 G27445 (.A1(W2500), .A2(W2297), .ZN(W3734));
  NANDX1 G27446 (.A1(W1341), .A2(W8203), .ZN(W12685));
  NANDX1 G27447 (.A1(W2809), .A2(I50), .ZN(W3735));
  NANDX1 G27448 (.A1(W673), .A2(W8791), .ZN(O1882));
  NANDX1 G27449 (.A1(W1740), .A2(W4400), .ZN(O1881));
  NANDX1 G27450 (.A1(W1249), .A2(W764), .ZN(W3737));
  NANDX1 G27451 (.A1(W17061), .A2(W10677), .ZN(W19909));
  NANDX1 G27452 (.A1(I875), .A2(I1224), .ZN(W3738));
  NANDX1 G27453 (.A1(W9045), .A2(W11555), .ZN(W19967));
  NANDX1 G27454 (.A1(W889), .A2(I1957), .ZN(W3739));
  NANDX1 G27455 (.A1(I1877), .A2(I1714), .ZN(W12686));
  NANDX1 G27456 (.A1(W978), .A2(W871), .ZN(O41));
  NANDX1 G27457 (.A1(W8300), .A2(W6602), .ZN(W8460));
  NANDX1 G27458 (.A1(I833), .A2(W3498), .ZN(W3746));
  NANDX1 G27459 (.A1(W4739), .A2(W6401), .ZN(W8458));
  NANDX1 G27460 (.A1(W192), .A2(W1235), .ZN(W19903));
  NANDX1 G27461 (.A1(W10152), .A2(W3491), .ZN(W19902));
  NANDX1 G27462 (.A1(W11986), .A2(I519), .ZN(W12639));
  NANDX1 G27463 (.A1(I1596), .A2(W17885), .ZN(W20023));
  NANDX1 G27464 (.A1(W9048), .A2(W3155), .ZN(W20022));
  NANDX1 G27465 (.A1(W15687), .A2(W11082), .ZN(W20020));
  NANDX1 G27466 (.A1(W937), .A2(W584), .ZN(W20019));
  NANDX1 G27467 (.A1(I1980), .A2(W2117), .ZN(W3658));
  NANDX1 G27468 (.A1(W1909), .A2(W2640), .ZN(W3662));
  NANDX1 G27469 (.A1(W5555), .A2(W2495), .ZN(W20017));
  NANDX1 G27470 (.A1(W6223), .A2(W1330), .ZN(W20016));
  NANDX1 G27471 (.A1(W3286), .A2(W256), .ZN(W3664));
  NANDX1 G27472 (.A1(W4534), .A2(W6379), .ZN(W20025));
  NANDX1 G27473 (.A1(W2181), .A2(W287), .ZN(W3666));
  NANDX1 G27474 (.A1(I706), .A2(W2449), .ZN(W3667));
  NANDX1 G27475 (.A1(W15818), .A2(W7605), .ZN(O1909));
  NANDX1 G27476 (.A1(W519), .A2(I777), .ZN(W8504));
  NANDX1 G27477 (.A1(I690), .A2(I1638), .ZN(W20013));
  NANDX1 G27478 (.A1(W4733), .A2(W3792), .ZN(W8503));
  NANDX1 G27479 (.A1(W510), .A2(W3990), .ZN(W8502));
  NANDX1 G27480 (.A1(W10809), .A2(W4826), .ZN(O1908));
  NANDX1 G27481 (.A1(W4896), .A2(W6921), .ZN(O626));
  NANDX1 G27482 (.A1(W5190), .A2(W17480), .ZN(O1915));
  NANDX1 G27483 (.A1(I132), .A2(W5338), .ZN(O1914));
  NANDX1 G27484 (.A1(W12686), .A2(W7870), .ZN(W20046));
  NANDX1 G27485 (.A1(W18283), .A2(W4821), .ZN(W20044));
  NANDX1 G27486 (.A1(W16200), .A2(W1668), .ZN(W20041));
  NANDX1 G27487 (.A1(W10201), .A2(W2014), .ZN(O625));
  NANDX1 G27488 (.A1(W14668), .A2(W15703), .ZN(W20039));
  NANDX1 G27489 (.A1(W3119), .A2(W5852), .ZN(O1912));
  NANDX1 G27490 (.A1(W8962), .A2(W11605), .ZN(W12644));
  NANDX1 G27491 (.A1(W18618), .A2(W4967), .ZN(W20035));
  NANDX1 G27492 (.A1(W564), .A2(W966), .ZN(W8508));
  NANDX1 G27493 (.A1(W12305), .A2(W18260), .ZN(O1910));
  NANDX1 G27494 (.A1(W12291), .A2(W5068), .ZN(W12635));
  NANDX1 G27495 (.A1(W7684), .A2(W16679), .ZN(W20029));
  NANDX1 G27496 (.A1(W3520), .A2(I1264), .ZN(W8507));
  NANDX1 G27497 (.A1(W2751), .A2(I1013), .ZN(W3655));
  NANDX1 G27498 (.A1(W3023), .A2(W1008), .ZN(W8506));
  NANDX1 G27499 (.A1(W3473), .A2(I1088), .ZN(W3693));
  NANDX1 G27500 (.A1(W11576), .A2(W7119), .ZN(W12657));
  NANDX1 G27501 (.A1(W13060), .A2(W4485), .ZN(W19985));
  NANDX1 G27502 (.A1(W14122), .A2(W16375), .ZN(W25342));
  NANDX1 G27503 (.A1(W2558), .A2(W1548), .ZN(W12661));
  NANDX1 G27504 (.A1(W2447), .A2(W8181), .ZN(O233));
  NANDX1 G27505 (.A1(W11171), .A2(W1802), .ZN(W12667));
  NANDX1 G27506 (.A1(W10866), .A2(W15189), .ZN(O1903));
  NANDX1 G27507 (.A1(W9262), .A2(W8235), .ZN(W12668));
  NANDX1 G27508 (.A1(W11874), .A2(I1458), .ZN(W12656));
  NANDX1 G27509 (.A1(W1218), .A2(I745), .ZN(W3694));
  NANDX1 G27510 (.A1(W8420), .A2(W9974), .ZN(W19974));
  NANDX1 G27511 (.A1(W1399), .A2(W2476), .ZN(W3695));
  NANDX1 G27512 (.A1(W2615), .A2(W2634), .ZN(W3697));
  NANDX1 G27513 (.A1(W8887), .A2(W8943), .ZN(O630));
  NANDX1 G27514 (.A1(W1078), .A2(W1220), .ZN(W3699));
  NANDX1 G27515 (.A1(W3388), .A2(W15812), .ZN(O1900));
  NANDX1 G27516 (.A1(I874), .A2(I1216), .ZN(W3701));
  NANDX1 G27517 (.A1(W13458), .A2(W4970), .ZN(W19997));
  NANDX1 G27518 (.A1(W2590), .A2(W3349), .ZN(W20009));
  NANDX1 G27519 (.A1(W10816), .A2(W4345), .ZN(W20008));
  NANDX1 G27520 (.A1(W999), .A2(W1253), .ZN(W3673));
  NANDX1 G27521 (.A1(W17466), .A2(W1074), .ZN(W20006));
  NANDX1 G27522 (.A1(I166), .A2(W3039), .ZN(W3674));
  NANDX1 G27523 (.A1(I1639), .A2(W9359), .ZN(W20004));
  NANDX1 G27524 (.A1(W1908), .A2(W7286), .ZN(W12645));
  NANDX1 G27525 (.A1(W7232), .A2(W6275), .ZN(W12646));
  NANDX1 G27526 (.A1(W4099), .A2(W7521), .ZN(W12696));
  NANDX1 G27527 (.A1(W10013), .A2(W11291), .ZN(W12650));
  NANDX1 G27528 (.A1(W129), .A2(W1385), .ZN(W3677));
  NANDX1 G27529 (.A1(W9070), .A2(W8660), .ZN(O1905));
  NANDX1 G27530 (.A1(W10910), .A2(W5325), .ZN(O628));
  NANDX1 G27531 (.A1(W5682), .A2(W305), .ZN(W8497));
  NANDX1 G27532 (.A1(I12), .A2(W5449), .ZN(W12652));
  NANDX1 G27533 (.A1(W12363), .A2(I268), .ZN(W19989));
  NANDX1 G27534 (.A1(W1604), .A2(I1800), .ZN(W8495));
  NANDX1 G27535 (.A1(W1340), .A2(I1529), .ZN(W3841));
  NANDX1 G27536 (.A1(W6665), .A2(W16568), .ZN(O1847));
  NANDX1 G27537 (.A1(W4963), .A2(W4628), .ZN(O645));
  NANDX1 G27538 (.A1(W2965), .A2(W5254), .ZN(W19765));
  NANDX1 G27539 (.A1(I1197), .A2(W4358), .ZN(W12761));
  NANDX1 G27540 (.A1(W3251), .A2(W16544), .ZN(W19764));
  NANDX1 G27541 (.A1(I1820), .A2(W6183), .ZN(W8420));
  NANDX1 G27542 (.A1(W879), .A2(I257), .ZN(W19761));
  NANDX1 G27543 (.A1(W8435), .A2(I1938), .ZN(W12762));
  NANDX1 G27544 (.A1(I1666), .A2(W5247), .ZN(W19759));
  NANDX1 G27545 (.A1(W3800), .A2(W4210), .ZN(W8422));
  NANDX1 G27546 (.A1(W2106), .A2(W1256), .ZN(W3842));
  NANDX1 G27547 (.A1(W8737), .A2(W10846), .ZN(W19757));
  NANDX1 G27548 (.A1(W6706), .A2(W11836), .ZN(O1846));
  NANDX1 G27549 (.A1(W19390), .A2(W6335), .ZN(W19753));
  NANDX1 G27550 (.A1(W14247), .A2(W13473), .ZN(W19751));
  NANDX1 G27551 (.A1(W2900), .A2(I1709), .ZN(O1843));
  NANDX1 G27552 (.A1(W1298), .A2(W6159), .ZN(W8417));
  NANDX1 G27553 (.A1(W10141), .A2(W14844), .ZN(W19745));
  NANDX1 G27554 (.A1(W5276), .A2(W6247), .ZN(W19787));
  NANDX1 G27555 (.A1(I1031), .A2(I827), .ZN(W8430));
  NANDX1 G27556 (.A1(I1271), .A2(W1599), .ZN(W3824));
  NANDX1 G27557 (.A1(W8689), .A2(W9445), .ZN(W19792));
  NANDX1 G27558 (.A1(W2388), .A2(I81), .ZN(W3825));
  NANDX1 G27559 (.A1(W4727), .A2(W11313), .ZN(W12745));
  NANDX1 G27560 (.A1(W615), .A2(W6109), .ZN(W12746));
  NANDX1 G27561 (.A1(W6130), .A2(W5438), .ZN(W12747));
  NANDX1 G27562 (.A1(W1262), .A2(W530), .ZN(W12748));
  NANDX1 G27563 (.A1(W17850), .A2(W3799), .ZN(W19744));
  NANDX1 G27564 (.A1(W9761), .A2(W5071), .ZN(W12749));
  NANDX1 G27565 (.A1(W3599), .A2(I675), .ZN(W12751));
  NANDX1 G27566 (.A1(W7511), .A2(W5496), .ZN(W8425));
  NANDX1 G27567 (.A1(W2201), .A2(W2471), .ZN(O46));
  NANDX1 G27568 (.A1(W4560), .A2(W11143), .ZN(O1850));
  NANDX1 G27569 (.A1(W13373), .A2(W19286), .ZN(W19780));
  NANDX1 G27570 (.A1(W10), .A2(W10487), .ZN(W19773));
  NANDX1 G27571 (.A1(W1557), .A2(W9256), .ZN(W12756));
  NANDX1 G27572 (.A1(W2728), .A2(W3707), .ZN(W3869));
  NANDX1 G27573 (.A1(W2938), .A2(W6349), .ZN(W12787));
  NANDX1 G27574 (.A1(I1021), .A2(I98), .ZN(W19714));
  NANDX1 G27575 (.A1(W7833), .A2(W18495), .ZN(W19713));
  NANDX1 G27576 (.A1(W760), .A2(W8822), .ZN(W12789));
  NANDX1 G27577 (.A1(W2405), .A2(W1226), .ZN(W3867));
  NANDX1 G27578 (.A1(W17220), .A2(W10513), .ZN(W19712));
  NANDX1 G27579 (.A1(W2783), .A2(W547), .ZN(W3868));
  NANDX1 G27580 (.A1(I1824), .A2(W13873), .ZN(O1832));
  NANDX1 G27581 (.A1(W3988), .A2(W2383), .ZN(O650));
  NANDX1 G27582 (.A1(W5182), .A2(W6736), .ZN(W12790));
  NANDX1 G27583 (.A1(W12021), .A2(W4851), .ZN(W19708));
  NANDX1 G27584 (.A1(W1595), .A2(W1500), .ZN(W12791));
  NANDX1 G27585 (.A1(W2297), .A2(W16441), .ZN(O1830));
  NANDX1 G27586 (.A1(W116), .A2(W2466), .ZN(W3879));
  NANDX1 G27587 (.A1(I846), .A2(W679), .ZN(W3880));
  NANDX1 G27588 (.A1(W14377), .A2(I1957), .ZN(O1829));
  NANDX1 G27589 (.A1(I12), .A2(I1299), .ZN(W3888));
  NANDX1 G27590 (.A1(I1013), .A2(W6878), .ZN(W8415));
  NANDX1 G27591 (.A1(W8135), .A2(W17102), .ZN(W19742));
  NANDX1 G27592 (.A1(W17540), .A2(W5656), .ZN(W19741));
  NANDX1 G27593 (.A1(W10032), .A2(W10385), .ZN(W12765));
  NANDX1 G27594 (.A1(W10978), .A2(W3606), .ZN(W12771));
  NANDX1 G27595 (.A1(W12362), .A2(W4369), .ZN(W12772));
  NANDX1 G27596 (.A1(W2734), .A2(I1216), .ZN(W3844));
  NANDX1 G27597 (.A1(W17519), .A2(I312), .ZN(W19735));
  NANDX1 G27598 (.A1(W8484), .A2(W1690), .ZN(W12777));
  NANDX1 G27599 (.A1(W3087), .A2(W1419), .ZN(W3819));
  NANDX1 G27600 (.A1(I1175), .A2(W535), .ZN(W12779));
  NANDX1 G27601 (.A1(W2171), .A2(W1322), .ZN(W3848));
  NANDX1 G27602 (.A1(W7433), .A2(W2933), .ZN(W12782));
  NANDX1 G27603 (.A1(W4034), .A2(W10793), .ZN(O1834));
  NANDX1 G27604 (.A1(W12876), .A2(W6842), .ZN(W19725));
  NANDX1 G27605 (.A1(W2629), .A2(W1201), .ZN(W12785));
  NANDX1 G27606 (.A1(W372), .A2(W48), .ZN(W3857));
  NANDX1 G27607 (.A1(I330), .A2(W2101), .ZN(W3860));
  NANDX1 G27608 (.A1(W13883), .A2(W9054), .ZN(W19844));
  NANDX1 G27609 (.A1(W3915), .A2(I1955), .ZN(W8450));
  NANDX1 G27610 (.A1(W17356), .A2(W18675), .ZN(W19853));
  NANDX1 G27611 (.A1(W17543), .A2(I1172), .ZN(W19850));
  NANDX1 G27612 (.A1(W17907), .A2(W15008), .ZN(W19848));
  NANDX1 G27613 (.A1(I1809), .A2(W2646), .ZN(W12707));
  NANDX1 G27614 (.A1(W2075), .A2(I924), .ZN(W3772));
  NANDX1 G27615 (.A1(W10132), .A2(W3643), .ZN(W12708));
  NANDX1 G27616 (.A1(I1386), .A2(I1851), .ZN(W8447));
  NANDX1 G27617 (.A1(W4882), .A2(W6814), .ZN(O637));
  NANDX1 G27618 (.A1(W3734), .A2(W869), .ZN(W3770));
  NANDX1 G27619 (.A1(W2407), .A2(W193), .ZN(W12715));
  NANDX1 G27620 (.A1(W306), .A2(W3400), .ZN(W3779));
  NANDX1 G27621 (.A1(I966), .A2(W3078), .ZN(W3780));
  NANDX1 G27622 (.A1(W1422), .A2(W7570), .ZN(W12716));
  NANDX1 G27623 (.A1(W16646), .A2(W17113), .ZN(W19842));
  NANDX1 G27624 (.A1(W3039), .A2(W209), .ZN(W19840));
  NANDX1 G27625 (.A1(W1413), .A2(W1626), .ZN(W3784));
  NANDX1 G27626 (.A1(W7288), .A2(W134), .ZN(W12721));
  NANDX1 G27627 (.A1(W15932), .A2(W12205), .ZN(W19865));
  NANDX1 G27628 (.A1(I220), .A2(W443), .ZN(W3758));
  NANDX1 G27629 (.A1(W6602), .A2(W10694), .ZN(W19873));
  NANDX1 G27630 (.A1(W644), .A2(W4920), .ZN(O636));
  NANDX1 G27631 (.A1(W2793), .A2(W1383), .ZN(W8453));
  NANDX1 G27632 (.A1(I1160), .A2(I1206), .ZN(W8452));
  NANDX1 G27633 (.A1(W4736), .A2(W3769), .ZN(W19869));
  NANDX1 G27634 (.A1(I1886), .A2(W2445), .ZN(W3762));
  NANDX1 G27635 (.A1(W2769), .A2(W11283), .ZN(W19867));
  NANDX1 G27636 (.A1(W3329), .A2(W2981), .ZN(O228));
  NANDX1 G27637 (.A1(W2823), .A2(W3318), .ZN(W3763));
  NANDX1 G27638 (.A1(W2842), .A2(I1935), .ZN(W8451));
  NANDX1 G27639 (.A1(W19054), .A2(W8921), .ZN(O1871));
  NANDX1 G27640 (.A1(I597), .A2(W939), .ZN(W3765));
  NANDX1 G27641 (.A1(W10098), .A2(W4885), .ZN(O1870));
  NANDX1 G27642 (.A1(W2142), .A2(W2892), .ZN(W3766));
  NANDX1 G27643 (.A1(I46), .A2(I764), .ZN(W3767));
  NANDX1 G27644 (.A1(I1519), .A2(I1393), .ZN(W3769));
  NANDX1 G27645 (.A1(W1717), .A2(I654), .ZN(W3813));
  NANDX1 G27646 (.A1(W93), .A2(W5956), .ZN(W8433));
  NANDX1 G27647 (.A1(W6877), .A2(W8944), .ZN(W19807));
  NANDX1 G27648 (.A1(W11606), .A2(W1295), .ZN(W19806));
  NANDX1 G27649 (.A1(W1118), .A2(W19684), .ZN(W19805));
  NANDX1 G27650 (.A1(I743), .A2(W7293), .ZN(O642));
  NANDX1 G27651 (.A1(W4634), .A2(W12724), .ZN(W12734));
  NANDX1 G27652 (.A1(I679), .A2(I1122), .ZN(W3809));
  NANDX1 G27653 (.A1(W1767), .A2(W2050), .ZN(W3812));
  NANDX1 G27654 (.A1(W5778), .A2(W5401), .ZN(W12731));
  NANDX1 G27655 (.A1(W16617), .A2(W5936), .ZN(W19802));
  NANDX1 G27656 (.A1(W770), .A2(W3138), .ZN(W3815));
  NANDX1 G27657 (.A1(W8862), .A2(I1707), .ZN(W19800));
  NANDX1 G27658 (.A1(W2840), .A2(W2422), .ZN(W3817));
  NANDX1 G27659 (.A1(W10549), .A2(I1283), .ZN(O1857));
  NANDX1 G27660 (.A1(W12564), .A2(W10310), .ZN(W12738));
  NANDX1 G27661 (.A1(W11819), .A2(W5903), .ZN(W12741));
  NANDX1 G27662 (.A1(W3015), .A2(I1160), .ZN(W3818));
  NANDX1 G27663 (.A1(W122), .A2(W3535), .ZN(W3799));
  NANDX1 G27664 (.A1(W2211), .A2(W2704), .ZN(W12724));
  NANDX1 G27665 (.A1(W2922), .A2(W1832), .ZN(O44));
  NANDX1 G27666 (.A1(W12362), .A2(W11584), .ZN(W19834));
  NANDX1 G27667 (.A1(W16538), .A2(W5577), .ZN(W19832));
  NANDX1 G27668 (.A1(W14143), .A2(W7109), .ZN(O1865));
  NANDX1 G27669 (.A1(W2094), .A2(I740), .ZN(W3794));
  NANDX1 G27670 (.A1(W7736), .A2(W19704), .ZN(W19828));
  NANDX1 G27671 (.A1(W809), .A2(W3428), .ZN(W8440));
  NANDX1 G27672 (.A1(W2353), .A2(W3460), .ZN(W5101));
  NANDX1 G27673 (.A1(I1510), .A2(W9175), .ZN(W19821));
  NANDX1 G27674 (.A1(W18499), .A2(I486), .ZN(O1863));
  NANDX1 G27675 (.A1(W104), .A2(W10760), .ZN(W19814));
  NANDX1 G27676 (.A1(W354), .A2(W11260), .ZN(W12728));
  NANDX1 G27677 (.A1(W6751), .A2(I690), .ZN(W8438));
  NANDX1 G27678 (.A1(W7447), .A2(W5997), .ZN(W8437));
  NANDX1 G27679 (.A1(W10067), .A2(W18047), .ZN(O1860));
  NANDX1 G27680 (.A1(W11630), .A2(W14710), .ZN(W19808));
  NANDX1 G27681 (.A1(W11157), .A2(W14126), .ZN(O1091));
  NANDX1 G27682 (.A1(W3542), .A2(W6144), .ZN(W6376));
  NANDX1 G27683 (.A1(W3169), .A2(W3145), .ZN(W6377));
  NANDX1 G27684 (.A1(W13363), .A2(W11), .ZN(W14518));
  NANDX1 G27685 (.A1(W2516), .A2(I921), .ZN(W7252));
  NANDX1 G27686 (.A1(W494), .A2(W3671), .ZN(W6379));
  NANDX1 G27687 (.A1(W1734), .A2(W13275), .ZN(O1092));
  NANDX1 G27688 (.A1(W13951), .A2(W6610), .ZN(W15918));
  NANDX1 G27689 (.A1(W12860), .A2(W3985), .ZN(W15917));
  NANDX1 G27690 (.A1(W2487), .A2(W6877), .ZN(W7248));
  NANDX1 G27691 (.A1(W5449), .A2(W9741), .ZN(W15928));
  NANDX1 G27692 (.A1(W220), .A2(I1079), .ZN(W6382));
  NANDX1 G27693 (.A1(W4463), .A2(W32), .ZN(W6384));
  NANDX1 G27694 (.A1(W3012), .A2(W2920), .ZN(O1090));
  NANDX1 G27695 (.A1(W10073), .A2(W8499), .ZN(W14522));
  NANDX1 G27696 (.A1(W14512), .A2(W3790), .ZN(W15907));
  NANDX1 G27697 (.A1(W5755), .A2(W663), .ZN(W7246));
  NANDX1 G27698 (.A1(W5665), .A2(W9540), .ZN(W14525));
  NANDX1 G27699 (.A1(W6380), .A2(W682), .ZN(W6393));
  NANDX1 G27700 (.A1(W1388), .A2(W5711), .ZN(W14499));
  NANDX1 G27701 (.A1(W11601), .A2(W5976), .ZN(W15952));
  NANDX1 G27702 (.A1(W6856), .A2(W4051), .ZN(W15951));
  NANDX1 G27703 (.A1(W5890), .A2(W3780), .ZN(W6349));
  NANDX1 G27704 (.A1(I1114), .A2(W361), .ZN(W7272));
  NANDX1 G27705 (.A1(W13420), .A2(W539), .ZN(W14493));
  NANDX1 G27706 (.A1(W14723), .A2(W9808), .ZN(W15946));
  NANDX1 G27707 (.A1(W6132), .A2(W193), .ZN(W6353));
  NANDX1 G27708 (.A1(W1360), .A2(I348), .ZN(W6359));
  NANDX1 G27709 (.A1(W795), .A2(W11481), .ZN(W15902));
  NANDX1 G27710 (.A1(W4387), .A2(W13000), .ZN(W14501));
  NANDX1 G27711 (.A1(W5116), .A2(W2009), .ZN(W6368));
  NANDX1 G27712 (.A1(W8765), .A2(W4732), .ZN(O879));
  NANDX1 G27713 (.A1(W11818), .A2(W4000), .ZN(W14510));
  NANDX1 G27714 (.A1(W380), .A2(W6964), .ZN(W14514));
  NANDX1 G27715 (.A1(W6904), .A2(I394), .ZN(W7260));
  NANDX1 G27716 (.A1(I72), .A2(W9029), .ZN(W15930));
  NANDX1 G27717 (.A1(W9818), .A2(W1858), .ZN(W15929));
  NANDX1 G27718 (.A1(I488), .A2(W11679), .ZN(O1077));
  NANDX1 G27719 (.A1(W5756), .A2(W6892), .ZN(W15871));
  NANDX1 G27720 (.A1(W4038), .A2(W737), .ZN(W15870));
  NANDX1 G27721 (.A1(W40), .A2(W1330), .ZN(W15869));
  NANDX1 G27722 (.A1(W4554), .A2(W1534), .ZN(O1080));
  NANDX1 G27723 (.A1(W13097), .A2(W8838), .ZN(W15864));
  NANDX1 G27724 (.A1(W4703), .A2(W8858), .ZN(W15863));
  NANDX1 G27725 (.A1(W7041), .A2(W11060), .ZN(W15862));
  NANDX1 G27726 (.A1(W2767), .A2(W10325), .ZN(W14536));
  NANDX1 G27727 (.A1(W579), .A2(W4344), .ZN(W6411));
  NANDX1 G27728 (.A1(W8667), .A2(W3241), .ZN(O1081));
  NANDX1 G27729 (.A1(W8191), .A2(W6241), .ZN(W15856));
  NANDX1 G27730 (.A1(W7117), .A2(W14709), .ZN(W15854));
  NANDX1 G27731 (.A1(W10798), .A2(I122), .ZN(W15853));
  NANDX1 G27732 (.A1(W828), .A2(W2158), .ZN(W6412));
  NANDX1 G27733 (.A1(W3772), .A2(W3274), .ZN(W6413));
  NANDX1 G27734 (.A1(W190), .A2(W12765), .ZN(W14539));
  NANDX1 G27735 (.A1(W2516), .A2(W14412), .ZN(O1075));
  NANDX1 G27736 (.A1(W4457), .A2(W1504), .ZN(W6415));
  NANDX1 G27737 (.A1(W3893), .A2(W10324), .ZN(O1086));
  NANDX1 G27738 (.A1(W3981), .A2(W4712), .ZN(W6398));
  NANDX1 G27739 (.A1(W9492), .A2(I895), .ZN(W14528));
  NANDX1 G27740 (.A1(W14878), .A2(W8134), .ZN(W15898));
  NANDX1 G27741 (.A1(W6798), .A2(W602), .ZN(W7243));
  NANDX1 G27742 (.A1(W5615), .A2(W6627), .ZN(W15894));
  NANDX1 G27743 (.A1(W3417), .A2(I873), .ZN(W7242));
  NANDX1 G27744 (.A1(W844), .A2(W3251), .ZN(W6404));
  NANDX1 G27745 (.A1(W6331), .A2(W5056), .ZN(W15891));
  NANDX1 G27746 (.A1(I1714), .A2(W4687), .ZN(W7273));
  NANDX1 G27747 (.A1(W4492), .A2(W13186), .ZN(W15888));
  NANDX1 G27748 (.A1(W7989), .A2(W10866), .ZN(W14533));
  NANDX1 G27749 (.A1(W6680), .A2(W6950), .ZN(W7241));
  NANDX1 G27750 (.A1(W3387), .A2(W13688), .ZN(W15882));
  NANDX1 G27751 (.A1(W4136), .A2(W209), .ZN(W6406));
  NANDX1 G27752 (.A1(W3968), .A2(W5034), .ZN(W15879));
  NANDX1 G27753 (.A1(W2743), .A2(W3625), .ZN(O1083));
  NANDX1 G27754 (.A1(W9936), .A2(W2749), .ZN(W15876));
  NANDX1 G27755 (.A1(W6397), .A2(W670), .ZN(W14474));
  NANDX1 G27756 (.A1(W3484), .A2(W2343), .ZN(W7290));
  NANDX1 G27757 (.A1(W1150), .A2(W14488), .ZN(O1102));
  NANDX1 G27758 (.A1(I446), .A2(W7196), .ZN(W7288));
  NANDX1 G27759 (.A1(W2270), .A2(W12063), .ZN(W14472));
  NANDX1 G27760 (.A1(W1945), .A2(W2352), .ZN(O128));
  NANDX1 G27761 (.A1(W4761), .A2(I1272), .ZN(W6307));
  NANDX1 G27762 (.A1(W13546), .A2(W4466), .ZN(W14473));
  NANDX1 G27763 (.A1(W1800), .A2(W5683), .ZN(W6308));
  NANDX1 G27764 (.A1(I1253), .A2(W12859), .ZN(O1101));
  NANDX1 G27765 (.A1(W1396), .A2(W1615), .ZN(W7291));
  NANDX1 G27766 (.A1(W12408), .A2(W6619), .ZN(W15995));
  NANDX1 G27767 (.A1(W4342), .A2(W5004), .ZN(W7283));
  NANDX1 G27768 (.A1(W5399), .A2(W14044), .ZN(W15994));
  NANDX1 G27769 (.A1(I51), .A2(W1586), .ZN(W6316));
  NANDX1 G27770 (.A1(W15619), .A2(W10259), .ZN(O1100));
  NANDX1 G27771 (.A1(W885), .A2(W4604), .ZN(W15989));
  NANDX1 G27772 (.A1(W4821), .A2(I350), .ZN(W6317));
  NANDX1 G27773 (.A1(I1770), .A2(W3896), .ZN(W6318));
  NANDX1 G27774 (.A1(W12701), .A2(W6461), .ZN(W16023));
  NANDX1 G27775 (.A1(W8546), .A2(W7487), .ZN(W14455));
  NANDX1 G27776 (.A1(W5614), .A2(W7406), .ZN(W14456));
  NANDX1 G27777 (.A1(W2696), .A2(W6889), .ZN(W14458));
  NANDX1 G27778 (.A1(W5414), .A2(W4713), .ZN(O126));
  NANDX1 G27779 (.A1(W5363), .A2(W3168), .ZN(W6283));
  NANDX1 G27780 (.A1(W612), .A2(W3039), .ZN(W6284));
  NANDX1 G27781 (.A1(W7961), .A2(W10353), .ZN(W14460));
  NANDX1 G27782 (.A1(W9402), .A2(W12695), .ZN(O1109));
  NANDX1 G27783 (.A1(W2750), .A2(I1862), .ZN(W6320));
  NANDX1 G27784 (.A1(W95), .A2(W4440), .ZN(W6288));
  NANDX1 G27785 (.A1(W8198), .A2(I168), .ZN(W16018));
  NANDX1 G27786 (.A1(W4024), .A2(I697), .ZN(W6289));
  NANDX1 G27787 (.A1(W3446), .A2(W1244), .ZN(W6290));
  NANDX1 G27788 (.A1(W507), .A2(I1338), .ZN(W6291));
  NANDX1 G27789 (.A1(W2988), .A2(I1630), .ZN(W6295));
  NANDX1 G27790 (.A1(W9691), .A2(W7138), .ZN(W14461));
  NANDX1 G27791 (.A1(W3695), .A2(W1381), .ZN(W7292));
  NANDX1 G27792 (.A1(W6158), .A2(W1245), .ZN(W7278));
  NANDX1 G27793 (.A1(W3909), .A2(W5873), .ZN(W6335));
  NANDX1 G27794 (.A1(W6420), .A2(W9711), .ZN(O1096));
  NANDX1 G27795 (.A1(I216), .A2(W6198), .ZN(W7280));
  NANDX1 G27796 (.A1(W7109), .A2(I1302), .ZN(W14485));
  NANDX1 G27797 (.A1(W8688), .A2(I1462), .ZN(W15963));
  NANDX1 G27798 (.A1(W7311), .A2(W13173), .ZN(W15962));
  NANDX1 G27799 (.A1(I1259), .A2(W5251), .ZN(W6338));
  NANDX1 G27800 (.A1(W1506), .A2(W3919), .ZN(W6340));
  NANDX1 G27801 (.A1(W13449), .A2(W14393), .ZN(W14484));
  NANDX1 G27802 (.A1(W4033), .A2(W9318), .ZN(W15958));
  NANDX1 G27803 (.A1(W965), .A2(W4018), .ZN(W14488));
  NANDX1 G27804 (.A1(I1274), .A2(I1640), .ZN(W7275));
  NANDX1 G27805 (.A1(W1387), .A2(W5739), .ZN(O876));
  NANDX1 G27806 (.A1(W1891), .A2(I531), .ZN(W6346));
  NANDX1 G27807 (.A1(W6575), .A2(W12417), .ZN(W15956));
  NANDX1 G27808 (.A1(W2398), .A2(W5605), .ZN(W6347));
  NANDX1 G27809 (.A1(I1110), .A2(W3885), .ZN(W6348));
  NANDX1 G27810 (.A1(W364), .A2(W3250), .ZN(W6328));
  NANDX1 G27811 (.A1(W8223), .A2(W8120), .ZN(W14476));
  NANDX1 G27812 (.A1(W509), .A2(I420), .ZN(W6321));
  NANDX1 G27813 (.A1(W11115), .A2(W8186), .ZN(W14477));
  NANDX1 G27814 (.A1(W1763), .A2(W1464), .ZN(O1098));
  NANDX1 G27815 (.A1(I1348), .A2(I1755), .ZN(W6322));
  NANDX1 G27816 (.A1(W2771), .A2(I970), .ZN(W15982));
  NANDX1 G27817 (.A1(W5556), .A2(W4061), .ZN(W6323));
  NANDX1 G27818 (.A1(W13203), .A2(W5398), .ZN(W14478));
  NANDX1 G27819 (.A1(W13443), .A2(W8736), .ZN(W15845));
  NANDX1 G27820 (.A1(W370), .A2(W7154), .ZN(W14479));
  NANDX1 G27821 (.A1(W5710), .A2(W6061), .ZN(W6331));
  NANDX1 G27822 (.A1(W10239), .A2(W6011), .ZN(W15976));
  NANDX1 G27823 (.A1(W2645), .A2(W4116), .ZN(W6332));
  NANDX1 G27824 (.A1(W12993), .A2(W9547), .ZN(W14482));
  NANDX1 G27825 (.A1(W14005), .A2(W3617), .ZN(W15972));
  NANDX1 G27826 (.A1(W12921), .A2(W8804), .ZN(W15971));
  NANDX1 G27827 (.A1(W9872), .A2(W13366), .ZN(W15969));
  NANDX1 G27828 (.A1(W11800), .A2(W5043), .ZN(W15726));
  NANDX1 G27829 (.A1(W2953), .A2(W7504), .ZN(W15744));
  NANDX1 G27830 (.A1(I1119), .A2(W5230), .ZN(W7214));
  NANDX1 G27831 (.A1(W3751), .A2(W4538), .ZN(W6489));
  NANDX1 G27832 (.A1(W14036), .A2(W3053), .ZN(W15739));
  NANDX1 G27833 (.A1(W13294), .A2(W11688), .ZN(W15737));
  NANDX1 G27834 (.A1(W11132), .A2(W1088), .ZN(W15734));
  NANDX1 G27835 (.A1(W5265), .A2(W5889), .ZN(W7211));
  NANDX1 G27836 (.A1(W3207), .A2(I1634), .ZN(W6493));
  NANDX1 G27837 (.A1(I610), .A2(W15372), .ZN(W15728));
  NANDX1 G27838 (.A1(W500), .A2(W10412), .ZN(W15746));
  NANDX1 G27839 (.A1(W1878), .A2(W2684), .ZN(W7210));
  NANDX1 G27840 (.A1(W2006), .A2(W5158), .ZN(W6494));
  NANDX1 G27841 (.A1(W2083), .A2(W6109), .ZN(W6496));
  NANDX1 G27842 (.A1(W5580), .A2(W15557), .ZN(W15721));
  NANDX1 G27843 (.A1(W4545), .A2(W12794), .ZN(O886));
  NANDX1 G27844 (.A1(W15027), .A2(W3019), .ZN(O1056));
  NANDX1 G27845 (.A1(I1800), .A2(I1075), .ZN(O1055));
  NANDX1 G27846 (.A1(W4025), .A2(I2), .ZN(W7208));
  NANDX1 G27847 (.A1(I165), .A2(W4804), .ZN(W6482));
  NANDX1 G27848 (.A1(W7210), .A2(W3001), .ZN(O1064));
  NANDX1 G27849 (.A1(W11533), .A2(W8964), .ZN(O1063));
  NANDX1 G27850 (.A1(W14345), .A2(W307), .ZN(W15765));
  NANDX1 G27851 (.A1(W11947), .A2(W4438), .ZN(W15762));
  NANDX1 G27852 (.A1(W1433), .A2(W1734), .ZN(O1062));
  NANDX1 G27853 (.A1(W165), .A2(I1072), .ZN(W15756));
  NANDX1 G27854 (.A1(W11895), .A2(W3487), .ZN(W15755));
  NANDX1 G27855 (.A1(I316), .A2(I864), .ZN(W14572));
  NANDX1 G27856 (.A1(W3487), .A2(W4783), .ZN(W15717));
  NANDX1 G27857 (.A1(W14679), .A2(W2507), .ZN(W15751));
  NANDX1 G27858 (.A1(W6187), .A2(W1794), .ZN(W14573));
  NANDX1 G27859 (.A1(W2559), .A2(W6583), .ZN(W15750));
  NANDX1 G27860 (.A1(W14297), .A2(W4976), .ZN(W15749));
  NANDX1 G27861 (.A1(W14851), .A2(I477), .ZN(O1061));
  NANDX1 G27862 (.A1(W5695), .A2(W1351), .ZN(W6485));
  NANDX1 G27863 (.A1(W2547), .A2(I278), .ZN(W6486));
  NANDX1 G27864 (.A1(W4480), .A2(W12455), .ZN(W14578));
  NANDX1 G27865 (.A1(W13604), .A2(W12139), .ZN(W15674));
  NANDX1 G27866 (.A1(I1072), .A2(W455), .ZN(W14597));
  NANDX1 G27867 (.A1(W1543), .A2(W13266), .ZN(W15685));
  NANDX1 G27868 (.A1(W978), .A2(W8435), .ZN(W15684));
  NANDX1 G27869 (.A1(W1529), .A2(W2894), .ZN(W6512));
  NANDX1 G27870 (.A1(I544), .A2(W3508), .ZN(W15681));
  NANDX1 G27871 (.A1(W1947), .A2(W1128), .ZN(W6514));
  NANDX1 G27872 (.A1(W6673), .A2(W3781), .ZN(W7198));
  NANDX1 G27873 (.A1(W691), .A2(W161), .ZN(O1049));
  NANDX1 G27874 (.A1(W8270), .A2(W2846), .ZN(W15689));
  NANDX1 G27875 (.A1(W12653), .A2(W6663), .ZN(W15673));
  NANDX1 G27876 (.A1(W873), .A2(W4109), .ZN(W14603));
  NANDX1 G27877 (.A1(W1111), .A2(W2935), .ZN(W6516));
  NANDX1 G27878 (.A1(I975), .A2(W12706), .ZN(W15669));
  NANDX1 G27879 (.A1(W3383), .A2(W3189), .ZN(W6518));
  NANDX1 G27880 (.A1(W5371), .A2(W1738), .ZN(O1047));
  NANDX1 G27881 (.A1(W3612), .A2(W5880), .ZN(W6522));
  NANDX1 G27882 (.A1(I884), .A2(W5236), .ZN(W6523));
  NANDX1 G27883 (.A1(W142), .A2(W9259), .ZN(W14594));
  NANDX1 G27884 (.A1(I1468), .A2(W5039), .ZN(W6498));
  NANDX1 G27885 (.A1(I1325), .A2(W987), .ZN(W15714));
  NANDX1 G27886 (.A1(I750), .A2(I1143), .ZN(W15710));
  NANDX1 G27887 (.A1(W4798), .A2(W4084), .ZN(W15708));
  NANDX1 G27888 (.A1(W189), .A2(W3202), .ZN(W6500));
  NANDX1 G27889 (.A1(W3033), .A2(W10661), .ZN(W15706));
  NANDX1 G27890 (.A1(W13053), .A2(W12602), .ZN(W14590));
  NANDX1 G27891 (.A1(W14060), .A2(W14199), .ZN(W15701));
  NANDX1 G27892 (.A1(W6097), .A2(W1128), .ZN(W6479));
  NANDX1 G27893 (.A1(W1249), .A2(W2566), .ZN(W14596));
  NANDX1 G27894 (.A1(W1909), .A2(W24), .ZN(W6507));
  NANDX1 G27895 (.A1(W1793), .A2(W6196), .ZN(W7200));
  NANDX1 G27896 (.A1(W4471), .A2(W763), .ZN(W6508));
  NANDX1 G27897 (.A1(W8083), .A2(W10579), .ZN(W15693));
  NANDX1 G27898 (.A1(W6030), .A2(W2377), .ZN(W15692));
  NANDX1 G27899 (.A1(W2325), .A2(W13675), .ZN(O1051));
  NANDX1 G27900 (.A1(W3740), .A2(I1282), .ZN(W6511));
  NANDX1 G27901 (.A1(W4630), .A2(W6562), .ZN(W7228));
  NANDX1 G27902 (.A1(W12842), .A2(W6413), .ZN(O1071));
  NANDX1 G27903 (.A1(W5345), .A2(W5222), .ZN(W6437));
  NANDX1 G27904 (.A1(W7825), .A2(W1543), .ZN(W15820));
  NANDX1 G27905 (.A1(W11705), .A2(W1848), .ZN(W14545));
  NANDX1 G27906 (.A1(I1154), .A2(I68), .ZN(W6439));
  NANDX1 G27907 (.A1(I1546), .A2(W14478), .ZN(W14546));
  NANDX1 G27908 (.A1(W2277), .A2(I657), .ZN(W6440));
  NANDX1 G27909 (.A1(I374), .A2(W3824), .ZN(W7229));
  NANDX1 G27910 (.A1(W4125), .A2(I424), .ZN(W6441));
  NANDX1 G27911 (.A1(W1265), .A2(W14384), .ZN(W14543));
  NANDX1 G27912 (.A1(I610), .A2(W273), .ZN(W6443));
  NANDX1 G27913 (.A1(W3209), .A2(I1780), .ZN(W6444));
  NANDX1 G27914 (.A1(W10504), .A2(W11867), .ZN(W15810));
  NANDX1 G27915 (.A1(W10541), .A2(W5097), .ZN(W15809));
  NANDX1 G27916 (.A1(W1470), .A2(W5626), .ZN(W14549));
  NANDX1 G27917 (.A1(W12430), .A2(W8046), .ZN(W15807));
  NANDX1 G27918 (.A1(W3110), .A2(W7236), .ZN(W15806));
  NANDX1 G27919 (.A1(W10098), .A2(W5447), .ZN(W15805));
  NANDX1 G27920 (.A1(W5423), .A2(W3390), .ZN(W7231));
  NANDX1 G27921 (.A1(W6386), .A2(W4352), .ZN(W6416));
  NANDX1 G27922 (.A1(W143), .A2(W500), .ZN(W6417));
  NANDX1 G27923 (.A1(W206), .A2(W3982), .ZN(W6419));
  NANDX1 G27924 (.A1(I1453), .A2(W13127), .ZN(W15843));
  NANDX1 G27925 (.A1(I104), .A2(W5711), .ZN(W15840));
  NANDX1 G27926 (.A1(W10415), .A2(W10249), .ZN(W15839));
  NANDX1 G27927 (.A1(W1168), .A2(W1581), .ZN(W6420));
  NANDX1 G27928 (.A1(W1778), .A2(W4029), .ZN(O130));
  NANDX1 G27929 (.A1(W83), .A2(W8143), .ZN(W15804));
  NANDX1 G27930 (.A1(W3404), .A2(W3834), .ZN(W6424));
  NANDX1 G27931 (.A1(W3103), .A2(I219), .ZN(W6426));
  NANDX1 G27932 (.A1(I1553), .A2(W1292), .ZN(W6429));
  NANDX1 G27933 (.A1(W6232), .A2(W7986), .ZN(W15830));
  NANDX1 G27934 (.A1(W5525), .A2(W10437), .ZN(W14541));
  NANDX1 G27935 (.A1(W12754), .A2(W3902), .ZN(W15829));
  NANDX1 G27936 (.A1(W2992), .A2(W1867), .ZN(W6431));
  NANDX1 G27937 (.A1(W6897), .A2(W9811), .ZN(W15828));
  NANDX1 G27938 (.A1(W14547), .A2(W1479), .ZN(W14568));
  NANDX1 G27939 (.A1(I471), .A2(I282), .ZN(W6461));
  NANDX1 G27940 (.A1(W1125), .A2(W6234), .ZN(W6462));
  NANDX1 G27941 (.A1(W3852), .A2(W4634), .ZN(W6465));
  NANDX1 G27942 (.A1(W8456), .A2(W12280), .ZN(W15782));
  NANDX1 G27943 (.A1(I331), .A2(W4558), .ZN(W6466));
  NANDX1 G27944 (.A1(W2741), .A2(W6668), .ZN(W7222));
  NANDX1 G27945 (.A1(W2278), .A2(W14616), .ZN(O1066));
  NANDX1 G27946 (.A1(W5666), .A2(I1452), .ZN(W15778));
  NANDX1 G27947 (.A1(W3434), .A2(W3111), .ZN(W6460));
  NANDX1 G27948 (.A1(I64), .A2(W2316), .ZN(W15775));
  NANDX1 G27949 (.A1(W10117), .A2(I255), .ZN(W15774));
  NANDX1 G27950 (.A1(W9328), .A2(W2207), .ZN(W14569));
  NANDX1 G27951 (.A1(I1945), .A2(W13622), .ZN(W15772));
  NANDX1 G27952 (.A1(W2781), .A2(I65), .ZN(W6468));
  NANDX1 G27953 (.A1(W1448), .A2(W4186), .ZN(W6474));
  NANDX1 G27954 (.A1(I1396), .A2(W6208), .ZN(W7219));
  NANDX1 G27955 (.A1(W4411), .A2(W1435), .ZN(W6478));
  NANDX1 G27956 (.A1(W5761), .A2(W3811), .ZN(W14554));
  NANDX1 G27957 (.A1(W4358), .A2(W5638), .ZN(W14550));
  NANDX1 G27958 (.A1(W962), .A2(W12367), .ZN(W15801));
  NANDX1 G27959 (.A1(I1990), .A2(W5842), .ZN(W15800));
  NANDX1 G27960 (.A1(I871), .A2(W7722), .ZN(W14551));
  NANDX1 G27961 (.A1(W856), .A2(W10671), .ZN(O882));
  NANDX1 G27962 (.A1(I1384), .A2(W810), .ZN(O132));
  NANDX1 G27963 (.A1(W13417), .A2(W14379), .ZN(W15799));
  NANDX1 G27964 (.A1(W11771), .A2(W331), .ZN(W15797));
  NANDX1 G27965 (.A1(W3524), .A2(W3400), .ZN(W6277));
  NANDX1 G27966 (.A1(W4622), .A2(I71), .ZN(W14555));
  NANDX1 G27967 (.A1(W3710), .A2(I45), .ZN(W6453));
  NANDX1 G27968 (.A1(W6429), .A2(W7480), .ZN(W14556));
  NANDX1 G27969 (.A1(W5906), .A2(W14743), .ZN(W15793));
  NANDX1 G27970 (.A1(I887), .A2(W2031), .ZN(W6457));
  NANDX1 G27971 (.A1(I970), .A2(W7171), .ZN(W7224));
  NANDX1 G27972 (.A1(W3517), .A2(W13462), .ZN(W15786));
  NANDX1 G27973 (.A1(W2240), .A2(W641), .ZN(W6459));
  NANDX1 G27974 (.A1(W1309), .A2(W4602), .ZN(W7364));
  NANDX1 G27975 (.A1(W4763), .A2(W876), .ZN(W6124));
  NANDX1 G27976 (.A1(W8284), .A2(W7183), .ZN(W14367));
  NANDX1 G27977 (.A1(I1591), .A2(W48), .ZN(W16311));
  NANDX1 G27978 (.A1(W6081), .A2(I562), .ZN(O858));
  NANDX1 G27979 (.A1(W5793), .A2(W3943), .ZN(W6132));
  NANDX1 G27980 (.A1(W12157), .A2(W10953), .ZN(W14374));
  NANDX1 G27981 (.A1(I1909), .A2(W6954), .ZN(W16298));
  NANDX1 G27982 (.A1(W6428), .A2(W2124), .ZN(W7365));
  NANDX1 G27983 (.A1(W11146), .A2(W5422), .ZN(W16296));
  NANDX1 G27984 (.A1(W7053), .A2(W1896), .ZN(W7368));
  NANDX1 G27985 (.A1(I1361), .A2(W3440), .ZN(W6136));
  NANDX1 G27986 (.A1(W10356), .A2(W10373), .ZN(W14375));
  NANDX1 G27987 (.A1(W2389), .A2(I1062), .ZN(W16292));
  NANDX1 G27988 (.A1(W13229), .A2(W12920), .ZN(W14377));
  NANDX1 G27989 (.A1(W7224), .A2(W8934), .ZN(W16291));
  NANDX1 G27990 (.A1(I1437), .A2(W4522), .ZN(W6141));
  NANDX1 G27991 (.A1(W1475), .A2(W13686), .ZN(W14378));
  NANDX1 G27992 (.A1(I872), .A2(W4506), .ZN(W6144));
  NANDX1 G27993 (.A1(W13533), .A2(W10007), .ZN(W14360));
  NANDX1 G27994 (.A1(W6972), .A2(W16311), .ZN(W16339));
  NANDX1 G27995 (.A1(W11793), .A2(W7208), .ZN(W16338));
  NANDX1 G27996 (.A1(W10396), .A2(W14588), .ZN(W16336));
  NANDX1 G27997 (.A1(I1400), .A2(W2009), .ZN(W14356));
  NANDX1 G27998 (.A1(I661), .A2(W12345), .ZN(W14358));
  NANDX1 G27999 (.A1(W4326), .A2(W15018), .ZN(W16331));
  NANDX1 G28000 (.A1(I421), .A2(W5605), .ZN(W6114));
  NANDX1 G28001 (.A1(W4254), .A2(W5015), .ZN(W6118));
  NANDX1 G28002 (.A1(W2601), .A2(W1424), .ZN(W6149));
  NANDX1 G28003 (.A1(W5783), .A2(W5124), .ZN(O119));
  NANDX1 G28004 (.A1(W8038), .A2(W3600), .ZN(W14361));
  NANDX1 G28005 (.A1(W10620), .A2(W2935), .ZN(W16324));
  NANDX1 G28006 (.A1(I1550), .A2(W9876), .ZN(W16323));
  NANDX1 G28007 (.A1(W3313), .A2(W5259), .ZN(W16321));
  NANDX1 G28008 (.A1(W5456), .A2(W5476), .ZN(W6122));
  NANDX1 G28009 (.A1(W4865), .A2(W6174), .ZN(W16317));
  NANDX1 G28010 (.A1(W163), .A2(W1057), .ZN(W6123));
  NANDX1 G28011 (.A1(W3054), .A2(W2649), .ZN(W6176));
  NANDX1 G28012 (.A1(W12424), .A2(W441), .ZN(O1148));
  NANDX1 G28013 (.A1(W4104), .A2(W16184), .ZN(W16260));
  NANDX1 G28014 (.A1(W5939), .A2(W1348), .ZN(W16259));
  NANDX1 G28015 (.A1(W2383), .A2(W3892), .ZN(W6173));
  NANDX1 G28016 (.A1(W3971), .A2(W1981), .ZN(W6174));
  NANDX1 G28017 (.A1(W1247), .A2(W9758), .ZN(W16255));
  NANDX1 G28018 (.A1(I1491), .A2(I1975), .ZN(W6175));
  NANDX1 G28019 (.A1(W2836), .A2(W15717), .ZN(W16247));
  NANDX1 G28020 (.A1(W5776), .A2(W2484), .ZN(W14384));
  NANDX1 G28021 (.A1(W1182), .A2(W11225), .ZN(W16246));
  NANDX1 G28022 (.A1(W15036), .A2(W10230), .ZN(O1144));
  NANDX1 G28023 (.A1(I1236), .A2(W2369), .ZN(W7347));
  NANDX1 G28024 (.A1(W5482), .A2(W736), .ZN(W6179));
  NANDX1 G28025 (.A1(W1358), .A2(W1192), .ZN(W7346));
  NANDX1 G28026 (.A1(W1119), .A2(W4972), .ZN(O121));
  NANDX1 G28027 (.A1(W4838), .A2(I706), .ZN(W6181));
  NANDX1 G28028 (.A1(W5733), .A2(W9527), .ZN(W16232));
  NANDX1 G28029 (.A1(W4146), .A2(W3064), .ZN(O120));
  NANDX1 G28030 (.A1(W7914), .A2(W11795), .ZN(W16285));
  NANDX1 G28031 (.A1(I1246), .A2(W1575), .ZN(W6152));
  NANDX1 G28032 (.A1(I1267), .A2(W2281), .ZN(W6153));
  NANDX1 G28033 (.A1(W2962), .A2(W4203), .ZN(W14379));
  NANDX1 G28034 (.A1(W5000), .A2(W14790), .ZN(O1153));
  NANDX1 G28035 (.A1(W3811), .A2(W589), .ZN(W16278));
  NANDX1 G28036 (.A1(W7463), .A2(W9086), .ZN(W16277));
  NANDX1 G28037 (.A1(I1447), .A2(W1235), .ZN(W14382));
  NANDX1 G28038 (.A1(W5194), .A2(I20), .ZN(W6108));
  NANDX1 G28039 (.A1(W5605), .A2(W632), .ZN(W16273));
  NANDX1 G28040 (.A1(W9224), .A2(I716), .ZN(O1150));
  NANDX1 G28041 (.A1(W2404), .A2(W6267), .ZN(W7356));
  NANDX1 G28042 (.A1(W58), .A2(I1998), .ZN(W16268));
  NANDX1 G28043 (.A1(W246), .A2(W488), .ZN(W6168));
  NANDX1 G28044 (.A1(W419), .A2(W545), .ZN(W6169));
  NANDX1 G28045 (.A1(W4588), .A2(W1178), .ZN(W6171));
  NANDX1 G28046 (.A1(W12646), .A2(I555), .ZN(W16262));
  NANDX1 G28047 (.A1(W4947), .A2(I1281), .ZN(W6067));
  NANDX1 G28048 (.A1(I7), .A2(W7301), .ZN(W7390));
  NANDX1 G28049 (.A1(W10164), .A2(W7667), .ZN(W14316));
  NANDX1 G28050 (.A1(W10188), .A2(W13005), .ZN(W14318));
  NANDX1 G28051 (.A1(W12480), .A2(W6534), .ZN(W14322));
  NANDX1 G28052 (.A1(W2141), .A2(W6310), .ZN(W16419));
  NANDX1 G28053 (.A1(W13014), .A2(W13465), .ZN(O1175));
  NANDX1 G28054 (.A1(W4319), .A2(W4248), .ZN(W6064));
  NANDX1 G28055 (.A1(W2965), .A2(W14519), .ZN(W16416));
  NANDX1 G28056 (.A1(W2250), .A2(I264), .ZN(O179));
  NANDX1 G28057 (.A1(W14921), .A2(W14558), .ZN(W16428));
  NANDX1 G28058 (.A1(W4002), .A2(W3693), .ZN(W14334));
  NANDX1 G28059 (.A1(W12384), .A2(W13932), .ZN(W14335));
  NANDX1 G28060 (.A1(W15214), .A2(I455), .ZN(W16401));
  NANDX1 G28061 (.A1(W520), .A2(W4239), .ZN(W7381));
  NANDX1 G28062 (.A1(W1267), .A2(W733), .ZN(W7380));
  NANDX1 G28063 (.A1(W6773), .A2(I524), .ZN(W16396));
  NANDX1 G28064 (.A1(W4771), .A2(W8811), .ZN(W16395));
  NANDX1 G28065 (.A1(I470), .A2(W5317), .ZN(W6078));
  NANDX1 G28066 (.A1(W8100), .A2(W12837), .ZN(W16436));
  NANDX1 G28067 (.A1(W12485), .A2(W158), .ZN(W16452));
  NANDX1 G28068 (.A1(W12349), .A2(W11577), .ZN(W16449));
  NANDX1 G28069 (.A1(W2784), .A2(W2813), .ZN(W16448));
  NANDX1 G28070 (.A1(W376), .A2(W4509), .ZN(O1179));
  NANDX1 G28071 (.A1(W6105), .A2(W11602), .ZN(W16442));
  NANDX1 G28072 (.A1(W11969), .A2(W4577), .ZN(W14306));
  NANDX1 G28073 (.A1(W2393), .A2(I441), .ZN(W16440));
  NANDX1 G28074 (.A1(W1920), .A2(W223), .ZN(W16439));
  NANDX1 G28075 (.A1(W2403), .A2(W5414), .ZN(W16389));
  NANDX1 G28076 (.A1(W533), .A2(I113), .ZN(W6053));
  NANDX1 G28077 (.A1(W15497), .A2(W14048), .ZN(W16433));
  NANDX1 G28078 (.A1(I552), .A2(W4475), .ZN(W16432));
  NANDX1 G28079 (.A1(W4220), .A2(W5505), .ZN(W6056));
  NANDX1 G28080 (.A1(I484), .A2(W3345), .ZN(W6057));
  NANDX1 G28081 (.A1(W4893), .A2(I660), .ZN(W7391));
  NANDX1 G28082 (.A1(W1744), .A2(W5852), .ZN(W6060));
  NANDX1 G28083 (.A1(W3549), .A2(W3390), .ZN(W16429));
  NANDX1 G28084 (.A1(I890), .A2(W6812), .ZN(O1162));
  NANDX1 G28085 (.A1(W136), .A2(W724), .ZN(O1167));
  NANDX1 G28086 (.A1(W4115), .A2(W205), .ZN(W6098));
  NANDX1 G28087 (.A1(W9192), .A2(W8136), .ZN(W16362));
  NANDX1 G28088 (.A1(W2779), .A2(W5541), .ZN(W6099));
  NANDX1 G28089 (.A1(W10931), .A2(W2313), .ZN(O1166));
  NANDX1 G28090 (.A1(W5079), .A2(W5455), .ZN(W14345));
  NANDX1 G28091 (.A1(W10485), .A2(W16087), .ZN(O1165));
  NANDX1 G28092 (.A1(W6106), .A2(W2968), .ZN(W14347));
  NANDX1 G28093 (.A1(W2864), .A2(W15564), .ZN(O1168));
  NANDX1 G28094 (.A1(I636), .A2(W5561), .ZN(W6104));
  NANDX1 G28095 (.A1(W8942), .A2(W10612), .ZN(W14351));
  NANDX1 G28096 (.A1(W671), .A2(I1858), .ZN(W7374));
  NANDX1 G28097 (.A1(W9740), .A2(W7709), .ZN(O1160));
  NANDX1 G28098 (.A1(W13001), .A2(W6244), .ZN(W16345));
  NANDX1 G28099 (.A1(W3874), .A2(W14235), .ZN(W14354));
  NANDX1 G28100 (.A1(W7529), .A2(W3686), .ZN(W16343));
  NANDX1 G28101 (.A1(W3874), .A2(W2866), .ZN(W6107));
  NANDX1 G28102 (.A1(W3718), .A2(W1840), .ZN(W6086));
  NANDX1 G28103 (.A1(W2538), .A2(W3915), .ZN(W6079));
  NANDX1 G28104 (.A1(W6144), .A2(W5203), .ZN(W7376));
  NANDX1 G28105 (.A1(W13655), .A2(W6129), .ZN(W16387));
  NANDX1 G28106 (.A1(W2652), .A2(I1985), .ZN(O118));
  NANDX1 G28107 (.A1(W3177), .A2(W1223), .ZN(W6084));
  NANDX1 G28108 (.A1(W14531), .A2(W7902), .ZN(W16381));
  NANDX1 G28109 (.A1(W4793), .A2(W12866), .ZN(W16379));
  NANDX1 G28110 (.A1(W829), .A2(W2683), .ZN(W6085));
  NANDX1 G28111 (.A1(W6222), .A2(W11671), .ZN(W14389));
  NANDX1 G28112 (.A1(I647), .A2(W5722), .ZN(W6087));
  NANDX1 G28113 (.A1(W7233), .A2(W5438), .ZN(W7375));
  NANDX1 G28114 (.A1(W16295), .A2(W7866), .ZN(W16374));
  NANDX1 G28115 (.A1(W5176), .A2(W663), .ZN(W6092));
  NANDX1 G28116 (.A1(W11137), .A2(W12532), .ZN(W16372));
  NANDX1 G28117 (.A1(W4115), .A2(W115), .ZN(W6095));
  NANDX1 G28118 (.A1(W3712), .A2(W5058), .ZN(W14341));
  NANDX1 G28119 (.A1(W9297), .A2(W721), .ZN(W14342));
  NANDX1 G28120 (.A1(W992), .A2(W6827), .ZN(W16090));
  NANDX1 G28121 (.A1(W5997), .A2(W12326), .ZN(W16095));
  NANDX1 G28122 (.A1(W317), .A2(W7007), .ZN(W7311));
  NANDX1 G28123 (.A1(I1770), .A2(W1913), .ZN(W6246));
  NANDX1 G28124 (.A1(W792), .A2(W3017), .ZN(W6247));
  NANDX1 G28125 (.A1(W1516), .A2(W36), .ZN(W16094));
  NANDX1 G28126 (.A1(I546), .A2(W2463), .ZN(O869));
  NANDX1 G28127 (.A1(I1430), .A2(W4377), .ZN(W6249));
  NANDX1 G28128 (.A1(I475), .A2(W4680), .ZN(W14431));
  NANDX1 G28129 (.A1(W2112), .A2(W4838), .ZN(W14434));
  NANDX1 G28130 (.A1(W3948), .A2(W13448), .ZN(W16097));
  NANDX1 G28131 (.A1(W2741), .A2(W736), .ZN(W14435));
  NANDX1 G28132 (.A1(W9589), .A2(W8668), .ZN(W16085));
  NANDX1 G28133 (.A1(I398), .A2(W5244), .ZN(W16084));
  NANDX1 G28134 (.A1(W4592), .A2(W5059), .ZN(W7309));
  NANDX1 G28135 (.A1(W279), .A2(W5531), .ZN(W6253));
  NANDX1 G28136 (.A1(I1819), .A2(W1279), .ZN(W6254));
  NANDX1 G28137 (.A1(W2061), .A2(W5285), .ZN(W6255));
  NANDX1 G28138 (.A1(I1414), .A2(W2775), .ZN(W14438));
  NANDX1 G28139 (.A1(W8231), .A2(W4409), .ZN(O868));
  NANDX1 G28140 (.A1(I1808), .A2(W3457), .ZN(W6229));
  NANDX1 G28141 (.A1(I1504), .A2(W11582), .ZN(W14418));
  NANDX1 G28142 (.A1(W4416), .A2(I720), .ZN(W6232));
  NANDX1 G28143 (.A1(I624), .A2(W8461), .ZN(W14419));
  NANDX1 G28144 (.A1(W4633), .A2(W651), .ZN(W6234));
  NANDX1 G28145 (.A1(W4471), .A2(I1712), .ZN(W6236));
  NANDX1 G28146 (.A1(I1516), .A2(W5775), .ZN(W16109));
  NANDX1 G28147 (.A1(W783), .A2(I1134), .ZN(W6237));
  NANDX1 G28148 (.A1(I168), .A2(W14032), .ZN(O1118));
  NANDX1 G28149 (.A1(W7773), .A2(W1393), .ZN(W16108));
  NANDX1 G28150 (.A1(W3299), .A2(W1324), .ZN(W6239));
  NANDX1 G28151 (.A1(W4013), .A2(I46), .ZN(W14423));
  NANDX1 G28152 (.A1(W10555), .A2(W9144), .ZN(W14424));
  NANDX1 G28153 (.A1(W6189), .A2(W1202), .ZN(W6243));
  NANDX1 G28154 (.A1(W4943), .A2(W3249), .ZN(W14425));
  NANDX1 G28155 (.A1(W5567), .A2(W11118), .ZN(W16100));
  NANDX1 G28156 (.A1(W13556), .A2(W8547), .ZN(W14428));
  NANDX1 G28157 (.A1(W12091), .A2(W6192), .ZN(W14453));
  NANDX1 G28158 (.A1(W3953), .A2(I360), .ZN(O124));
  NANDX1 G28159 (.A1(W13816), .A2(W2667), .ZN(W16049));
  NANDX1 G28160 (.A1(W15433), .A2(W1110), .ZN(W16048));
  NANDX1 G28161 (.A1(W2996), .A2(W4523), .ZN(O175));
  NANDX1 G28162 (.A1(W3547), .A2(W2523), .ZN(W14452));
  NANDX1 G28163 (.A1(W10436), .A2(W10545), .ZN(W16046));
  NANDX1 G28164 (.A1(W13938), .A2(W14052), .ZN(O1113));
  NANDX1 G28165 (.A1(W3991), .A2(W11998), .ZN(O1112));
  NANDX1 G28166 (.A1(W4447), .A2(W14401), .ZN(W16053));
  NANDX1 G28167 (.A1(W5553), .A2(W5986), .ZN(W6274));
  NANDX1 G28168 (.A1(W273), .A2(I1322), .ZN(W6275));
  NANDX1 G28169 (.A1(I982), .A2(W8674), .ZN(W16039));
  NANDX1 G28170 (.A1(W4354), .A2(I299), .ZN(O125));
  NANDX1 G28171 (.A1(I1474), .A2(I519), .ZN(W16037));
  NANDX1 G28172 (.A1(W5272), .A2(W11620), .ZN(W16036));
  NANDX1 G28173 (.A1(W8236), .A2(W9639), .ZN(W16035));
  NANDX1 G28174 (.A1(I1685), .A2(W11794), .ZN(W16033));
  NANDX1 G28175 (.A1(W3594), .A2(W1951), .ZN(W6264));
  NANDX1 G28176 (.A1(W12253), .A2(W7611), .ZN(W14439));
  NANDX1 G28177 (.A1(W2728), .A2(W12121), .ZN(W16073));
  NANDX1 G28178 (.A1(W2687), .A2(I745), .ZN(W6256));
  NANDX1 G28179 (.A1(W737), .A2(W3610), .ZN(W6257));
  NANDX1 G28180 (.A1(W6698), .A2(I918), .ZN(W7308));
  NANDX1 G28181 (.A1(W10905), .A2(W4358), .ZN(W14444));
  NANDX1 G28182 (.A1(W10646), .A2(W13443), .ZN(W16069));
  NANDX1 G28183 (.A1(I1409), .A2(I1221), .ZN(W6261));
  NANDX1 G28184 (.A1(W14100), .A2(W7336), .ZN(W14417));
  NANDX1 G28185 (.A1(I1187), .A2(W4841), .ZN(O872));
  NANDX1 G28186 (.A1(W2546), .A2(W1437), .ZN(W6265));
  NANDX1 G28187 (.A1(W3839), .A2(W1016), .ZN(W16061));
  NANDX1 G28188 (.A1(W2519), .A2(W1220), .ZN(W7298));
  NANDX1 G28189 (.A1(W741), .A2(W7980), .ZN(W14447));
  NANDX1 G28190 (.A1(W3891), .A2(W2625), .ZN(W6269));
  NANDX1 G28191 (.A1(W3433), .A2(W343), .ZN(O1115));
  NANDX1 G28192 (.A1(W523), .A2(W6602), .ZN(W7297));
  NANDX1 G28193 (.A1(I928), .A2(W2348), .ZN(W6197));
  NANDX1 G28194 (.A1(W8079), .A2(I905), .ZN(W16205));
  NANDX1 G28195 (.A1(I782), .A2(W1941), .ZN(W6193));
  NANDX1 G28196 (.A1(W1380), .A2(W3656), .ZN(W6194));
  NANDX1 G28197 (.A1(W8863), .A2(W11838), .ZN(W16201));
  NANDX1 G28198 (.A1(I1874), .A2(W11719), .ZN(W14393));
  NANDX1 G28199 (.A1(W5898), .A2(W7920), .ZN(W16198));
  NANDX1 G28200 (.A1(W1194), .A2(W567), .ZN(W7336));
  NANDX1 G28201 (.A1(W6795), .A2(I164), .ZN(W16196));
  NANDX1 G28202 (.A1(W11821), .A2(W1391), .ZN(W14395));
  NANDX1 G28203 (.A1(W2005), .A2(I1197), .ZN(W6192));
  NANDX1 G28204 (.A1(W3214), .A2(W2808), .ZN(W6198));
  NANDX1 G28205 (.A1(W2871), .A2(W5495), .ZN(W6199));
  NANDX1 G28206 (.A1(W8784), .A2(I1112), .ZN(W16183));
  NANDX1 G28207 (.A1(W5362), .A2(W1951), .ZN(W16180));
  NANDX1 G28208 (.A1(W15532), .A2(W2054), .ZN(W16179));
  NANDX1 G28209 (.A1(I1367), .A2(W495), .ZN(W6200));
  NANDX1 G28210 (.A1(W3490), .A2(W3210), .ZN(W7329));
  NANDX1 G28211 (.A1(W1662), .A2(W2156), .ZN(W16175));
  NANDX1 G28212 (.A1(W5731), .A2(W9276), .ZN(W16221));
  NANDX1 G28213 (.A1(I1584), .A2(W5047), .ZN(W6184));
  NANDX1 G28214 (.A1(W1064), .A2(W4842), .ZN(W16231));
  NANDX1 G28215 (.A1(W5191), .A2(W10405), .ZN(O864));
  NANDX1 G28216 (.A1(W2853), .A2(W5319), .ZN(W6188));
  NANDX1 G28217 (.A1(W6573), .A2(W5059), .ZN(W7339));
  NANDX1 G28218 (.A1(W12841), .A2(W2079), .ZN(W16227));
  NANDX1 G28219 (.A1(W7219), .A2(W3272), .ZN(W16226));
  NANDX1 G28220 (.A1(W7276), .A2(W10006), .ZN(W16223));
  NANDX1 G28221 (.A1(W11525), .A2(I1064), .ZN(W16172));
  NANDX1 G28222 (.A1(I1454), .A2(I1131), .ZN(W16218));
  NANDX1 G28223 (.A1(W12693), .A2(W4479), .ZN(W16216));
  NANDX1 G28224 (.A1(W2950), .A2(W2732), .ZN(W16215));
  NANDX1 G28225 (.A1(W3432), .A2(W10081), .ZN(O1140));
  NANDX1 G28226 (.A1(I714), .A2(W287), .ZN(W6189));
  NANDX1 G28227 (.A1(W10393), .A2(W2381), .ZN(W16212));
  NANDX1 G28228 (.A1(W246), .A2(W2), .ZN(O1139));
  NANDX1 G28229 (.A1(W10277), .A2(W2202), .ZN(W14392));
  NANDX1 G28230 (.A1(W7524), .A2(W12267), .ZN(W14411));
  NANDX1 G28231 (.A1(I1333), .A2(W6143), .ZN(W16138));
  NANDX1 G28232 (.A1(W12820), .A2(W13681), .ZN(O867));
  NANDX1 G28233 (.A1(W5444), .A2(W7524), .ZN(W14409));
  NANDX1 G28234 (.A1(W13747), .A2(W8795), .ZN(O1129));
  NANDX1 G28235 (.A1(W2896), .A2(W7145), .ZN(O1128));
  NANDX1 G28236 (.A1(W3026), .A2(W2807), .ZN(W6215));
  NANDX1 G28237 (.A1(W5611), .A2(W3821), .ZN(W6217));
  NANDX1 G28238 (.A1(I1326), .A2(W13380), .ZN(W16131));
  NANDX1 G28239 (.A1(W11645), .A2(W8980), .ZN(W16139));
  NANDX1 G28240 (.A1(I1639), .A2(W303), .ZN(W6221));
  NANDX1 G28241 (.A1(I396), .A2(W2566), .ZN(W7317));
  NANDX1 G28242 (.A1(W4578), .A2(W38), .ZN(W6222));
  NANDX1 G28243 (.A1(I197), .A2(W3282), .ZN(W6223));
  NANDX1 G28244 (.A1(W5297), .A2(W2409), .ZN(W6225));
  NANDX1 G28245 (.A1(W1864), .A2(W138), .ZN(W6226));
  NANDX1 G28246 (.A1(W2272), .A2(W4474), .ZN(W7315));
  NANDX1 G28247 (.A1(W1396), .A2(W11768), .ZN(W14416));
  NANDX1 G28248 (.A1(I410), .A2(W5175), .ZN(W6205));
  NANDX1 G28249 (.A1(W11794), .A2(I866), .ZN(W16171));
  NANDX1 G28250 (.A1(W1787), .A2(W1505), .ZN(W7325));
  NANDX1 G28251 (.A1(W11814), .A2(W15963), .ZN(W16160));
  NANDX1 G28252 (.A1(W9993), .A2(W5886), .ZN(W16156));
  NANDX1 G28253 (.A1(W7538), .A2(W14215), .ZN(W14407));
  NANDX1 G28254 (.A1(W5872), .A2(I1263), .ZN(W16151));
  NANDX1 G28255 (.A1(W1601), .A2(I232), .ZN(W16150));
  NANDX1 G28256 (.A1(W45), .A2(I1744), .ZN(W6204));
  NANDX1 G28257 (.A1(W1660), .A2(W6365), .ZN(W14610));
  NANDX1 G28258 (.A1(I1464), .A2(W5622), .ZN(W6206));
  NANDX1 G28259 (.A1(W2176), .A2(W4970), .ZN(W6208));
  NANDX1 G28260 (.A1(W11763), .A2(W12584), .ZN(W16147));
  NANDX1 G28261 (.A1(W13749), .A2(W6834), .ZN(W16144));
  NANDX1 G28262 (.A1(W13758), .A2(I144), .ZN(O1130));
  NANDX1 G28263 (.A1(W2385), .A2(W2890), .ZN(W6209));
  NANDX1 G28264 (.A1(I1906), .A2(W11541), .ZN(W16142));
  NANDX1 G28265 (.A1(W12849), .A2(I915), .ZN(W16141));
  NANDX1 G28266 (.A1(W8302), .A2(W6926), .ZN(W14819));
  NANDX1 G28267 (.A1(W8146), .A2(W12793), .ZN(W15167));
  NANDX1 G28268 (.A1(W3983), .A2(W5243), .ZN(W6830));
  NANDX1 G28269 (.A1(I474), .A2(W121), .ZN(W15166));
  NANDX1 G28270 (.A1(W2542), .A2(I1839), .ZN(W15164));
  NANDX1 G28271 (.A1(W3741), .A2(I432), .ZN(W15163));
  NANDX1 G28272 (.A1(W3371), .A2(W5139), .ZN(W6831));
  NANDX1 G28273 (.A1(W2811), .A2(W8453), .ZN(O970));
  NANDX1 G28274 (.A1(W5678), .A2(W9673), .ZN(W15157));
  NANDX1 G28275 (.A1(W830), .A2(W4309), .ZN(W7034));
  NANDX1 G28276 (.A1(W1807), .A2(I71), .ZN(W6829));
  NANDX1 G28277 (.A1(W9900), .A2(W7153), .ZN(W15154));
  NANDX1 G28278 (.A1(I1578), .A2(W8182), .ZN(W15153));
  NANDX1 G28279 (.A1(W14439), .A2(I272), .ZN(W15152));
  NANDX1 G28280 (.A1(I1846), .A2(I331), .ZN(W6834));
  NANDX1 G28281 (.A1(W10746), .A2(W54), .ZN(W14821));
  NANDX1 G28282 (.A1(W6435), .A2(I1901), .ZN(W7028));
  NANDX1 G28283 (.A1(W9865), .A2(W4278), .ZN(W14822));
  NANDX1 G28284 (.A1(W12296), .A2(I1602), .ZN(O923));
  NANDX1 G28285 (.A1(W5954), .A2(W11327), .ZN(W15184));
  NANDX1 G28286 (.A1(W5828), .A2(W4290), .ZN(W6814));
  NANDX1 G28287 (.A1(W125), .A2(W1627), .ZN(W6816));
  NANDX1 G28288 (.A1(W1035), .A2(I1130), .ZN(W6818));
  NANDX1 G28289 (.A1(W3978), .A2(W13379), .ZN(W14810));
  NANDX1 G28290 (.A1(W6699), .A2(W4471), .ZN(W7043));
  NANDX1 G28291 (.A1(W405), .A2(W5677), .ZN(W7042));
  NANDX1 G28292 (.A1(W6021), .A2(W3361), .ZN(W6824));
  NANDX1 G28293 (.A1(W483), .A2(W8522), .ZN(O920));
  NANDX1 G28294 (.A1(W6035), .A2(W3491), .ZN(W6841));
  NANDX1 G28295 (.A1(I901), .A2(W54), .ZN(W6825));
  NANDX1 G28296 (.A1(W2314), .A2(W2338), .ZN(O162));
  NANDX1 G28297 (.A1(W3647), .A2(W2125), .ZN(W15179));
  NANDX1 G28298 (.A1(W6134), .A2(W9330), .ZN(O972));
  NANDX1 G28299 (.A1(W14825), .A2(W197), .ZN(W15176));
  NANDX1 G28300 (.A1(W3019), .A2(I1609), .ZN(O971));
  NANDX1 G28301 (.A1(W6546), .A2(W1522), .ZN(W15171));
  NANDX1 G28302 (.A1(W6048), .A2(W4089), .ZN(W15170));
  NANDX1 G28303 (.A1(I537), .A2(W1919), .ZN(W14839));
  NANDX1 G28304 (.A1(W14075), .A2(W12795), .ZN(W15120));
  NANDX1 G28305 (.A1(W5517), .A2(I884), .ZN(W6856));
  NANDX1 G28306 (.A1(W9049), .A2(W913), .ZN(W14837));
  NANDX1 G28307 (.A1(W6701), .A2(W14027), .ZN(W15118));
  NANDX1 G28308 (.A1(W4071), .A2(W297), .ZN(W15117));
  NANDX1 G28309 (.A1(I535), .A2(W71), .ZN(W6859));
  NANDX1 G28310 (.A1(W1663), .A2(W12500), .ZN(O962));
  NANDX1 G28311 (.A1(W4842), .A2(W956), .ZN(W7024));
  NANDX1 G28312 (.A1(W8679), .A2(W3796), .ZN(O964));
  NANDX1 G28313 (.A1(W5962), .A2(W1920), .ZN(W7022));
  NANDX1 G28314 (.A1(W6587), .A2(I1209), .ZN(W6861));
  NANDX1 G28315 (.A1(W1160), .A2(W2338), .ZN(W6862));
  NANDX1 G28316 (.A1(W1443), .A2(W5625), .ZN(W15104));
  NANDX1 G28317 (.A1(I1639), .A2(I1883), .ZN(W6864));
  NANDX1 G28318 (.A1(W59), .A2(W5960), .ZN(W6866));
  NANDX1 G28319 (.A1(W1090), .A2(W5508), .ZN(W14840));
  NANDX1 G28320 (.A1(W1169), .A2(I714), .ZN(W6868));
  NANDX1 G28321 (.A1(W2201), .A2(W1834), .ZN(W6844));
  NANDX1 G28322 (.A1(I1412), .A2(W13437), .ZN(W15144));
  NANDX1 G28323 (.A1(W2489), .A2(W6165), .ZN(W6843));
  NANDX1 G28324 (.A1(W8561), .A2(W10880), .ZN(W15139));
  NANDX1 G28325 (.A1(W3856), .A2(W7701), .ZN(O967));
  NANDX1 G28326 (.A1(W6524), .A2(W6118), .ZN(O966));
  NANDX1 G28327 (.A1(W1893), .A2(W7009), .ZN(W7027));
  NANDX1 G28328 (.A1(W10225), .A2(W3639), .ZN(W14828));
  NANDX1 G28329 (.A1(W8312), .A2(W6081), .ZN(W15134));
  NANDX1 G28330 (.A1(W793), .A2(I310), .ZN(W6813));
  NANDX1 G28331 (.A1(W5749), .A2(W150), .ZN(W14830));
  NANDX1 G28332 (.A1(W10316), .A2(W9360), .ZN(W14832));
  NANDX1 G28333 (.A1(I1974), .A2(W5827), .ZN(W7026));
  NANDX1 G28334 (.A1(W3637), .A2(I446), .ZN(W6852));
  NANDX1 G28335 (.A1(W203), .A2(W2948), .ZN(W15129));
  NANDX1 G28336 (.A1(W14779), .A2(W3557), .ZN(W15127));
  NANDX1 G28337 (.A1(W3908), .A2(W6023), .ZN(O153));
  NANDX1 G28338 (.A1(W3649), .A2(W10946), .ZN(W15124));
  NANDX1 G28339 (.A1(W11728), .A2(W665), .ZN(W14787));
  NANDX1 G28340 (.A1(W8382), .A2(W6467), .ZN(W14782));
  NANDX1 G28341 (.A1(I704), .A2(I1150), .ZN(W6763));
  NANDX1 G28342 (.A1(W4462), .A2(W3300), .ZN(W6766));
  NANDX1 G28343 (.A1(W745), .A2(W5761), .ZN(W6767));
  NANDX1 G28344 (.A1(W1058), .A2(W4228), .ZN(O981));
  NANDX1 G28345 (.A1(W13629), .A2(W1620), .ZN(W15252));
  NANDX1 G28346 (.A1(W13), .A2(W3558), .ZN(W6768));
  NANDX1 G28347 (.A1(W12082), .A2(W11852), .ZN(W14784));
  NANDX1 G28348 (.A1(W575), .A2(W14403), .ZN(W14786));
  NANDX1 G28349 (.A1(I1308), .A2(W1608), .ZN(W7068));
  NANDX1 G28350 (.A1(I96), .A2(W3679), .ZN(W6775));
  NANDX1 G28351 (.A1(I200), .A2(W8313), .ZN(O977));
  NANDX1 G28352 (.A1(W12256), .A2(W10745), .ZN(W15243));
  NANDX1 G28353 (.A1(W7284), .A2(W9383), .ZN(W15242));
  NANDX1 G28354 (.A1(W6667), .A2(W5336), .ZN(O976));
  NANDX1 G28355 (.A1(I702), .A2(W5450), .ZN(W14790));
  NANDX1 G28356 (.A1(W2721), .A2(W5362), .ZN(W6781));
  NANDX1 G28357 (.A1(W1472), .A2(W12666), .ZN(O916));
  NANDX1 G28358 (.A1(W14839), .A2(W3681), .ZN(W15266));
  NANDX1 G28359 (.A1(W12188), .A2(W4846), .ZN(W15273));
  NANDX1 G28360 (.A1(W7540), .A2(W3318), .ZN(W14768));
  NANDX1 G28361 (.A1(W5061), .A2(W1736), .ZN(W15272));
  NANDX1 G28362 (.A1(W1395), .A2(W5667), .ZN(W7071));
  NANDX1 G28363 (.A1(W8136), .A2(I1255), .ZN(W15271));
  NANDX1 G28364 (.A1(W15031), .A2(W3317), .ZN(W15270));
  NANDX1 G28365 (.A1(I137), .A2(I1276), .ZN(W15269));
  NANDX1 G28366 (.A1(W3520), .A2(W6673), .ZN(W14770));
  NANDX1 G28367 (.A1(W6681), .A2(W1345), .ZN(W6785));
  NANDX1 G28368 (.A1(W10978), .A2(W5117), .ZN(W14774));
  NANDX1 G28369 (.A1(W14161), .A2(I958), .ZN(W14776));
  NANDX1 G28370 (.A1(W8279), .A2(W14989), .ZN(W15264));
  NANDX1 G28371 (.A1(W4022), .A2(W7512), .ZN(W15263));
  NANDX1 G28372 (.A1(W3913), .A2(W1058), .ZN(W6757));
  NANDX1 G28373 (.A1(W10894), .A2(W6507), .ZN(W15261));
  NANDX1 G28374 (.A1(W6014), .A2(W6702), .ZN(W7070));
  NANDX1 G28375 (.A1(W3259), .A2(I1671), .ZN(W15259));
  NANDX1 G28376 (.A1(W1474), .A2(W4231), .ZN(W14805));
  NANDX1 G28377 (.A1(I1690), .A2(W2551), .ZN(W7051));
  NANDX1 G28378 (.A1(W7292), .A2(W13875), .ZN(W15210));
  NANDX1 G28379 (.A1(W5505), .A2(W8814), .ZN(W15209));
  NANDX1 G28380 (.A1(W3401), .A2(W1052), .ZN(O152));
  NANDX1 G28381 (.A1(W465), .A2(W5622), .ZN(W15206));
  NANDX1 G28382 (.A1(W446), .A2(W7499), .ZN(W15203));
  NANDX1 G28383 (.A1(W716), .A2(W219), .ZN(W6802));
  NANDX1 G28384 (.A1(W5522), .A2(W2675), .ZN(W6803));
  NANDX1 G28385 (.A1(W1214), .A2(W13999), .ZN(W15215));
  NANDX1 G28386 (.A1(W13638), .A2(W5373), .ZN(W14806));
  NANDX1 G28387 (.A1(W1715), .A2(W2145), .ZN(W7047));
  NANDX1 G28388 (.A1(W606), .A2(W9991), .ZN(W15200));
  NANDX1 G28389 (.A1(W4217), .A2(W1342), .ZN(W6809));
  NANDX1 G28390 (.A1(I1104), .A2(W13951), .ZN(W15196));
  NANDX1 G28391 (.A1(W7952), .A2(I476), .ZN(W15195));
  NANDX1 G28392 (.A1(W2726), .A2(W14353), .ZN(W15194));
  NANDX1 G28393 (.A1(W1340), .A2(W1651), .ZN(W15193));
  NANDX1 G28394 (.A1(W7574), .A2(W2327), .ZN(W15226));
  NANDX1 G28395 (.A1(W5107), .A2(W3369), .ZN(W14793));
  NANDX1 G28396 (.A1(W4464), .A2(I1338), .ZN(W7060));
  NANDX1 G28397 (.A1(W5507), .A2(I764), .ZN(W6789));
  NANDX1 G28398 (.A1(W5380), .A2(W1771), .ZN(W15233));
  NANDX1 G28399 (.A1(W4822), .A2(W5442), .ZN(W14796));
  NANDX1 G28400 (.A1(W3794), .A2(W1358), .ZN(W15228));
  NANDX1 G28401 (.A1(W4704), .A2(I887), .ZN(W6792));
  NANDX1 G28402 (.A1(W10272), .A2(W2697), .ZN(W15227));
  NANDX1 G28403 (.A1(I1100), .A2(W4848), .ZN(W6869));
  NANDX1 G28404 (.A1(I662), .A2(W7422), .ZN(W15224));
  NANDX1 G28405 (.A1(I697), .A2(W9167), .ZN(O975));
  NANDX1 G28406 (.A1(W9051), .A2(W6627), .ZN(W15220));
  NANDX1 G28407 (.A1(I849), .A2(W1277), .ZN(W6796));
  NANDX1 G28408 (.A1(I1411), .A2(W5593), .ZN(W7054));
  NANDX1 G28409 (.A1(I1586), .A2(W1299), .ZN(W15218));
  NANDX1 G28410 (.A1(I1865), .A2(I1306), .ZN(W6798));
  NANDX1 G28411 (.A1(W1674), .A2(W4744), .ZN(W7053));
  NANDX1 G28412 (.A1(W10940), .A2(W82), .ZN(W14950));
  NANDX1 G28413 (.A1(W115), .A2(W584), .ZN(W6953));
  NANDX1 G28414 (.A1(W11670), .A2(W7575), .ZN(W14960));
  NANDX1 G28415 (.A1(W1452), .A2(I1909), .ZN(W14959));
  NANDX1 G28416 (.A1(W6200), .A2(I1448), .ZN(W6954));
  NANDX1 G28417 (.A1(W9855), .A2(I687), .ZN(O929));
  NANDX1 G28418 (.A1(W14464), .A2(W6487), .ZN(W14954));
  NANDX1 G28419 (.A1(W3373), .A2(W6199), .ZN(W14953));
  NANDX1 G28420 (.A1(W7476), .A2(I422), .ZN(W14887));
  NANDX1 G28421 (.A1(W3016), .A2(W6698), .ZN(W6991));
  NANDX1 G28422 (.A1(W3330), .A2(W5138), .ZN(W14962));
  NANDX1 G28423 (.A1(I723), .A2(W4727), .ZN(W6957));
  NANDX1 G28424 (.A1(W11820), .A2(I445), .ZN(W14889));
  NANDX1 G28425 (.A1(W6102), .A2(W8028), .ZN(W14949));
  NANDX1 G28426 (.A1(W13254), .A2(W3540), .ZN(O935));
  NANDX1 G28427 (.A1(W178), .A2(W9855), .ZN(W14947));
  NANDX1 G28428 (.A1(I248), .A2(W3116), .ZN(W6989));
  NANDX1 G28429 (.A1(W8727), .A2(W4672), .ZN(W14891));
  NANDX1 G28430 (.A1(W4848), .A2(W14543), .ZN(O934));
  NANDX1 G28431 (.A1(W9201), .A2(W13689), .ZN(O940));
  NANDX1 G28432 (.A1(W654), .A2(W229), .ZN(W6938));
  NANDX1 G28433 (.A1(W1007), .A2(W11600), .ZN(W14984));
  NANDX1 G28434 (.A1(W5728), .A2(W474), .ZN(W6940));
  NANDX1 G28435 (.A1(W1790), .A2(W8767), .ZN(W14876));
  NANDX1 G28436 (.A1(W11341), .A2(W2668), .ZN(W14982));
  NANDX1 G28437 (.A1(W3918), .A2(W2844), .ZN(O157));
  NANDX1 G28438 (.A1(W138), .A2(W499), .ZN(W6948));
  NANDX1 G28439 (.A1(I1255), .A2(W2266), .ZN(W6949));
  NANDX1 G28440 (.A1(W1601), .A2(W14641), .ZN(W14940));
  NANDX1 G28441 (.A1(I444), .A2(W4869), .ZN(W14973));
  NANDX1 G28442 (.A1(W10419), .A2(W5283), .ZN(W14972));
  NANDX1 G28443 (.A1(W2882), .A2(W5028), .ZN(W14969));
  NANDX1 G28444 (.A1(W2481), .A2(W6676), .ZN(W6995));
  NANDX1 G28445 (.A1(I200), .A2(W3832), .ZN(W14968));
  NANDX1 G28446 (.A1(W12599), .A2(W6286), .ZN(W14966));
  NANDX1 G28447 (.A1(W14064), .A2(I1148), .ZN(W14883));
  NANDX1 G28448 (.A1(W4140), .A2(W3098), .ZN(W6952));
  NANDX1 G28449 (.A1(W1525), .A2(W4845), .ZN(W6985));
  NANDX1 G28450 (.A1(W4424), .A2(W18), .ZN(W14921));
  NANDX1 G28451 (.A1(W3323), .A2(W1524), .ZN(W14920));
  NANDX1 G28452 (.A1(W397), .A2(W1530), .ZN(W6975));
  NANDX1 G28453 (.A1(W1647), .A2(W14194), .ZN(W14899));
  NANDX1 G28454 (.A1(W4385), .A2(W2650), .ZN(W6979));
  NANDX1 G28455 (.A1(W4066), .A2(W165), .ZN(W6980));
  NANDX1 G28456 (.A1(W12334), .A2(W627), .ZN(W14916));
  NANDX1 G28457 (.A1(I1032), .A2(W5818), .ZN(W6981));
  NANDX1 G28458 (.A1(W3480), .A2(W1568), .ZN(W6973));
  NANDX1 G28459 (.A1(W12965), .A2(W344), .ZN(O931));
  NANDX1 G28460 (.A1(W9768), .A2(W11193), .ZN(W14902));
  NANDX1 G28461 (.A1(W14883), .A2(I1293), .ZN(W14906));
  NANDX1 G28462 (.A1(W2332), .A2(W6826), .ZN(W6982));
  NANDX1 G28463 (.A1(W620), .A2(I285), .ZN(W6983));
  NANDX1 G28464 (.A1(W2845), .A2(W5826), .ZN(W6984));
  NANDX1 G28465 (.A1(W11711), .A2(W9008), .ZN(W14903));
  NANDX1 G28466 (.A1(W9485), .A2(W13153), .ZN(W14904));
  NANDX1 G28467 (.A1(W1441), .A2(W5878), .ZN(W14894));
  NANDX1 G28468 (.A1(W3113), .A2(W6022), .ZN(W14939));
  NANDX1 G28469 (.A1(W4547), .A2(W6523), .ZN(W6958));
  NANDX1 G28470 (.A1(W12920), .A2(W13298), .ZN(W14937));
  NANDX1 G28471 (.A1(W10244), .A2(W2555), .ZN(W14892));
  NANDX1 G28472 (.A1(W8575), .A2(W4668), .ZN(W14936));
  NANDX1 G28473 (.A1(W12016), .A2(W5978), .ZN(W14893));
  NANDX1 G28474 (.A1(W3984), .A2(I413), .ZN(W6961));
  NANDX1 G28475 (.A1(W5838), .A2(W5674), .ZN(W6962));
  NANDX1 G28476 (.A1(W6594), .A2(W1153), .ZN(W14989));
  NANDX1 G28477 (.A1(W1557), .A2(W12850), .ZN(W14895));
  NANDX1 G28478 (.A1(W5750), .A2(W617), .ZN(W6964));
  NANDX1 G28479 (.A1(W2910), .A2(I791), .ZN(W14896));
  NANDX1 G28480 (.A1(W1505), .A2(W6267), .ZN(W14933));
  NANDX1 G28481 (.A1(W14474), .A2(W10916), .ZN(W14926));
  NANDX1 G28482 (.A1(W3679), .A2(W3371), .ZN(W6988));
  NANDX1 G28483 (.A1(W7305), .A2(W2147), .ZN(W14898));
  NANDX1 G28484 (.A1(W4910), .A2(W6617), .ZN(W14923));
  NANDX1 G28485 (.A1(W1801), .A2(W5132), .ZN(W6894));
  NANDX1 G28486 (.A1(W11716), .A2(W10171), .ZN(W15071));
  NANDX1 G28487 (.A1(W10267), .A2(W2753), .ZN(W14843));
  NANDX1 G28488 (.A1(W1749), .A2(W589), .ZN(W14848));
  NANDX1 G28489 (.A1(W3714), .A2(I701), .ZN(W6889));
  NANDX1 G28490 (.A1(W727), .A2(W1685), .ZN(W14850));
  NANDX1 G28491 (.A1(W1006), .A2(W4346), .ZN(W6890));
  NANDX1 G28492 (.A1(W6081), .A2(W3370), .ZN(W7014));
  NANDX1 G28493 (.A1(W228), .A2(I1432), .ZN(W6891));
  NANDX1 G28494 (.A1(I670), .A2(W3957), .ZN(W6893));
  NANDX1 G28495 (.A1(W5705), .A2(W6081), .ZN(W6886));
  NANDX1 G28496 (.A1(I1629), .A2(W9731), .ZN(W14855));
  NANDX1 G28497 (.A1(I225), .A2(W541), .ZN(W6897));
  NANDX1 G28498 (.A1(W869), .A2(W9868), .ZN(O954));
  NANDX1 G28499 (.A1(W14924), .A2(W482), .ZN(W15049));
  NANDX1 G28500 (.A1(W113), .A2(W12376), .ZN(W15046));
  NANDX1 G28501 (.A1(I754), .A2(W5853), .ZN(W15045));
  NANDX1 G28502 (.A1(W3260), .A2(I913), .ZN(W6903));
  NANDX1 G28503 (.A1(W1433), .A2(W6499), .ZN(W6905));
  NANDX1 G28504 (.A1(W10198), .A2(W1316), .ZN(W15083));
  NANDX1 G28505 (.A1(W4677), .A2(W6678), .ZN(W6870));
  NANDX1 G28506 (.A1(W11294), .A2(W9933), .ZN(W15094));
  NANDX1 G28507 (.A1(W3796), .A2(W6082), .ZN(W15092));
  NANDX1 G28508 (.A1(I458), .A2(W8294), .ZN(W15090));
  NANDX1 G28509 (.A1(W10664), .A2(W13583), .ZN(W15089));
  NANDX1 G28510 (.A1(W1913), .A2(W14029), .ZN(O959));
  NANDX1 G28511 (.A1(W3346), .A2(W1011), .ZN(W7019));
  NANDX1 G28512 (.A1(W5476), .A2(W2577), .ZN(W6873));
  NANDX1 G28513 (.A1(W7404), .A2(I1886), .ZN(W15040));
  NANDX1 G28514 (.A1(W3729), .A2(W8828), .ZN(W14841));
  NANDX1 G28515 (.A1(W4461), .A2(W234), .ZN(W6878));
  NANDX1 G28516 (.A1(W6410), .A2(W7695), .ZN(W15080));
  NANDX1 G28517 (.A1(W1771), .A2(W6139), .ZN(W6879));
  NANDX1 G28518 (.A1(W8184), .A2(W6595), .ZN(O958));
  NANDX1 G28519 (.A1(W3389), .A2(W1690), .ZN(W6881));
  NANDX1 G28520 (.A1(W191), .A2(W4698), .ZN(W6882));
  NANDX1 G28521 (.A1(W2861), .A2(W5749), .ZN(W7017));
  NANDX1 G28522 (.A1(W6760), .A2(W9075), .ZN(W14868));
  NANDX1 G28523 (.A1(W5236), .A2(W14237), .ZN(W15016));
  NANDX1 G28524 (.A1(W7428), .A2(W4139), .ZN(W15014));
  NANDX1 G28525 (.A1(W1104), .A2(W5868), .ZN(W7003));
  NANDX1 G28526 (.A1(W11320), .A2(W13286), .ZN(O943));
  NANDX1 G28527 (.A1(W3860), .A2(W50), .ZN(W6927));
  NANDX1 G28528 (.A1(W12290), .A2(W13599), .ZN(W15004));
  NANDX1 G28529 (.A1(W941), .A2(I814), .ZN(W6930));
  NANDX1 G28530 (.A1(W1973), .A2(W10459), .ZN(W14998));
  NANDX1 G28531 (.A1(W8720), .A2(W6270), .ZN(W15019));
  NANDX1 G28532 (.A1(W6951), .A2(W9210), .ZN(W14996));
  NANDX1 G28533 (.A1(W6400), .A2(W6122), .ZN(W14995));
  NANDX1 G28534 (.A1(W11355), .A2(W5817), .ZN(W14994));
  NANDX1 G28535 (.A1(W13106), .A2(W7497), .ZN(W14871));
  NANDX1 G28536 (.A1(I878), .A2(W11205), .ZN(W14874));
  NANDX1 G28537 (.A1(W9987), .A2(W6464), .ZN(W14991));
  NANDX1 G28538 (.A1(W12775), .A2(W13295), .ZN(W14990));
  NANDX1 G28539 (.A1(W6847), .A2(I720), .ZN(W6935));
  NANDX1 G28540 (.A1(W6162), .A2(W2234), .ZN(W15027));
  NANDX1 G28541 (.A1(W8448), .A2(W8591), .ZN(W14856));
  NANDX1 G28542 (.A1(W1928), .A2(W341), .ZN(W15039));
  NANDX1 G28543 (.A1(W8992), .A2(W2066), .ZN(W14857));
  NANDX1 G28544 (.A1(W4902), .A2(W2186), .ZN(W7008));
  NANDX1 G28545 (.A1(I6), .A2(W13721), .ZN(O950));
  NANDX1 G28546 (.A1(W392), .A2(I166), .ZN(W6907));
  NANDX1 G28547 (.A1(W5331), .A2(W7902), .ZN(W14858));
  NANDX1 G28548 (.A1(I1314), .A2(W6155), .ZN(W6911));
  NANDX1 G28549 (.A1(I1939), .A2(I1220), .ZN(W7073));
  NANDX1 G28550 (.A1(W371), .A2(W6172), .ZN(W6912));
  NANDX1 G28551 (.A1(W6577), .A2(W3630), .ZN(W7007));
  NANDX1 G28552 (.A1(W5217), .A2(W803), .ZN(W6915));
  NANDX1 G28553 (.A1(W5654), .A2(W5128), .ZN(W14860));
  NANDX1 G28554 (.A1(W1553), .A2(W984), .ZN(W6920));
  NANDX1 G28555 (.A1(W1381), .A2(W859), .ZN(W7005));
  NANDX1 G28556 (.A1(W7481), .A2(W11317), .ZN(O945));
  NANDX1 G28557 (.A1(W10050), .A2(W1653), .ZN(O944));
  NANDX1 G28558 (.A1(W9190), .A2(W3339), .ZN(W15538));
  NANDX1 G28559 (.A1(W761), .A2(W2362), .ZN(W15551));
  NANDX1 G28560 (.A1(I917), .A2(W2153), .ZN(W15549));
  NANDX1 G28561 (.A1(W2872), .A2(W6366), .ZN(W6606));
  NANDX1 G28562 (.A1(W3345), .A2(W13050), .ZN(W15545));
  NANDX1 G28563 (.A1(W1097), .A2(W9842), .ZN(W15544));
  NANDX1 G28564 (.A1(W13602), .A2(W11792), .ZN(W14652));
  NANDX1 G28565 (.A1(W11289), .A2(W3036), .ZN(W15542));
  NANDX1 G28566 (.A1(W580), .A2(W14558), .ZN(W14654));
  NANDX1 G28567 (.A1(W1735), .A2(W9010), .ZN(O1026));
  NANDX1 G28568 (.A1(W3148), .A2(W3772), .ZN(O1027));
  NANDX1 G28569 (.A1(W6870), .A2(W14545), .ZN(W15536));
  NANDX1 G28570 (.A1(W2642), .A2(I135), .ZN(O1024));
  NANDX1 G28571 (.A1(W8273), .A2(W12855), .ZN(W15533));
  NANDX1 G28572 (.A1(I1053), .A2(I1956), .ZN(W7169));
  NANDX1 G28573 (.A1(W12771), .A2(W3900), .ZN(W15528));
  NANDX1 G28574 (.A1(W6267), .A2(I1346), .ZN(W15527));
  NANDX1 G28575 (.A1(W6672), .A2(W2665), .ZN(W15526));
  NANDX1 G28576 (.A1(W2927), .A2(W3699), .ZN(W7168));
  NANDX1 G28577 (.A1(W5516), .A2(I1186), .ZN(W14639));
  NANDX1 G28578 (.A1(W475), .A2(W3974), .ZN(W6590));
  NANDX1 G28579 (.A1(W6010), .A2(I1294), .ZN(W7175));
  NANDX1 G28580 (.A1(W13740), .A2(W1952), .ZN(W15567));
  NANDX1 G28581 (.A1(W3779), .A2(W3666), .ZN(W15566));
  NANDX1 G28582 (.A1(W1107), .A2(W7237), .ZN(W15565));
  NANDX1 G28583 (.A1(W2049), .A2(W8271), .ZN(W15564));
  NANDX1 G28584 (.A1(W4310), .A2(W1327), .ZN(W6595));
  NANDX1 G28585 (.A1(W3973), .A2(W14424), .ZN(W15563));
  NANDX1 G28586 (.A1(W8975), .A2(W1755), .ZN(W14662));
  NANDX1 G28587 (.A1(W11538), .A2(W7229), .ZN(W14640));
  NANDX1 G28588 (.A1(W1622), .A2(W12555), .ZN(W15561));
  NANDX1 G28589 (.A1(I1392), .A2(W6925), .ZN(W15560));
  NANDX1 G28590 (.A1(I126), .A2(W2943), .ZN(W6597));
  NANDX1 G28591 (.A1(W1833), .A2(W6299), .ZN(W15559));
  NANDX1 G28592 (.A1(W8782), .A2(W12424), .ZN(W14642));
  NANDX1 G28593 (.A1(I1816), .A2(W5764), .ZN(W6600));
  NANDX1 G28594 (.A1(W5822), .A2(W4637), .ZN(W15554));
  NANDX1 G28595 (.A1(W10040), .A2(W8810), .ZN(W14677));
  NANDX1 G28596 (.A1(W1420), .A2(W6611), .ZN(W6625));
  NANDX1 G28597 (.A1(W6230), .A2(W5761), .ZN(W6627));
  NANDX1 G28598 (.A1(W584), .A2(W1850), .ZN(W14670));
  NANDX1 G28599 (.A1(W13225), .A2(W11300), .ZN(W14672));
  NANDX1 G28600 (.A1(W4350), .A2(W6408), .ZN(W7163));
  NANDX1 G28601 (.A1(I1718), .A2(W10291), .ZN(W15488));
  NANDX1 G28602 (.A1(W3789), .A2(W2276), .ZN(O139));
  NANDX1 G28603 (.A1(W5211), .A2(W282), .ZN(W15487));
  NANDX1 G28604 (.A1(W2442), .A2(W4408), .ZN(W15495));
  NANDX1 G28605 (.A1(W2368), .A2(W14361), .ZN(W15485));
  NANDX1 G28606 (.A1(W11358), .A2(W9268), .ZN(W14678));
  NANDX1 G28607 (.A1(W4954), .A2(W5164), .ZN(W6640));
  NANDX1 G28608 (.A1(I502), .A2(I32), .ZN(W7158));
  NANDX1 G28609 (.A1(W6476), .A2(W7964), .ZN(W14679));
  NANDX1 G28610 (.A1(W6432), .A2(W6737), .ZN(W7156));
  NANDX1 G28611 (.A1(I1495), .A2(I597), .ZN(W6641));
  NANDX1 G28612 (.A1(W7679), .A2(W689), .ZN(W15479));
  NANDX1 G28613 (.A1(W1009), .A2(W788), .ZN(W15516));
  NANDX1 G28614 (.A1(I825), .A2(W11748), .ZN(W15524));
  NANDX1 G28615 (.A1(W14238), .A2(W13407), .ZN(W14663));
  NANDX1 G28616 (.A1(I1377), .A2(W825), .ZN(W7167));
  NANDX1 G28617 (.A1(W2521), .A2(W929), .ZN(W14667));
  NANDX1 G28618 (.A1(W2270), .A2(W5873), .ZN(W6617));
  NANDX1 G28619 (.A1(I537), .A2(W4370), .ZN(O1021));
  NANDX1 G28620 (.A1(W4482), .A2(I1694), .ZN(W6619));
  NANDX1 G28621 (.A1(W12874), .A2(W7503), .ZN(W15517));
  NANDX1 G28622 (.A1(W8328), .A2(W135), .ZN(W15569));
  NANDX1 G28623 (.A1(W12206), .A2(W47), .ZN(W15513));
  NANDX1 G28624 (.A1(W1124), .A2(W6397), .ZN(W15508));
  NANDX1 G28625 (.A1(W9491), .A2(I1656), .ZN(W15507));
  NANDX1 G28626 (.A1(W3928), .A2(I549), .ZN(W15504));
  NANDX1 G28627 (.A1(W5615), .A2(I358), .ZN(W6621));
  NANDX1 G28628 (.A1(W11128), .A2(I72), .ZN(W15501));
  NANDX1 G28629 (.A1(W5545), .A2(W5413), .ZN(W6624));
  NANDX1 G28630 (.A1(W11780), .A2(W238), .ZN(W15497));
  NANDX1 G28631 (.A1(W7889), .A2(W5555), .ZN(W15633));
  NANDX1 G28632 (.A1(W160), .A2(W13134), .ZN(W14620));
  NANDX1 G28633 (.A1(W9122), .A2(W10100), .ZN(W15641));
  NANDX1 G28634 (.A1(W4608), .A2(I531), .ZN(W6553));
  NANDX1 G28635 (.A1(W205), .A2(W1297), .ZN(W15639));
  NANDX1 G28636 (.A1(W10828), .A2(W12142), .ZN(W15638));
  NANDX1 G28637 (.A1(I1088), .A2(W2817), .ZN(W6556));
  NANDX1 G28638 (.A1(W3239), .A2(I1550), .ZN(W6558));
  NANDX1 G28639 (.A1(I1720), .A2(W5717), .ZN(W6561));
  NANDX1 G28640 (.A1(W3667), .A2(W8401), .ZN(W15634));
  NANDX1 G28641 (.A1(I1264), .A2(W15631), .ZN(W15644));
  NANDX1 G28642 (.A1(W2195), .A2(W5030), .ZN(W15632));
  NANDX1 G28643 (.A1(W1712), .A2(W14163), .ZN(W15630));
  NANDX1 G28644 (.A1(W5779), .A2(W3776), .ZN(O1041));
  NANDX1 G28645 (.A1(W343), .A2(I198), .ZN(O169));
  NANDX1 G28646 (.A1(W6038), .A2(W3939), .ZN(W15628));
  NANDX1 G28647 (.A1(W15489), .A2(W13406), .ZN(W15626));
  NANDX1 G28648 (.A1(I267), .A2(W3118), .ZN(W6562));
  NANDX1 G28649 (.A1(W4407), .A2(W10914), .ZN(W15623));
  NANDX1 G28650 (.A1(W661), .A2(W5176), .ZN(W14616));
  NANDX1 G28651 (.A1(W13585), .A2(W13406), .ZN(O889));
  NANDX1 G28652 (.A1(W13400), .A2(W6370), .ZN(W15660));
  NANDX1 G28653 (.A1(W3998), .A2(W5261), .ZN(W6525));
  NANDX1 G28654 (.A1(W744), .A2(W1621), .ZN(O1044));
  NANDX1 G28655 (.A1(W584), .A2(W4111), .ZN(W7193));
  NANDX1 G28656 (.A1(W703), .A2(W4010), .ZN(W7191));
  NANDX1 G28657 (.A1(W3794), .A2(W1614), .ZN(W6528));
  NANDX1 G28658 (.A1(W12846), .A2(W6556), .ZN(W15652));
  NANDX1 G28659 (.A1(W3683), .A2(W959), .ZN(W6565));
  NANDX1 G28660 (.A1(W125), .A2(I208), .ZN(W6531));
  NANDX1 G28661 (.A1(W8063), .A2(I492), .ZN(W15650));
  NANDX1 G28662 (.A1(W1616), .A2(W10744), .ZN(W14618));
  NANDX1 G28663 (.A1(W840), .A2(W3743), .ZN(W6545));
  NANDX1 G28664 (.A1(I1482), .A2(W1932), .ZN(W6546));
  NANDX1 G28665 (.A1(W5536), .A2(W13498), .ZN(W15646));
  NANDX1 G28666 (.A1(W1711), .A2(W2995), .ZN(W6547));
  NANDX1 G28667 (.A1(W5480), .A2(W3625), .ZN(W6550));
  NANDX1 G28668 (.A1(W8849), .A2(W3413), .ZN(W15580));
  NANDX1 G28669 (.A1(W3446), .A2(I1798), .ZN(W15593));
  NANDX1 G28670 (.A1(W5649), .A2(I1972), .ZN(W6574));
  NANDX1 G28671 (.A1(W4447), .A2(W3740), .ZN(W6575));
  NANDX1 G28672 (.A1(W2690), .A2(W829), .ZN(W14631));
  NANDX1 G28673 (.A1(W1498), .A2(I1634), .ZN(W6576));
  NANDX1 G28674 (.A1(W6405), .A2(W1755), .ZN(W15591));
  NANDX1 G28675 (.A1(W3121), .A2(W1781), .ZN(W7179));
  NANDX1 G28676 (.A1(W14157), .A2(W10838), .ZN(W15585));
  NANDX1 G28677 (.A1(W8472), .A2(W1340), .ZN(O891));
  NANDX1 G28678 (.A1(W10883), .A2(W7501), .ZN(W14632));
  NANDX1 G28679 (.A1(W4882), .A2(W2785), .ZN(O892));
  NANDX1 G28680 (.A1(W8837), .A2(W3732), .ZN(W14636));
  NANDX1 G28681 (.A1(W4766), .A2(W3211), .ZN(W6586));
  NANDX1 G28682 (.A1(W1929), .A2(W10488), .ZN(W15575));
  NANDX1 G28683 (.A1(W2172), .A2(W14843), .ZN(O1031));
  NANDX1 G28684 (.A1(W1662), .A2(I1177), .ZN(W7176));
  NANDX1 G28685 (.A1(W3521), .A2(W11375), .ZN(W14638));
  NANDX1 G28686 (.A1(W308), .A2(W15064), .ZN(W15605));
  NANDX1 G28687 (.A1(W2437), .A2(W6746), .ZN(O1040));
  NANDX1 G28688 (.A1(W2788), .A2(W14199), .ZN(W15621));
  NANDX1 G28689 (.A1(W1210), .A2(W15564), .ZN(W15619));
  NANDX1 G28690 (.A1(W5595), .A2(W3745), .ZN(W7183));
  NANDX1 G28691 (.A1(W12662), .A2(I1078), .ZN(W15615));
  NANDX1 G28692 (.A1(W1030), .A2(I238), .ZN(W6568));
  NANDX1 G28693 (.A1(W3190), .A2(W3044), .ZN(O1036));
  NANDX1 G28694 (.A1(W8692), .A2(W2189), .ZN(O1034));
  NANDX1 G28695 (.A1(W7344), .A2(W13251), .ZN(W15478));
  NANDX1 G28696 (.A1(W11278), .A2(W911), .ZN(W14628));
  NANDX1 G28697 (.A1(I927), .A2(W3038), .ZN(W7182));
  NANDX1 G28698 (.A1(W3251), .A2(W6696), .ZN(W15603));
  NANDX1 G28699 (.A1(W446), .A2(W4781), .ZN(W6571));
  NANDX1 G28700 (.A1(W4072), .A2(W13018), .ZN(W15602));
  NANDX1 G28701 (.A1(I382), .A2(W7866), .ZN(O1033));
  NANDX1 G28702 (.A1(W8513), .A2(W4236), .ZN(W15597));
  NANDX1 G28703 (.A1(W4004), .A2(W2167), .ZN(W6572));
  NANDX1 G28704 (.A1(I1820), .A2(W13479), .ZN(O992));
  NANDX1 G28705 (.A1(W13552), .A2(W4591), .ZN(W14733));
  NANDX1 G28706 (.A1(W4452), .A2(W8240), .ZN(W14734));
  NANDX1 G28707 (.A1(W4020), .A2(W6872), .ZN(O994));
  NANDX1 G28708 (.A1(W1657), .A2(W4203), .ZN(W6708));
  NANDX1 G28709 (.A1(W10780), .A2(I1669), .ZN(W15339));
  NANDX1 G28710 (.A1(W306), .A2(W11714), .ZN(W15338));
  NANDX1 G28711 (.A1(W506), .A2(I255), .ZN(W14736));
  NANDX1 G28712 (.A1(W1643), .A2(I778), .ZN(W15337));
  NANDX1 G28713 (.A1(I1628), .A2(W1412), .ZN(O144));
  NANDX1 G28714 (.A1(W2392), .A2(W4949), .ZN(W6705));
  NANDX1 G28715 (.A1(W4368), .A2(W3713), .ZN(O145));
  NANDX1 G28716 (.A1(W3351), .A2(W12382), .ZN(O991));
  NANDX1 G28717 (.A1(I592), .A2(W3803), .ZN(W7091));
  NANDX1 G28718 (.A1(W7732), .A2(W11891), .ZN(W15325));
  NANDX1 G28719 (.A1(W2391), .A2(W5110), .ZN(W6718));
  NANDX1 G28720 (.A1(I539), .A2(W5956), .ZN(W7087));
  NANDX1 G28721 (.A1(W1158), .A2(W7845), .ZN(O989));
  NANDX1 G28722 (.A1(W7686), .A2(W8137), .ZN(W15317));
  NANDX1 G28723 (.A1(W66), .A2(I1114), .ZN(W7097));
  NANDX1 G28724 (.A1(W9855), .A2(W5262), .ZN(W15367));
  NANDX1 G28725 (.A1(W483), .A2(W3061), .ZN(W15366));
  NANDX1 G28726 (.A1(W4185), .A2(W3758), .ZN(W15365));
  NANDX1 G28727 (.A1(W1759), .A2(W8574), .ZN(W15361));
  NANDX1 G28728 (.A1(W324), .A2(I1795), .ZN(W7099));
  NANDX1 G28729 (.A1(W1785), .A2(W6576), .ZN(W6693));
  NANDX1 G28730 (.A1(W4874), .A2(I1432), .ZN(W6697));
  NANDX1 G28731 (.A1(I347), .A2(W4448), .ZN(W6699));
  NANDX1 G28732 (.A1(W6769), .A2(I1984), .ZN(W14741));
  NANDX1 G28733 (.A1(W6171), .A2(W2530), .ZN(W15351));
  NANDX1 G28734 (.A1(W290), .A2(W5607), .ZN(W6701));
  NANDX1 G28735 (.A1(W1377), .A2(W13361), .ZN(W15350));
  NANDX1 G28736 (.A1(W662), .A2(W658), .ZN(W6703));
  NANDX1 G28737 (.A1(W5815), .A2(W3766), .ZN(W7093));
  NANDX1 G28738 (.A1(W6285), .A2(W7929), .ZN(W15346));
  NANDX1 G28739 (.A1(W826), .A2(W7969), .ZN(W15345));
  NANDX1 G28740 (.A1(W3456), .A2(I420), .ZN(W6704));
  NANDX1 G28741 (.A1(W12578), .A2(W14034), .ZN(O984));
  NANDX1 G28742 (.A1(W14428), .A2(W12138), .ZN(W14752));
  NANDX1 G28743 (.A1(W878), .A2(I456), .ZN(W14756));
  NANDX1 G28744 (.A1(W9661), .A2(W11511), .ZN(W15290));
  NANDX1 G28745 (.A1(W13279), .A2(W12495), .ZN(W14757));
  NANDX1 G28746 (.A1(W249), .A2(W8628), .ZN(W15286));
  NANDX1 G28747 (.A1(W1422), .A2(W5800), .ZN(W6742));
  NANDX1 G28748 (.A1(W5695), .A2(W14070), .ZN(W14762));
  NANDX1 G28749 (.A1(W4791), .A2(W6572), .ZN(W6745));
  NANDX1 G28750 (.A1(W11), .A2(W12806), .ZN(W15293));
  NANDX1 G28751 (.A1(W4335), .A2(I1202), .ZN(W14765));
  NANDX1 G28752 (.A1(W8764), .A2(W12075), .ZN(W15279));
  NANDX1 G28753 (.A1(W5144), .A2(W6506), .ZN(W6746));
  NANDX1 G28754 (.A1(W13690), .A2(W3263), .ZN(W15278));
  NANDX1 G28755 (.A1(W2171), .A2(I1600), .ZN(O983));
  NANDX1 G28756 (.A1(W443), .A2(W2642), .ZN(W14766));
  NANDX1 G28757 (.A1(W4247), .A2(W401), .ZN(W6747));
  NANDX1 G28758 (.A1(W3316), .A2(W14569), .ZN(W14767));
  NANDX1 G28759 (.A1(W3088), .A2(W1169), .ZN(W6734));
  NANDX1 G28760 (.A1(W8608), .A2(W11270), .ZN(O911));
  NANDX1 G28761 (.A1(W2960), .A2(I170), .ZN(W6722));
  NANDX1 G28762 (.A1(W1192), .A2(W1457), .ZN(W6723));
  NANDX1 G28763 (.A1(W1004), .A2(W14450), .ZN(W15315));
  NANDX1 G28764 (.A1(W7736), .A2(W4507), .ZN(W15309));
  NANDX1 G28765 (.A1(W2178), .A2(W4291), .ZN(W6728));
  NANDX1 G28766 (.A1(W3815), .A2(W3879), .ZN(W6730));
  NANDX1 G28767 (.A1(W3421), .A2(W3940), .ZN(W6733));
  NANDX1 G28768 (.A1(W3703), .A2(W2123), .ZN(W15368));
  NANDX1 G28769 (.A1(W4940), .A2(W5688), .ZN(O912));
  NANDX1 G28770 (.A1(W5508), .A2(W1924), .ZN(W14745));
  NANDX1 G28771 (.A1(W4934), .A2(I1934), .ZN(W6735));
  NANDX1 G28772 (.A1(W4765), .A2(W5245), .ZN(W15303));
  NANDX1 G28773 (.A1(W5636), .A2(W4484), .ZN(W15299));
  NANDX1 G28774 (.A1(W4238), .A2(W4296), .ZN(W6736));
  NANDX1 G28775 (.A1(W5479), .A2(W3896), .ZN(W7078));
  NANDX1 G28776 (.A1(W6069), .A2(W5870), .ZN(O148));
  NANDX1 G28777 (.A1(W1019), .A2(W362), .ZN(W15428));
  NANDX1 G28778 (.A1(I186), .A2(W5821), .ZN(W7139));
  NANDX1 G28779 (.A1(W6644), .A2(W2138), .ZN(W6659));
  NANDX1 G28780 (.A1(W3162), .A2(W3768), .ZN(W7137));
  NANDX1 G28781 (.A1(W4899), .A2(W1748), .ZN(O141));
  NANDX1 G28782 (.A1(I203), .A2(W722), .ZN(W7135));
  NANDX1 G28783 (.A1(W4389), .A2(I1996), .ZN(W7134));
  NANDX1 G28784 (.A1(W12541), .A2(I466), .ZN(O1006));
  NANDX1 G28785 (.A1(W9509), .A2(W433), .ZN(W15434));
  NANDX1 G28786 (.A1(W14570), .A2(W2647), .ZN(W15430));
  NANDX1 G28787 (.A1(W1924), .A2(W11033), .ZN(W15440));
  NANDX1 G28788 (.A1(W11989), .A2(W7001), .ZN(O902));
  NANDX1 G28789 (.A1(W1423), .A2(W8190), .ZN(W14695));
  NANDX1 G28790 (.A1(W812), .A2(W3416), .ZN(W7131));
  NANDX1 G28791 (.A1(W10015), .A2(W7254), .ZN(W15419));
  NANDX1 G28792 (.A1(W855), .A2(W12181), .ZN(W15416));
  NANDX1 G28793 (.A1(W12687), .A2(I1622), .ZN(W15415));
  NANDX1 G28794 (.A1(W6452), .A2(W6254), .ZN(W6668));
  NANDX1 G28795 (.A1(W9211), .A2(W3398), .ZN(W14699));
  NANDX1 G28796 (.A1(W9316), .A2(W9350), .ZN(W15461));
  NANDX1 G28797 (.A1(W5200), .A2(W4084), .ZN(W7155));
  NANDX1 G28798 (.A1(W2278), .A2(W2035), .ZN(W6643));
  NANDX1 G28799 (.A1(W798), .A2(W7068), .ZN(W7152));
  NANDX1 G28800 (.A1(W14164), .A2(W2113), .ZN(O901));
  NANDX1 G28801 (.A1(W3743), .A2(W2740), .ZN(O1013));
  NANDX1 G28802 (.A1(W7268), .A2(W15155), .ZN(O1011));
  NANDX1 G28803 (.A1(W5486), .A2(W5362), .ZN(W15465));
  NANDX1 G28804 (.A1(W5011), .A2(W10371), .ZN(W15464));
  NANDX1 G28805 (.A1(W14444), .A2(W14532), .ZN(O903));
  NANDX1 G28806 (.A1(W1327), .A2(I1877), .ZN(O140));
  NANDX1 G28807 (.A1(W6780), .A2(W5643), .ZN(W7149));
  NANDX1 G28808 (.A1(W3977), .A2(W6589), .ZN(W6654));
  NANDX1 G28809 (.A1(W14371), .A2(W8790), .ZN(W15452));
  NANDX1 G28810 (.A1(I1213), .A2(W2284), .ZN(W6657));
  NANDX1 G28811 (.A1(W6251), .A2(W296), .ZN(W7143));
  NANDX1 G28812 (.A1(W11956), .A2(W8969), .ZN(W15441));
  NANDX1 G28813 (.A1(W1139), .A2(W3018), .ZN(W7142));
  NANDX1 G28814 (.A1(W14630), .A2(I1177), .ZN(W15384));
  NANDX1 G28815 (.A1(W7487), .A2(W13005), .ZN(W15393));
  NANDX1 G28816 (.A1(W4696), .A2(W4337), .ZN(W6677));
  NANDX1 G28817 (.A1(W5569), .A2(W1607), .ZN(W7116));
  NANDX1 G28818 (.A1(W2958), .A2(W5416), .ZN(W7115));
  NANDX1 G28819 (.A1(W2951), .A2(W10534), .ZN(W15391));
  NANDX1 G28820 (.A1(I102), .A2(I946), .ZN(O908));
  NANDX1 G28821 (.A1(W6592), .A2(W8652), .ZN(W15389));
  NANDX1 G28822 (.A1(I1229), .A2(W8354), .ZN(W15385));
  NANDX1 G28823 (.A1(W15345), .A2(W2823), .ZN(W15394));
  NANDX1 G28824 (.A1(W4876), .A2(I846), .ZN(W6683));
  NANDX1 G28825 (.A1(W4912), .A2(W5405), .ZN(W6685));
  NANDX1 G28826 (.A1(I1184), .A2(W2459), .ZN(W14722));
  NANDX1 G28827 (.A1(W55), .A2(W5722), .ZN(W14723));
  NANDX1 G28828 (.A1(I1918), .A2(I289), .ZN(O996));
  NANDX1 G28829 (.A1(W9926), .A2(W9132), .ZN(W15373));
  NANDX1 G28830 (.A1(W4076), .A2(W4550), .ZN(W7104));
  NANDX1 G28831 (.A1(W703), .A2(W13979), .ZN(W15369));
  NANDX1 G28832 (.A1(W9182), .A2(W2829), .ZN(W15409));
  NANDX1 G28833 (.A1(W2002), .A2(W3283), .ZN(W7124));
  NANDX1 G28834 (.A1(W1609), .A2(W13422), .ZN(O904));
  NANDX1 G28835 (.A1(W1411), .A2(W12639), .ZN(W15413));
  NANDX1 G28836 (.A1(W5829), .A2(W2646), .ZN(W7122));
  NANDX1 G28837 (.A1(W10253), .A2(W4402), .ZN(W14709));
  NANDX1 G28838 (.A1(W4322), .A2(W6168), .ZN(W6672));
  NANDX1 G28839 (.A1(W2865), .A2(W9150), .ZN(W14711));
  NANDX1 G28840 (.A1(W4822), .A2(W7327), .ZN(W15410));
  NANDX1 G28841 (.A1(W14704), .A2(W2769), .ZN(W16453));
  NANDX1 G28842 (.A1(W8721), .A2(W5718), .ZN(W15408));
  NANDX1 G28843 (.A1(W2972), .A2(W5131), .ZN(W7118));
  NANDX1 G28844 (.A1(W8935), .A2(W3802), .ZN(W15406));
  NANDX1 G28845 (.A1(I978), .A2(W6765), .ZN(W15405));
  NANDX1 G28846 (.A1(W925), .A2(W6806), .ZN(W14713));
  NANDX1 G28847 (.A1(W325), .A2(W14015), .ZN(W15401));
  NANDX1 G28848 (.A1(W322), .A2(I1232), .ZN(W6676));
  NANDX1 G28849 (.A1(W13011), .A2(W636), .ZN(W15398));
  NANDX1 G28850 (.A1(W11131), .A2(W3746), .ZN(W13885));
  NANDX1 G28851 (.A1(I1709), .A2(W14001), .ZN(W17473));
  NANDX1 G28852 (.A1(I1193), .A2(W6801), .ZN(W7696));
  NANDX1 G28853 (.A1(W1949), .A2(W4188), .ZN(W5402));
  NANDX1 G28854 (.A1(W6214), .A2(I1441), .ZN(W7694));
  NANDX1 G28855 (.A1(W4289), .A2(I406), .ZN(W5406));
  NANDX1 G28856 (.A1(W6810), .A2(I923), .ZN(W7693));
  NANDX1 G28857 (.A1(W14), .A2(W2527), .ZN(W7691));
  NANDX1 G28858 (.A1(W11629), .A2(W554), .ZN(W13880));
  NANDX1 G28859 (.A1(W2753), .A2(W2967), .ZN(W17464));
  NANDX1 G28860 (.A1(W4624), .A2(W1312), .ZN(O1398));
  NANDX1 G28861 (.A1(W4645), .A2(W16202), .ZN(W17461));
  NANDX1 G28862 (.A1(W6621), .A2(W1448), .ZN(W13886));
  NANDX1 G28863 (.A1(W1503), .A2(W4068), .ZN(W5415));
  NANDX1 G28864 (.A1(W8375), .A2(W6669), .ZN(W17458));
  NANDX1 G28865 (.A1(W5228), .A2(I1289), .ZN(W7688));
  NANDX1 G28866 (.A1(W6616), .A2(W6565), .ZN(W7685));
  NANDX1 G28867 (.A1(W2957), .A2(W1440), .ZN(W7684));
  NANDX1 G28868 (.A1(W8490), .A2(I290), .ZN(W17451));
  NANDX1 G28869 (.A1(W6685), .A2(W9692), .ZN(O797));
  NANDX1 G28870 (.A1(W5134), .A2(W2057), .ZN(W17494));
  NANDX1 G28871 (.A1(W2741), .A2(W5283), .ZN(W13875));
  NANDX1 G28872 (.A1(W3006), .A2(W1686), .ZN(W5394));
  NANDX1 G28873 (.A1(W3880), .A2(W5584), .ZN(W7699));
  NANDX1 G28874 (.A1(W12818), .A2(W12388), .ZN(W17491));
  NANDX1 G28875 (.A1(W96), .A2(W2552), .ZN(W5395));
  NANDX1 G28876 (.A1(W15208), .A2(W9528), .ZN(W17487));
  NANDX1 G28877 (.A1(I154), .A2(W13546), .ZN(W17484));
  NANDX1 G28878 (.A1(W11812), .A2(W12620), .ZN(W17450));
  NANDX1 G28879 (.A1(W5500), .A2(I1047), .ZN(W17483));
  NANDX1 G28880 (.A1(W6139), .A2(W7590), .ZN(O195));
  NANDX1 G28881 (.A1(W2730), .A2(W761), .ZN(W17482));
  NANDX1 G28882 (.A1(W16244), .A2(W6159), .ZN(W17481));
  NANDX1 G28883 (.A1(W2678), .A2(W2005), .ZN(W5397));
  NANDX1 G28884 (.A1(W8965), .A2(W15131), .ZN(O1399));
  NANDX1 G28885 (.A1(W2570), .A2(I941), .ZN(W5399));
  NANDX1 G28886 (.A1(W6259), .A2(W7495), .ZN(W7697));
  NANDX1 G28887 (.A1(I1332), .A2(W1552), .ZN(W5436));
  NANDX1 G28888 (.A1(W1136), .A2(W12956), .ZN(W17414));
  NANDX1 G28889 (.A1(W1943), .A2(W3997), .ZN(W5427));
  NANDX1 G28890 (.A1(W4704), .A2(W2369), .ZN(W17413));
  NANDX1 G28891 (.A1(W3474), .A2(W1395), .ZN(W7674));
  NANDX1 G28892 (.A1(W782), .A2(W2565), .ZN(W17411));
  NANDX1 G28893 (.A1(W822), .A2(W959), .ZN(W7673));
  NANDX1 G28894 (.A1(W4332), .A2(I1571), .ZN(W5430));
  NANDX1 G28895 (.A1(W5456), .A2(W300), .ZN(W17405));
  NANDX1 G28896 (.A1(W14376), .A2(W10091), .ZN(W17416));
  NANDX1 G28897 (.A1(W2951), .A2(W3439), .ZN(W7669));
  NANDX1 G28898 (.A1(W5100), .A2(W13226), .ZN(O1382));
  NANDX1 G28899 (.A1(W13566), .A2(W15080), .ZN(W17402));
  NANDX1 G28900 (.A1(W13772), .A2(W4934), .ZN(W13904));
  NANDX1 G28901 (.A1(I103), .A2(W3820), .ZN(W5437));
  NANDX1 G28902 (.A1(W1041), .A2(W2895), .ZN(W5438));
  NANDX1 G28903 (.A1(W12299), .A2(W14738), .ZN(W17391));
  NANDX1 G28904 (.A1(W16226), .A2(I326), .ZN(W17390));
  NANDX1 G28905 (.A1(W2804), .A2(W9345), .ZN(W17434));
  NANDX1 G28906 (.A1(W17387), .A2(W3153), .ZN(W17449));
  NANDX1 G28907 (.A1(W16620), .A2(W248), .ZN(W17447));
  NANDX1 G28908 (.A1(W1006), .A2(W5657), .ZN(W17445));
  NANDX1 G28909 (.A1(W9276), .A2(W4696), .ZN(W17444));
  NANDX1 G28910 (.A1(W3551), .A2(W895), .ZN(W17441));
  NANDX1 G28911 (.A1(W2267), .A2(W2535), .ZN(W7680));
  NANDX1 G28912 (.A1(I1637), .A2(W1780), .ZN(W5421));
  NANDX1 G28913 (.A1(W6124), .A2(W16619), .ZN(O1389));
  NANDX1 G28914 (.A1(W2103), .A2(W4923), .ZN(W5390));
  NANDX1 G28915 (.A1(W8315), .A2(W2155), .ZN(O1388));
  NANDX1 G28916 (.A1(W15660), .A2(W3109), .ZN(W17431));
  NANDX1 G28917 (.A1(W4735), .A2(W8143), .ZN(W17430));
  NANDX1 G28918 (.A1(W2499), .A2(I1836), .ZN(W5423));
  NANDX1 G28919 (.A1(W16690), .A2(W1220), .ZN(W17425));
  NANDX1 G28920 (.A1(W8616), .A2(W1063), .ZN(O1385));
  NANDX1 G28921 (.A1(W4230), .A2(W1305), .ZN(W5424));
  NANDX1 G28922 (.A1(W13180), .A2(W5499), .ZN(W17418));
  NANDX1 G28923 (.A1(W8320), .A2(W11535), .ZN(W17535));
  NANDX1 G28924 (.A1(W5994), .A2(W11338), .ZN(O791));
  NANDX1 G28925 (.A1(W2945), .A2(W3283), .ZN(W5345));
  NANDX1 G28926 (.A1(W1319), .A2(W1032), .ZN(W5347));
  NANDX1 G28927 (.A1(I1325), .A2(W12033), .ZN(W17543));
  NANDX1 G28928 (.A1(W11747), .A2(W5242), .ZN(O792));
  NANDX1 G28929 (.A1(I348), .A2(W2146), .ZN(W7713));
  NANDX1 G28930 (.A1(W14206), .A2(W12726), .ZN(W17539));
  NANDX1 G28931 (.A1(W4516), .A2(W1049), .ZN(W5352));
  NANDX1 G28932 (.A1(W1861), .A2(W12084), .ZN(W17536));
  NANDX1 G28933 (.A1(W10627), .A2(W3677), .ZN(W13847));
  NANDX1 G28934 (.A1(W5162), .A2(I716), .ZN(W13853));
  NANDX1 G28935 (.A1(W6325), .A2(W1263), .ZN(W17534));
  NANDX1 G28936 (.A1(I145), .A2(W1389), .ZN(W5357));
  NANDX1 G28937 (.A1(W15651), .A2(W7169), .ZN(W17531));
  NANDX1 G28938 (.A1(W589), .A2(W195), .ZN(O83));
  NANDX1 G28939 (.A1(W108), .A2(W7354), .ZN(W13855));
  NANDX1 G28940 (.A1(I501), .A2(W2931), .ZN(W7709));
  NANDX1 G28941 (.A1(W5717), .A2(W9246), .ZN(W13857));
  NANDX1 G28942 (.A1(W813), .A2(W4887), .ZN(W7715));
  NANDX1 G28943 (.A1(W2016), .A2(I414), .ZN(W7721));
  NANDX1 G28944 (.A1(W5841), .A2(W12998), .ZN(W17566));
  NANDX1 G28945 (.A1(W12646), .A2(W11481), .ZN(W17563));
  NANDX1 G28946 (.A1(W13115), .A2(W13064), .ZN(W13835));
  NANDX1 G28947 (.A1(W1036), .A2(W1503), .ZN(W7718));
  NANDX1 G28948 (.A1(W5380), .A2(W6148), .ZN(W7716));
  NANDX1 G28949 (.A1(W7071), .A2(W3960), .ZN(W13838));
  NANDX1 G28950 (.A1(W904), .A2(W17060), .ZN(W17561));
  NANDX1 G28951 (.A1(W3975), .A2(I1370), .ZN(W5362));
  NANDX1 G28952 (.A1(W16196), .A2(I919), .ZN(W17557));
  NANDX1 G28953 (.A1(W3330), .A2(W10610), .ZN(W13840));
  NANDX1 G28954 (.A1(I1277), .A2(I1078), .ZN(W5338));
  NANDX1 G28955 (.A1(W2946), .A2(W7973), .ZN(W17555));
  NANDX1 G28956 (.A1(W9596), .A2(W452), .ZN(W17554));
  NANDX1 G28957 (.A1(W1448), .A2(W12693), .ZN(W17553));
  NANDX1 G28958 (.A1(W1432), .A2(W11575), .ZN(W13843));
  NANDX1 G28959 (.A1(W2904), .A2(I409), .ZN(W7714));
  NANDX1 G28960 (.A1(W1641), .A2(W9619), .ZN(W13872));
  NANDX1 G28961 (.A1(W2623), .A2(W3316), .ZN(W13870));
  NANDX1 G28962 (.A1(W2473), .A2(W2272), .ZN(W17504));
  NANDX1 G28963 (.A1(W4850), .A2(W2090), .ZN(W5374));
  NANDX1 G28964 (.A1(W2819), .A2(I992), .ZN(W7704));
  NANDX1 G28965 (.A1(W3358), .A2(W1119), .ZN(W5375));
  NANDX1 G28966 (.A1(W4715), .A2(W6905), .ZN(W7703));
  NANDX1 G28967 (.A1(W1721), .A2(W1123), .ZN(W5380));
  NANDX1 G28968 (.A1(W6978), .A2(I914), .ZN(W7701));
  NANDX1 G28969 (.A1(W3227), .A2(W13098), .ZN(O1403));
  NANDX1 G28970 (.A1(W471), .A2(W8202), .ZN(W17501));
  NANDX1 G28971 (.A1(W16494), .A2(W5745), .ZN(W17500));
  NANDX1 G28972 (.A1(W1196), .A2(W7544), .ZN(W17499));
  NANDX1 G28973 (.A1(I387), .A2(W2012), .ZN(W5388));
  NANDX1 G28974 (.A1(I1603), .A2(W2988), .ZN(W17498));
  NANDX1 G28975 (.A1(W13304), .A2(W12945), .ZN(W13873));
  NANDX1 G28976 (.A1(W7022), .A2(W10046), .ZN(W17496));
  NANDX1 G28977 (.A1(I1889), .A2(W3607), .ZN(W5389));
  NANDX1 G28978 (.A1(W9586), .A2(W9331), .ZN(W17513));
  NANDX1 G28979 (.A1(W846), .A2(W8314), .ZN(W17525));
  NANDX1 G28980 (.A1(W7019), .A2(W1756), .ZN(O1408));
  NANDX1 G28981 (.A1(W1660), .A2(W2480), .ZN(W5364));
  NANDX1 G28982 (.A1(W2004), .A2(W4288), .ZN(W5366));
  NANDX1 G28983 (.A1(W3242), .A2(I707), .ZN(W13862));
  NANDX1 G28984 (.A1(W13646), .A2(W12548), .ZN(W17516));
  NANDX1 G28985 (.A1(W473), .A2(W3838), .ZN(W5367));
  NANDX1 G28986 (.A1(W10207), .A2(W847), .ZN(O795));
  NANDX1 G28987 (.A1(W5258), .A2(W5730), .ZN(W7666));
  NANDX1 G28988 (.A1(W6159), .A2(W955), .ZN(O1405));
  NANDX1 G28989 (.A1(I724), .A2(I787), .ZN(W5369));
  NANDX1 G28990 (.A1(W8139), .A2(W3693), .ZN(O796));
  NANDX1 G28991 (.A1(W5254), .A2(W1531), .ZN(W5372));
  NANDX1 G28992 (.A1(W11825), .A2(W4650), .ZN(W13866));
  NANDX1 G28993 (.A1(W11160), .A2(I70), .ZN(W17508));
  NANDX1 G28994 (.A1(I735), .A2(W2027), .ZN(W17507));
  NANDX1 G28995 (.A1(W1376), .A2(I818), .ZN(W5373));
  NANDX1 G28996 (.A1(W3909), .A2(W797), .ZN(W5512));
  NANDX1 G28997 (.A1(W3666), .A2(W1443), .ZN(W5504));
  NANDX1 G28998 (.A1(W1180), .A2(I1743), .ZN(W5505));
  NANDX1 G28999 (.A1(W1858), .A2(W10901), .ZN(W17284));
  NANDX1 G29000 (.A1(W13899), .A2(W12758), .ZN(W13951));
  NANDX1 G29001 (.A1(I1198), .A2(W14967), .ZN(W17277));
  NANDX1 G29002 (.A1(W2579), .A2(W1392), .ZN(W5507));
  NANDX1 G29003 (.A1(W5285), .A2(W585), .ZN(W17273));
  NANDX1 G29004 (.A1(W304), .A2(W158), .ZN(W5511));
  NANDX1 G29005 (.A1(W9969), .A2(W15448), .ZN(W17271));
  NANDX1 G29006 (.A1(W5249), .A2(W2706), .ZN(W5503));
  NANDX1 G29007 (.A1(W10591), .A2(W14479), .ZN(O1359));
  NANDX1 G29008 (.A1(W17043), .A2(W15621), .ZN(W17268));
  NANDX1 G29009 (.A1(W728), .A2(W4043), .ZN(W5513));
  NANDX1 G29010 (.A1(W1194), .A2(W2509), .ZN(W5514));
  NANDX1 G29011 (.A1(W4403), .A2(W4784), .ZN(W7624));
  NANDX1 G29012 (.A1(W13829), .A2(W12452), .ZN(W13956));
  NANDX1 G29013 (.A1(W542), .A2(W1358), .ZN(W5516));
  NANDX1 G29014 (.A1(W7396), .A2(W3669), .ZN(O810));
  NANDX1 G29015 (.A1(W1433), .A2(W5403), .ZN(W5499));
  NANDX1 G29016 (.A1(W11611), .A2(W4091), .ZN(W13947));
  NANDX1 G29017 (.A1(W4010), .A2(W16450), .ZN(W17307));
  NANDX1 G29018 (.A1(W10183), .A2(W5273), .ZN(W17305));
  NANDX1 G29019 (.A1(I1894), .A2(W16636), .ZN(W17304));
  NANDX1 G29020 (.A1(W4944), .A2(W11212), .ZN(O1366));
  NANDX1 G29021 (.A1(W4680), .A2(W15041), .ZN(O1365));
  NANDX1 G29022 (.A1(W5402), .A2(W1432), .ZN(W7629));
  NANDX1 G29023 (.A1(I1652), .A2(I1215), .ZN(W17298));
  NANDX1 G29024 (.A1(W5271), .A2(I475), .ZN(W17266));
  NANDX1 G29025 (.A1(W14120), .A2(W5525), .ZN(W17296));
  NANDX1 G29026 (.A1(W11178), .A2(W1154), .ZN(W17293));
  NANDX1 G29027 (.A1(W11226), .A2(W7288), .ZN(W17291));
  NANDX1 G29028 (.A1(W12742), .A2(I600), .ZN(W17290));
  NANDX1 G29029 (.A1(W9340), .A2(W4866), .ZN(W17289));
  NANDX1 G29030 (.A1(W7367), .A2(W2729), .ZN(W7628));
  NANDX1 G29031 (.A1(W8270), .A2(W9990), .ZN(W13950));
  NANDX1 G29032 (.A1(W14919), .A2(W15926), .ZN(W17286));
  NANDX1 G29033 (.A1(W4928), .A2(I1136), .ZN(W17234));
  NANDX1 G29034 (.A1(W796), .A2(W10012), .ZN(O1353));
  NANDX1 G29035 (.A1(I1535), .A2(W8083), .ZN(W13973));
  NANDX1 G29036 (.A1(I1654), .A2(W3895), .ZN(W5535));
  NANDX1 G29037 (.A1(W840), .A2(W2974), .ZN(W17242));
  NANDX1 G29038 (.A1(W2313), .A2(W4914), .ZN(W5536));
  NANDX1 G29039 (.A1(I760), .A2(W1075), .ZN(W17241));
  NANDX1 G29040 (.A1(W3180), .A2(W13710), .ZN(W13977));
  NANDX1 G29041 (.A1(W3512), .A2(I420), .ZN(W5538));
  NANDX1 G29042 (.A1(W758), .A2(W14219), .ZN(O1354));
  NANDX1 G29043 (.A1(W2713), .A2(W6424), .ZN(W17233));
  NANDX1 G29044 (.A1(W5878), .A2(W5641), .ZN(W7616));
  NANDX1 G29045 (.A1(I1380), .A2(W3534), .ZN(W7615));
  NANDX1 G29046 (.A1(W1039), .A2(W4802), .ZN(W5544));
  NANDX1 G29047 (.A1(W7462), .A2(W7661), .ZN(W17231));
  NANDX1 G29048 (.A1(I793), .A2(W4889), .ZN(W7614));
  NANDX1 G29049 (.A1(I194), .A2(W6536), .ZN(W17229));
  NANDX1 G29050 (.A1(W14266), .A2(W2794), .ZN(W17228));
  NANDX1 G29051 (.A1(I1232), .A2(W4461), .ZN(W5521));
  NANDX1 G29052 (.A1(W650), .A2(W2275), .ZN(W17265));
  NANDX1 G29053 (.A1(W2266), .A2(I1459), .ZN(O89));
  NANDX1 G29054 (.A1(W10221), .A2(W8812), .ZN(W13958));
  NANDX1 G29055 (.A1(W4566), .A2(W2222), .ZN(W5520));
  NANDX1 G29056 (.A1(W15526), .A2(W13332), .ZN(W17261));
  NANDX1 G29057 (.A1(W6965), .A2(I920), .ZN(W17260));
  NANDX1 G29058 (.A1(W8110), .A2(W4012), .ZN(W17259));
  NANDX1 G29059 (.A1(W13762), .A2(W45), .ZN(W13960));
  NANDX1 G29060 (.A1(W1079), .A2(W3126), .ZN(W5496));
  NANDX1 G29061 (.A1(W13127), .A2(W5123), .ZN(W13961));
  NANDX1 G29062 (.A1(W6925), .A2(I1889), .ZN(O1357));
  NANDX1 G29063 (.A1(W13056), .A2(W11619), .ZN(W17253));
  NANDX1 G29064 (.A1(W4304), .A2(I1005), .ZN(W5526));
  NANDX1 G29065 (.A1(W3322), .A2(W6468), .ZN(W7618));
  NANDX1 G29066 (.A1(W13), .A2(W564), .ZN(W5529));
  NANDX1 G29067 (.A1(W9246), .A2(W11139), .ZN(W17249));
  NANDX1 G29068 (.A1(W1081), .A2(I1277), .ZN(W5532));
  NANDX1 G29069 (.A1(W3654), .A2(I1937), .ZN(W5464));
  NANDX1 G29070 (.A1(W3080), .A2(W4752), .ZN(O85));
  NANDX1 G29071 (.A1(W1602), .A2(W5463), .ZN(W13915));
  NANDX1 G29072 (.A1(W1133), .A2(I978), .ZN(W13920));
  NANDX1 G29073 (.A1(W10943), .A2(W661), .ZN(W13921));
  NANDX1 G29074 (.A1(W5251), .A2(I9), .ZN(W17359));
  NANDX1 G29075 (.A1(W909), .A2(W3237), .ZN(W5463));
  NANDX1 G29076 (.A1(W8500), .A2(W6272), .ZN(W17354));
  NANDX1 G29077 (.A1(W4626), .A2(W2672), .ZN(W17353));
  NANDX1 G29078 (.A1(W11008), .A2(I229), .ZN(W17351));
  NANDX1 G29079 (.A1(W3759), .A2(W1017), .ZN(W17363));
  NANDX1 G29080 (.A1(W8066), .A2(W2004), .ZN(W17350));
  NANDX1 G29081 (.A1(W6672), .A2(W3684), .ZN(W13922));
  NANDX1 G29082 (.A1(W3074), .A2(W3626), .ZN(O1376));
  NANDX1 G29083 (.A1(W16698), .A2(W4861), .ZN(W17348));
  NANDX1 G29084 (.A1(W4555), .A2(I642), .ZN(W7647));
  NANDX1 G29085 (.A1(W12477), .A2(W471), .ZN(W13923));
  NANDX1 G29086 (.A1(I1255), .A2(W4567), .ZN(W5467));
  NANDX1 G29087 (.A1(W5557), .A2(W5587), .ZN(W7646));
  NANDX1 G29088 (.A1(W2417), .A2(W1669), .ZN(W5454));
  NANDX1 G29089 (.A1(W14928), .A2(W4476), .ZN(W17389));
  NANDX1 G29090 (.A1(W1379), .A2(W1879), .ZN(W5443));
  NANDX1 G29091 (.A1(W10334), .A2(W9284), .ZN(W13910));
  NANDX1 G29092 (.A1(W1866), .A2(W3687), .ZN(W7659));
  NANDX1 G29093 (.A1(W7652), .A2(W3434), .ZN(W7656));
  NANDX1 G29094 (.A1(I792), .A2(W1033), .ZN(W7654));
  NANDX1 G29095 (.A1(W16912), .A2(W4039), .ZN(W17382));
  NANDX1 G29096 (.A1(W5052), .A2(W1168), .ZN(W7653));
  NANDX1 G29097 (.A1(W4688), .A2(W3481), .ZN(W5470));
  NANDX1 G29098 (.A1(W432), .A2(W5018), .ZN(W5455));
  NANDX1 G29099 (.A1(W7941), .A2(W1624), .ZN(W17379));
  NANDX1 G29100 (.A1(W15312), .A2(W14789), .ZN(W17377));
  NANDX1 G29101 (.A1(I1429), .A2(W4552), .ZN(W5456));
  NANDX1 G29102 (.A1(W15988), .A2(W14328), .ZN(W17375));
  NANDX1 G29103 (.A1(W501), .A2(W3475), .ZN(W17374));
  NANDX1 G29104 (.A1(W7720), .A2(W14357), .ZN(W17371));
  NANDX1 G29105 (.A1(W1935), .A2(W15161), .ZN(W17370));
  NANDX1 G29106 (.A1(W8994), .A2(W7222), .ZN(W17319));
  NANDX1 G29107 (.A1(W1632), .A2(I992), .ZN(W5483));
  NANDX1 G29108 (.A1(W14707), .A2(W571), .ZN(W17329));
  NANDX1 G29109 (.A1(W4079), .A2(W4710), .ZN(O87));
  NANDX1 G29110 (.A1(W4974), .A2(I1788), .ZN(W5487));
  NANDX1 G29111 (.A1(W11656), .A2(W11725), .ZN(W17327));
  NANDX1 G29112 (.A1(W8573), .A2(W6325), .ZN(W13935));
  NANDX1 G29113 (.A1(W418), .A2(W169), .ZN(W5490));
  NANDX1 G29114 (.A1(I509), .A2(W14703), .ZN(W17320));
  NANDX1 G29115 (.A1(W7299), .A2(W6209), .ZN(W13933));
  NANDX1 G29116 (.A1(W2650), .A2(W3896), .ZN(W17318));
  NANDX1 G29117 (.A1(W4964), .A2(W441), .ZN(W5491));
  NANDX1 G29118 (.A1(W14388), .A2(W4498), .ZN(W17316));
  NANDX1 G29119 (.A1(W2205), .A2(W2059), .ZN(W7632));
  NANDX1 G29120 (.A1(W1513), .A2(W9479), .ZN(W13942));
  NANDX1 G29121 (.A1(W3753), .A2(W8191), .ZN(W13943));
  NANDX1 G29122 (.A1(W4767), .A2(W1211), .ZN(W5493));
  NANDX1 G29123 (.A1(W6425), .A2(W13172), .ZN(W13946));
  NANDX1 G29124 (.A1(W3027), .A2(W5922), .ZN(W17335));
  NANDX1 G29125 (.A1(W5313), .A2(W3480), .ZN(W5471));
  NANDX1 G29126 (.A1(W10176), .A2(W13587), .ZN(W17343));
  NANDX1 G29127 (.A1(I1398), .A2(W994), .ZN(W5474));
  NANDX1 G29128 (.A1(W4712), .A2(W4702), .ZN(W5475));
  NANDX1 G29129 (.A1(W8962), .A2(W9432), .ZN(W17340));
  NANDX1 G29130 (.A1(W13664), .A2(W11432), .ZN(W13928));
  NANDX1 G29131 (.A1(W5306), .A2(W174), .ZN(W5476));
  NANDX1 G29132 (.A1(W2117), .A2(W353), .ZN(W7644));
  NANDX1 G29133 (.A1(W2600), .A2(W685), .ZN(W5329));
  NANDX1 G29134 (.A1(W10230), .A2(W9206), .ZN(W13929));
  NANDX1 G29135 (.A1(W13378), .A2(W10124), .ZN(W17334));
  NANDX1 G29136 (.A1(W2725), .A2(W4089), .ZN(W5478));
  NANDX1 G29137 (.A1(W7851), .A2(W3786), .ZN(W17332));
  NANDX1 G29138 (.A1(I1552), .A2(W6834), .ZN(W7643));
  NANDX1 G29139 (.A1(I1547), .A2(W3934), .ZN(W5480));
  NANDX1 G29140 (.A1(W1347), .A2(W511), .ZN(O191));
  NANDX1 G29141 (.A1(W7388), .A2(W5744), .ZN(W13932));
  NANDX1 G29142 (.A1(W4789), .A2(W692), .ZN(W7810));
  NANDX1 G29143 (.A1(I819), .A2(W8055), .ZN(W13713));
  NANDX1 G29144 (.A1(I1565), .A2(W12238), .ZN(W13715));
  NANDX1 G29145 (.A1(W1843), .A2(W3079), .ZN(W7817));
  NANDX1 G29146 (.A1(W13365), .A2(W6723), .ZN(W17814));
  NANDX1 G29147 (.A1(W7391), .A2(W3834), .ZN(W7816));
  NANDX1 G29148 (.A1(W1228), .A2(W78), .ZN(W5180));
  NANDX1 G29149 (.A1(W4732), .A2(I151), .ZN(W5181));
  NANDX1 G29150 (.A1(W3224), .A2(W3915), .ZN(W7811));
  NANDX1 G29151 (.A1(I690), .A2(W1284), .ZN(W5183));
  NANDX1 G29152 (.A1(W3316), .A2(W3785), .ZN(W5177));
  NANDX1 G29153 (.A1(W10601), .A2(W11021), .ZN(W17806));
  NANDX1 G29154 (.A1(W13207), .A2(W403), .ZN(W13722));
  NANDX1 G29155 (.A1(W6242), .A2(W7769), .ZN(W7809));
  NANDX1 G29156 (.A1(W6943), .A2(W7897), .ZN(W17801));
  NANDX1 G29157 (.A1(I398), .A2(W7859), .ZN(W13727));
  NANDX1 G29158 (.A1(W14833), .A2(I1686), .ZN(W17798));
  NANDX1 G29159 (.A1(W8687), .A2(W6640), .ZN(W17794));
  NANDX1 G29160 (.A1(W1106), .A2(W1546), .ZN(W5188));
  NANDX1 G29161 (.A1(W11852), .A2(W15305), .ZN(W17831));
  NANDX1 G29162 (.A1(W12089), .A2(W3789), .ZN(W17837));
  NANDX1 G29163 (.A1(W1313), .A2(W811), .ZN(W5164));
  NANDX1 G29164 (.A1(W14996), .A2(W12167), .ZN(W17835));
  NANDX1 G29165 (.A1(I1319), .A2(W3324), .ZN(W5166));
  NANDX1 G29166 (.A1(W6426), .A2(W8013), .ZN(W13706));
  NANDX1 G29167 (.A1(W6391), .A2(W10424), .ZN(W17832));
  NANDX1 G29168 (.A1(W637), .A2(W3064), .ZN(W5167));
  NANDX1 G29169 (.A1(W5346), .A2(I1956), .ZN(W7825));
  NANDX1 G29170 (.A1(W17275), .A2(I1400), .ZN(O1444));
  NANDX1 G29171 (.A1(I1812), .A2(W4281), .ZN(W5170));
  NANDX1 G29172 (.A1(I267), .A2(I1421), .ZN(W17829));
  NANDX1 G29173 (.A1(I690), .A2(I370), .ZN(W5171));
  NANDX1 G29174 (.A1(I120), .A2(I876), .ZN(W7824));
  NANDX1 G29175 (.A1(I1945), .A2(W1302), .ZN(W5173));
  NANDX1 G29176 (.A1(I84), .A2(W3716), .ZN(W7820));
  NANDX1 G29177 (.A1(W9124), .A2(W4323), .ZN(W13712));
  NANDX1 G29178 (.A1(W51), .A2(I914), .ZN(W5176));
  NANDX1 G29179 (.A1(W14302), .A2(W2833), .ZN(W17756));
  NANDX1 G29180 (.A1(W13155), .A2(I1477), .ZN(W17766));
  NANDX1 G29181 (.A1(W4087), .A2(W4043), .ZN(O1440));
  NANDX1 G29182 (.A1(I770), .A2(I445), .ZN(W5203));
  NANDX1 G29183 (.A1(W2399), .A2(W3111), .ZN(W17763));
  NANDX1 G29184 (.A1(W1172), .A2(W6478), .ZN(W7797));
  NANDX1 G29185 (.A1(W43), .A2(I674), .ZN(W5205));
  NANDX1 G29186 (.A1(W16956), .A2(W9568), .ZN(W17759));
  NANDX1 G29187 (.A1(W2618), .A2(W2499), .ZN(W17758));
  NANDX1 G29188 (.A1(W9853), .A2(W954), .ZN(O780));
  NANDX1 G29189 (.A1(W6842), .A2(W15359), .ZN(W17754));
  NANDX1 G29190 (.A1(W193), .A2(W4653), .ZN(W13739));
  NANDX1 G29191 (.A1(W4045), .A2(W1935), .ZN(W5208));
  NANDX1 G29192 (.A1(W13142), .A2(W4365), .ZN(W13741));
  NANDX1 G29193 (.A1(W10675), .A2(W2166), .ZN(W13743));
  NANDX1 G29194 (.A1(W1223), .A2(I550), .ZN(W5209));
  NANDX1 G29195 (.A1(W5039), .A2(W3141), .ZN(W5214));
  NANDX1 G29196 (.A1(I161), .A2(W5883), .ZN(O201));
  NANDX1 G29197 (.A1(W7092), .A2(W8898), .ZN(W17777));
  NANDX1 G29198 (.A1(W1360), .A2(W6367), .ZN(O1443));
  NANDX1 G29199 (.A1(I1181), .A2(W3731), .ZN(W5190));
  NANDX1 G29200 (.A1(I527), .A2(W5670), .ZN(W7805));
  NANDX1 G29201 (.A1(I236), .A2(W8852), .ZN(W17784));
  NANDX1 G29202 (.A1(W5039), .A2(W13240), .ZN(W17782));
  NANDX1 G29203 (.A1(W2150), .A2(W540), .ZN(W5192));
  NANDX1 G29204 (.A1(W6282), .A2(W5981), .ZN(W7804));
  NANDX1 G29205 (.A1(W329), .A2(W3593), .ZN(W17780));
  NANDX1 G29206 (.A1(W193), .A2(I1404), .ZN(W17840));
  NANDX1 G29207 (.A1(W797), .A2(W4094), .ZN(W5196));
  NANDX1 G29208 (.A1(W4993), .A2(W8574), .ZN(W17775));
  NANDX1 G29209 (.A1(W16662), .A2(W1889), .ZN(W17774));
  NANDX1 G29210 (.A1(W13669), .A2(I698), .ZN(W13730));
  NANDX1 G29211 (.A1(I1058), .A2(W3683), .ZN(W5199));
  NANDX1 G29212 (.A1(I1656), .A2(W109), .ZN(W5201));
  NANDX1 G29213 (.A1(W13362), .A2(W10846), .ZN(W17770));
  NANDX1 G29214 (.A1(W3510), .A2(I705), .ZN(W7799));
  NANDX1 G29215 (.A1(I1133), .A2(W7847), .ZN(W17886));
  NANDX1 G29216 (.A1(W4412), .A2(W29), .ZN(W5123));
  NANDX1 G29217 (.A1(W4183), .A2(W2962), .ZN(W5124));
  NANDX1 G29218 (.A1(I774), .A2(W802), .ZN(W5125));
  NANDX1 G29219 (.A1(I1164), .A2(W7044), .ZN(W7835));
  NANDX1 G29220 (.A1(I1794), .A2(I544), .ZN(W5128));
  NANDX1 G29221 (.A1(W15147), .A2(W8452), .ZN(O1465));
  NANDX1 G29222 (.A1(W8886), .A2(W2285), .ZN(W17890));
  NANDX1 G29223 (.A1(I661), .A2(W5880), .ZN(W13676));
  NANDX1 G29224 (.A1(W16754), .A2(W950), .ZN(W17889));
  NANDX1 G29225 (.A1(I1959), .A2(W110), .ZN(W5122));
  NANDX1 G29226 (.A1(I692), .A2(W3300), .ZN(W17884));
  NANDX1 G29227 (.A1(I1087), .A2(W164), .ZN(W7834));
  NANDX1 G29228 (.A1(W6476), .A2(W3240), .ZN(O774));
  NANDX1 G29229 (.A1(I586), .A2(W3193), .ZN(W5130));
  NANDX1 G29230 (.A1(W12082), .A2(W9290), .ZN(W17881));
  NANDX1 G29231 (.A1(W2957), .A2(W14323), .ZN(W17879));
  NANDX1 G29232 (.A1(I1127), .A2(W110), .ZN(W5132));
  NANDX1 G29233 (.A1(W3669), .A2(W3661), .ZN(W5133));
  NANDX1 G29234 (.A1(W4631), .A2(W2719), .ZN(W13667));
  NANDX1 G29235 (.A1(W4083), .A2(W7899), .ZN(W13661));
  NANDX1 G29236 (.A1(I1087), .A2(W4924), .ZN(W5106));
  NANDX1 G29237 (.A1(W373), .A2(W17773), .ZN(W17916));
  NANDX1 G29238 (.A1(W13537), .A2(W3085), .ZN(W13662));
  NANDX1 G29239 (.A1(W5140), .A2(W6590), .ZN(W17915));
  NANDX1 G29240 (.A1(W3913), .A2(W4857), .ZN(W13663));
  NANDX1 G29241 (.A1(W2723), .A2(I674), .ZN(W5114));
  NANDX1 G29242 (.A1(W6990), .A2(W6687), .ZN(W17913));
  NANDX1 G29243 (.A1(W4212), .A2(W16865), .ZN(O1460));
  NANDX1 G29244 (.A1(W5153), .A2(W9232), .ZN(W13670));
  NANDX1 G29245 (.A1(W4076), .A2(W2611), .ZN(W17909));
  NANDX1 G29246 (.A1(W3457), .A2(W4118), .ZN(W7840));
  NANDX1 G29247 (.A1(W151), .A2(W10897), .ZN(W17904));
  NANDX1 G29248 (.A1(W7633), .A2(W1668), .ZN(W13674));
  NANDX1 G29249 (.A1(W17530), .A2(W17192), .ZN(W17903));
  NANDX1 G29250 (.A1(I151), .A2(W3376), .ZN(W5121));
  NANDX1 G29251 (.A1(W4086), .A2(W5448), .ZN(W7836));
  NANDX1 G29252 (.A1(W1276), .A2(W3726), .ZN(W17847));
  NANDX1 G29253 (.A1(W3936), .A2(W5131), .ZN(W13690));
  NANDX1 G29254 (.A1(W5611), .A2(W9020), .ZN(W13694));
  NANDX1 G29255 (.A1(I393), .A2(W7509), .ZN(O1455));
  NANDX1 G29256 (.A1(W6481), .A2(W6673), .ZN(W13695));
  NANDX1 G29257 (.A1(W1587), .A2(W3388), .ZN(W5157));
  NANDX1 G29258 (.A1(W10430), .A2(W15349), .ZN(W17850));
  NANDX1 G29259 (.A1(W9971), .A2(W3678), .ZN(W17849));
  NANDX1 G29260 (.A1(W12837), .A2(W16477), .ZN(W17848));
  NANDX1 G29261 (.A1(I1336), .A2(W884), .ZN(W5153));
  NANDX1 G29262 (.A1(W11383), .A2(W10806), .ZN(W17846));
  NANDX1 G29263 (.A1(W2920), .A2(W15803), .ZN(W17845));
  NANDX1 G29264 (.A1(W13979), .A2(I291), .ZN(O1454));
  NANDX1 G29265 (.A1(W8885), .A2(W1011), .ZN(O1453));
  NANDX1 G29266 (.A1(W2293), .A2(W230), .ZN(W5160));
  NANDX1 G29267 (.A1(W8161), .A2(W11348), .ZN(O777));
  NANDX1 G29268 (.A1(I1400), .A2(W12949), .ZN(W13705));
  NANDX1 G29269 (.A1(W6247), .A2(W4524), .ZN(W17841));
  NANDX1 G29270 (.A1(W14894), .A2(W8158), .ZN(W17866));
  NANDX1 G29271 (.A1(W10581), .A2(I1392), .ZN(W17873));
  NANDX1 G29272 (.A1(W1780), .A2(I20), .ZN(W5136));
  NANDX1 G29273 (.A1(I1084), .A2(I1036), .ZN(W5137));
  NANDX1 G29274 (.A1(W5031), .A2(W1236), .ZN(W7831));
  NANDX1 G29275 (.A1(W4078), .A2(W14026), .ZN(W17870));
  NANDX1 G29276 (.A1(W7241), .A2(W2505), .ZN(O1458));
  NANDX1 G29277 (.A1(W5668), .A2(W9275), .ZN(W17867));
  NANDX1 G29278 (.A1(W8875), .A2(W8094), .ZN(W13684));
  NANDX1 G29279 (.A1(W16142), .A2(W14232), .ZN(W17738));
  NANDX1 G29280 (.A1(I1358), .A2(W12286), .ZN(W17865));
  NANDX1 G29281 (.A1(W17422), .A2(W9868), .ZN(W17863));
  NANDX1 G29282 (.A1(I1712), .A2(W12134), .ZN(O776));
  NANDX1 G29283 (.A1(W15311), .A2(W16929), .ZN(W17857));
  NANDX1 G29284 (.A1(W4512), .A2(W242), .ZN(W7829));
  NANDX1 G29285 (.A1(I1642), .A2(W2327), .ZN(W5148));
  NANDX1 G29286 (.A1(W10326), .A2(W10773), .ZN(W13689));
  NANDX1 G29287 (.A1(W5902), .A2(W304), .ZN(W17855));
  NANDX1 G29288 (.A1(W4892), .A2(W673), .ZN(W5296));
  NANDX1 G29289 (.A1(W980), .A2(I870), .ZN(W7738));
  NANDX1 G29290 (.A1(I1941), .A2(W1592), .ZN(W5287));
  NANDX1 G29291 (.A1(W1625), .A2(W16234), .ZN(W17641));
  NANDX1 G29292 (.A1(W3174), .A2(W385), .ZN(W5290));
  NANDX1 G29293 (.A1(W5480), .A2(W16240), .ZN(W17640));
  NANDX1 G29294 (.A1(W1078), .A2(W4771), .ZN(W5291));
  NANDX1 G29295 (.A1(W2572), .A2(I956), .ZN(W5293));
  NANDX1 G29296 (.A1(W15532), .A2(W16592), .ZN(W17636));
  NANDX1 G29297 (.A1(I271), .A2(W355), .ZN(W5294));
  NANDX1 G29298 (.A1(W2112), .A2(W1014), .ZN(W5285));
  NANDX1 G29299 (.A1(W7351), .A2(W6136), .ZN(W17631));
  NANDX1 G29300 (.A1(W3582), .A2(W6863), .ZN(W7737));
  NANDX1 G29301 (.A1(W10174), .A2(W14862), .ZN(W17628));
  NANDX1 G29302 (.A1(I1784), .A2(W5317), .ZN(O198));
  NANDX1 G29303 (.A1(W9742), .A2(W5383), .ZN(W17626));
  NANDX1 G29304 (.A1(W2261), .A2(W3073), .ZN(W7733));
  NANDX1 G29305 (.A1(W3804), .A2(I1482), .ZN(W5302));
  NANDX1 G29306 (.A1(W1822), .A2(W3602), .ZN(W13813));
  NANDX1 G29307 (.A1(W2386), .A2(W140), .ZN(W5273));
  NANDX1 G29308 (.A1(W539), .A2(W2806), .ZN(W7755));
  NANDX1 G29309 (.A1(I1695), .A2(W4313), .ZN(W5265));
  NANDX1 G29310 (.A1(W1395), .A2(W8857), .ZN(O1423));
  NANDX1 G29311 (.A1(W15827), .A2(W4589), .ZN(W17653));
  NANDX1 G29312 (.A1(W1441), .A2(W2185), .ZN(W5268));
  NANDX1 G29313 (.A1(W16565), .A2(W13940), .ZN(W17651));
  NANDX1 G29314 (.A1(W2124), .A2(W4826), .ZN(W5271));
  NANDX1 G29315 (.A1(W3254), .A2(W7235), .ZN(W7752));
  NANDX1 G29316 (.A1(W3789), .A2(W16128), .ZN(W17621));
  NANDX1 G29317 (.A1(W3341), .A2(W7744), .ZN(W7748));
  NANDX1 G29318 (.A1(W3456), .A2(W1155), .ZN(W5279));
  NANDX1 G29319 (.A1(W7408), .A2(I1368), .ZN(W7747));
  NANDX1 G29320 (.A1(I812), .A2(I1960), .ZN(O80));
  NANDX1 G29321 (.A1(W4793), .A2(W4770), .ZN(W5283));
  NANDX1 G29322 (.A1(W2057), .A2(W5784), .ZN(W7746));
  NANDX1 G29323 (.A1(I134), .A2(W7732), .ZN(O199));
  NANDX1 G29324 (.A1(W3380), .A2(W2016), .ZN(W5284));
  NANDX1 G29325 (.A1(W7439), .A2(W10427), .ZN(W17580));
  NANDX1 G29326 (.A1(W4983), .A2(I519), .ZN(W17589));
  NANDX1 G29327 (.A1(W8134), .A2(I1161), .ZN(W13832));
  NANDX1 G29328 (.A1(I1876), .A2(W2118), .ZN(W5316));
  NANDX1 G29329 (.A1(W16441), .A2(W7622), .ZN(W17587));
  NANDX1 G29330 (.A1(I565), .A2(I1591), .ZN(O81));
  NANDX1 G29331 (.A1(W13300), .A2(W8827), .ZN(W17584));
  NANDX1 G29332 (.A1(I1336), .A2(W13489), .ZN(W17583));
  NANDX1 G29333 (.A1(W1473), .A2(I1324), .ZN(W7722));
  NANDX1 G29334 (.A1(W4885), .A2(W5153), .ZN(W7723));
  NANDX1 G29335 (.A1(W11373), .A2(W8042), .ZN(W17579));
  NANDX1 G29336 (.A1(W9537), .A2(W12138), .ZN(W17578));
  NANDX1 G29337 (.A1(I385), .A2(I1824), .ZN(W5326));
  NANDX1 G29338 (.A1(W12721), .A2(W14169), .ZN(W17575));
  NANDX1 G29339 (.A1(W51), .A2(I1472), .ZN(W5327));
  NANDX1 G29340 (.A1(W11512), .A2(W17498), .ZN(W17572));
  NANDX1 G29341 (.A1(W11839), .A2(W4279), .ZN(W17571));
  NANDX1 G29342 (.A1(W8235), .A2(W2315), .ZN(W17568));
  NANDX1 G29343 (.A1(W14875), .A2(W11126), .ZN(W17601));
  NANDX1 G29344 (.A1(W3625), .A2(W821), .ZN(W13814));
  NANDX1 G29345 (.A1(I696), .A2(W2624), .ZN(W17615));
  NANDX1 G29346 (.A1(I494), .A2(W5591), .ZN(W17614));
  NANDX1 G29347 (.A1(W14174), .A2(W4007), .ZN(W17613));
  NANDX1 G29348 (.A1(I1173), .A2(W3003), .ZN(O197));
  NANDX1 G29349 (.A1(W16966), .A2(W4524), .ZN(W17607));
  NANDX1 G29350 (.A1(W11778), .A2(W17211), .ZN(W17606));
  NANDX1 G29351 (.A1(W3240), .A2(I782), .ZN(W5306));
  NANDX1 G29352 (.A1(W57), .A2(W5252), .ZN(W5262));
  NANDX1 G29353 (.A1(W11144), .A2(W3189), .ZN(O1414));
  NANDX1 G29354 (.A1(W847), .A2(W187), .ZN(W13818));
  NANDX1 G29355 (.A1(W5777), .A2(W717), .ZN(W13820));
  NANDX1 G29356 (.A1(I1579), .A2(W7331), .ZN(W7726));
  NANDX1 G29357 (.A1(W15721), .A2(W1998), .ZN(W17595));
  NANDX1 G29358 (.A1(I598), .A2(W4821), .ZN(W5313));
  NANDX1 G29359 (.A1(W5110), .A2(W2912), .ZN(W5314));
  NANDX1 G29360 (.A1(W512), .A2(W1161), .ZN(W13827));
  NANDX1 G29361 (.A1(W332), .A2(W4272), .ZN(W7776));
  NANDX1 G29362 (.A1(W3835), .A2(W4296), .ZN(W17716));
  NANDX1 G29363 (.A1(W6762), .A2(W4487), .ZN(W13758));
  NANDX1 G29364 (.A1(W6471), .A2(W13329), .ZN(W17712));
  NANDX1 G29365 (.A1(W11610), .A2(W1378), .ZN(W13759));
  NANDX1 G29366 (.A1(W5908), .A2(W13907), .ZN(W17709));
  NANDX1 G29367 (.A1(W4519), .A2(W4225), .ZN(W7778));
  NANDX1 G29368 (.A1(I1398), .A2(W569), .ZN(W17708));
  NANDX1 G29369 (.A1(W49), .A2(W4704), .ZN(W5228));
  NANDX1 G29370 (.A1(W2402), .A2(W1968), .ZN(W5229));
  NANDX1 G29371 (.A1(W1814), .A2(W5081), .ZN(W7780));
  NANDX1 G29372 (.A1(W4601), .A2(I1492), .ZN(W5232));
  NANDX1 G29373 (.A1(W7061), .A2(I481), .ZN(W17701));
  NANDX1 G29374 (.A1(I1894), .A2(W4247), .ZN(W5234));
  NANDX1 G29375 (.A1(I909), .A2(W437), .ZN(W5236));
  NANDX1 G29376 (.A1(W16436), .A2(I964), .ZN(W17697));
  NANDX1 G29377 (.A1(W17594), .A2(W12093), .ZN(W17694));
  NANDX1 G29378 (.A1(W6639), .A2(W488), .ZN(O200));
  NANDX1 G29379 (.A1(W2920), .A2(W16664), .ZN(W17693));
  NANDX1 G29380 (.A1(W4410), .A2(W2150), .ZN(W7788));
  NANDX1 G29381 (.A1(I707), .A2(W6272), .ZN(W7791));
  NANDX1 G29382 (.A1(W9030), .A2(W6207), .ZN(W17736));
  NANDX1 G29383 (.A1(W3964), .A2(W7383), .ZN(W7789));
  NANDX1 G29384 (.A1(W11573), .A2(W2370), .ZN(W17732));
  NANDX1 G29385 (.A1(W9613), .A2(W15868), .ZN(W17730));
  NANDX1 G29386 (.A1(W9454), .A2(W1486), .ZN(W17728));
  NANDX1 G29387 (.A1(W1965), .A2(W12384), .ZN(W17727));
  NANDX1 G29388 (.A1(W1999), .A2(W10006), .ZN(W13750));
  NANDX1 G29389 (.A1(W8753), .A2(W12353), .ZN(O1433));
  NANDX1 G29390 (.A1(I472), .A2(W3476), .ZN(W5216));
  NANDX1 G29391 (.A1(I874), .A2(W6241), .ZN(W7786));
  NANDX1 G29392 (.A1(I1614), .A2(W7554), .ZN(W7785));
  NANDX1 G29393 (.A1(W205), .A2(W6869), .ZN(W7784));
  NANDX1 G29394 (.A1(W2063), .A2(W7275), .ZN(W7782));
  NANDX1 G29395 (.A1(W5123), .A2(W4816), .ZN(W5220));
  NANDX1 G29396 (.A1(W1075), .A2(W6708), .ZN(W7781));
  NANDX1 G29397 (.A1(W3062), .A2(W3144), .ZN(W5221));
  NANDX1 G29398 (.A1(W2495), .A2(W6464), .ZN(W17668));
  NANDX1 G29399 (.A1(W9948), .A2(I975), .ZN(W17674));
  NANDX1 G29400 (.A1(W6126), .A2(W2230), .ZN(W7761));
  NANDX1 G29401 (.A1(W3232), .A2(W6786), .ZN(W7759));
  NANDX1 G29402 (.A1(W1646), .A2(W1789), .ZN(W5255));
  NANDX1 G29403 (.A1(I930), .A2(W9421), .ZN(W13784));
  NANDX1 G29404 (.A1(W7152), .A2(W12289), .ZN(W17672));
  NANDX1 G29405 (.A1(W4837), .A2(W1687), .ZN(W17671));
  NANDX1 G29406 (.A1(W13245), .A2(W10335), .ZN(O1427));
  NANDX1 G29407 (.A1(W10929), .A2(W11580), .ZN(O1429));
  NANDX1 G29408 (.A1(W1075), .A2(W4971), .ZN(W5256));
  NANDX1 G29409 (.A1(I1298), .A2(I1367), .ZN(W5257));
  NANDX1 G29410 (.A1(W15218), .A2(W9056), .ZN(W17665));
  NANDX1 G29411 (.A1(I1153), .A2(W7351), .ZN(W13791));
  NANDX1 G29412 (.A1(W9258), .A2(I250), .ZN(W17663));
  NANDX1 G29413 (.A1(W7758), .A2(W13131), .ZN(W17661));
  NANDX1 G29414 (.A1(W2603), .A2(W2638), .ZN(W5260));
  NANDX1 G29415 (.A1(I705), .A2(W779), .ZN(W5261));
  NANDX1 G29416 (.A1(I514), .A2(W15474), .ZN(W17681));
  NANDX1 G29417 (.A1(W1328), .A2(W14318), .ZN(W17691));
  NANDX1 G29418 (.A1(W7752), .A2(W12322), .ZN(W17690));
  NANDX1 G29419 (.A1(W2530), .A2(W11528), .ZN(W13770));
  NANDX1 G29420 (.A1(W16516), .A2(W10453), .ZN(W17688));
  NANDX1 G29421 (.A1(I503), .A2(W5338), .ZN(W13771));
  NANDX1 G29422 (.A1(W4502), .A2(W9748), .ZN(W17685));
  NANDX1 G29423 (.A1(I186), .A2(I1675), .ZN(W13774));
  NANDX1 G29424 (.A1(W1188), .A2(W3160), .ZN(W7764));
  NANDX1 G29425 (.A1(W2479), .A2(W614), .ZN(W13983));
  NANDX1 G29426 (.A1(W7125), .A2(W1527), .ZN(W7763));
  NANDX1 G29427 (.A1(W11633), .A2(W12264), .ZN(W17680));
  NANDX1 G29428 (.A1(W475), .A2(W3708), .ZN(W5242));
  NANDX1 G29429 (.A1(W16819), .A2(W6967), .ZN(W17679));
  NANDX1 G29430 (.A1(W13641), .A2(W577), .ZN(W13777));
  NANDX1 G29431 (.A1(W5168), .A2(W7906), .ZN(W13778));
  NANDX1 G29432 (.A1(W1529), .A2(W4061), .ZN(W5245));
  NANDX1 G29433 (.A1(W619), .A2(W2194), .ZN(W17677));
  NANDX1 G29434 (.A1(W7353), .A2(W4152), .ZN(W16705));
  NANDX1 G29435 (.A1(W2361), .A2(I856), .ZN(W5890));
  NANDX1 G29436 (.A1(W4814), .A2(W4745), .ZN(W5894));
  NANDX1 G29437 (.A1(W4387), .A2(W11290), .ZN(W16716));
  NANDX1 G29438 (.A1(I1036), .A2(W4608), .ZN(W5895));
  NANDX1 G29439 (.A1(W1965), .A2(W9490), .ZN(W16715));
  NANDX1 G29440 (.A1(W4973), .A2(W4731), .ZN(W16713));
  NANDX1 G29441 (.A1(W3633), .A2(W13562), .ZN(O1234));
  NANDX1 G29442 (.A1(I109), .A2(W8546), .ZN(W16710));
  NANDX1 G29443 (.A1(W3500), .A2(W5468), .ZN(W7462));
  NANDX1 G29444 (.A1(W4512), .A2(W2062), .ZN(W14207));
  NANDX1 G29445 (.A1(W13768), .A2(I1305), .ZN(W14210));
  NANDX1 G29446 (.A1(I679), .A2(W1941), .ZN(W7459));
  NANDX1 G29447 (.A1(W13290), .A2(W7030), .ZN(W16704));
  NANDX1 G29448 (.A1(W9093), .A2(W8730), .ZN(W16703));
  NANDX1 G29449 (.A1(W13323), .A2(I310), .ZN(W14216));
  NANDX1 G29450 (.A1(W7837), .A2(W4838), .ZN(W16699));
  NANDX1 G29451 (.A1(W15598), .A2(W11689), .ZN(W16698));
  NANDX1 G29452 (.A1(W3735), .A2(W4676), .ZN(W7455));
  NANDX1 G29453 (.A1(W4096), .A2(W11575), .ZN(W14206));
  NANDX1 G29454 (.A1(W14501), .A2(W12019), .ZN(O1244));
  NANDX1 G29455 (.A1(I876), .A2(W10933), .ZN(W14200));
  NANDX1 G29456 (.A1(W1827), .A2(W2440), .ZN(W7468));
  NANDX1 G29457 (.A1(I1794), .A2(W3405), .ZN(W5879));
  NANDX1 G29458 (.A1(W5577), .A2(W4002), .ZN(W14202));
  NANDX1 G29459 (.A1(I1664), .A2(W9212), .ZN(W16735));
  NANDX1 G29460 (.A1(W6475), .A2(W5066), .ZN(O1243));
  NANDX1 G29461 (.A1(W1553), .A2(W5246), .ZN(W5880));
  NANDX1 G29462 (.A1(W3295), .A2(W12133), .ZN(W14219));
  NANDX1 G29463 (.A1(W5865), .A2(W13205), .ZN(W16733));
  NANDX1 G29464 (.A1(W13122), .A2(W12392), .ZN(O1242));
  NANDX1 G29465 (.A1(W3380), .A2(W4768), .ZN(W5883));
  NANDX1 G29466 (.A1(W2854), .A2(W2417), .ZN(W5884));
  NANDX1 G29467 (.A1(W2243), .A2(W426), .ZN(W5885));
  NANDX1 G29468 (.A1(W4694), .A2(I1782), .ZN(W5886));
  NANDX1 G29469 (.A1(W6661), .A2(W4679), .ZN(W7466));
  NANDX1 G29470 (.A1(W4597), .A2(W16671), .ZN(W16724));
  NANDX1 G29471 (.A1(W2512), .A2(I354), .ZN(W5922));
  NANDX1 G29472 (.A1(W1361), .A2(W1762), .ZN(W7450));
  NANDX1 G29473 (.A1(I18), .A2(W13083), .ZN(O1226));
  NANDX1 G29474 (.A1(W924), .A2(I316), .ZN(W5917));
  NANDX1 G29475 (.A1(W5735), .A2(W1370), .ZN(O846));
  NANDX1 G29476 (.A1(I26), .A2(W6744), .ZN(O847));
  NANDX1 G29477 (.A1(W3407), .A2(W999), .ZN(W5921));
  NANDX1 G29478 (.A1(W3872), .A2(W1904), .ZN(O1224));
  NANDX1 G29479 (.A1(I191), .A2(W12594), .ZN(W14232));
  NANDX1 G29480 (.A1(W1584), .A2(W456), .ZN(W5914));
  NANDX1 G29481 (.A1(I856), .A2(W1562), .ZN(W5924));
  NANDX1 G29482 (.A1(W12757), .A2(W2260), .ZN(W16659));
  NANDX1 G29483 (.A1(W3323), .A2(W5358), .ZN(W14234));
  NANDX1 G29484 (.A1(I606), .A2(W4051), .ZN(W5926));
  NANDX1 G29485 (.A1(W2299), .A2(W5342), .ZN(O107));
  NANDX1 G29486 (.A1(W532), .A2(I1412), .ZN(W5930));
  NANDX1 G29487 (.A1(W4335), .A2(I1304), .ZN(W5931));
  NANDX1 G29488 (.A1(I1080), .A2(I202), .ZN(W7448));
  NANDX1 G29489 (.A1(I831), .A2(I575), .ZN(W16689));
  NANDX1 G29490 (.A1(W3580), .A2(I1385), .ZN(W16696));
  NANDX1 G29491 (.A1(W3026), .A2(W5856), .ZN(W5902));
  NANDX1 G29492 (.A1(W12649), .A2(W6117), .ZN(W14220));
  NANDX1 G29493 (.A1(W12958), .A2(W10394), .ZN(O843));
  NANDX1 G29494 (.A1(W770), .A2(W3776), .ZN(W5906));
  NANDX1 G29495 (.A1(W7298), .A2(W3516), .ZN(W7453));
  NANDX1 G29496 (.A1(W6722), .A2(W587), .ZN(W7452));
  NANDX1 G29497 (.A1(W6188), .A2(I1132), .ZN(W16690));
  NANDX1 G29498 (.A1(W3674), .A2(W783), .ZN(W7469));
  NANDX1 G29499 (.A1(W1278), .A2(W4162), .ZN(W5908));
  NANDX1 G29500 (.A1(W1882), .A2(W4420), .ZN(W5910));
  NANDX1 G29501 (.A1(W14050), .A2(W2800), .ZN(W14225));
  NANDX1 G29502 (.A1(W12498), .A2(I1883), .ZN(W14227));
  NANDX1 G29503 (.A1(W1341), .A2(W6761), .ZN(O1227));
  NANDX1 G29504 (.A1(W4279), .A2(W5088), .ZN(W5913));
  NANDX1 G29505 (.A1(W3135), .A2(W4227), .ZN(W16680));
  NANDX1 G29506 (.A1(W2432), .A2(W399), .ZN(W16679));
  NANDX1 G29507 (.A1(W12475), .A2(W15476), .ZN(W16807));
  NANDX1 G29508 (.A1(I787), .A2(W5566), .ZN(W5826));
  NANDX1 G29509 (.A1(W623), .A2(W438), .ZN(W7499));
  NANDX1 G29510 (.A1(W3861), .A2(I1055), .ZN(W5828));
  NANDX1 G29511 (.A1(W2884), .A2(W4998), .ZN(W5829));
  NANDX1 G29512 (.A1(W9258), .A2(W7050), .ZN(W16814));
  NANDX1 G29513 (.A1(W12444), .A2(W3836), .ZN(W16813));
  NANDX1 G29514 (.A1(W9701), .A2(W6297), .ZN(W14165));
  NANDX1 G29515 (.A1(W15703), .A2(W15829), .ZN(W16810));
  NANDX1 G29516 (.A1(W12377), .A2(W5539), .ZN(W14167));
  NANDX1 G29517 (.A1(W3940), .A2(W3548), .ZN(W14161));
  NANDX1 G29518 (.A1(W1865), .A2(W4246), .ZN(O105));
  NANDX1 G29519 (.A1(W8004), .A2(W13620), .ZN(W16806));
  NANDX1 G29520 (.A1(W9493), .A2(I457), .ZN(W14168));
  NANDX1 G29521 (.A1(I370), .A2(W2093), .ZN(W5837));
  NANDX1 G29522 (.A1(W3579), .A2(W16568), .ZN(O1267));
  NANDX1 G29523 (.A1(W4302), .A2(W880), .ZN(W16800));
  NANDX1 G29524 (.A1(W4565), .A2(W4432), .ZN(W5846));
  NANDX1 G29525 (.A1(W4805), .A2(W9997), .ZN(W14170));
  NANDX1 G29526 (.A1(I738), .A2(W4738), .ZN(W5815));
  NANDX1 G29527 (.A1(W11021), .A2(W4165), .ZN(W14154));
  NANDX1 G29528 (.A1(W7127), .A2(W15217), .ZN(W16841));
  NANDX1 G29529 (.A1(W3727), .A2(W3384), .ZN(W16840));
  NANDX1 G29530 (.A1(I1186), .A2(W5380), .ZN(W16839));
  NANDX1 G29531 (.A1(W8680), .A2(W1317), .ZN(W16838));
  NANDX1 G29532 (.A1(W3247), .A2(W1674), .ZN(W5812));
  NANDX1 G29533 (.A1(W2066), .A2(W6670), .ZN(W14155));
  NANDX1 G29534 (.A1(W11716), .A2(W3990), .ZN(W16836));
  NANDX1 G29535 (.A1(W8065), .A2(W1274), .ZN(O1262));
  NANDX1 G29536 (.A1(I678), .A2(I178), .ZN(W16833));
  NANDX1 G29537 (.A1(W3314), .A2(W886), .ZN(W5818));
  NANDX1 G29538 (.A1(W1984), .A2(W751), .ZN(W16827));
  NANDX1 G29539 (.A1(I1483), .A2(W12570), .ZN(W16826));
  NANDX1 G29540 (.A1(W5319), .A2(I1375), .ZN(W5819));
  NANDX1 G29541 (.A1(W12789), .A2(W358), .ZN(O1269));
  NANDX1 G29542 (.A1(W12756), .A2(W16610), .ZN(W16821));
  NANDX1 G29543 (.A1(I1442), .A2(I1895), .ZN(W5821));
  NANDX1 G29544 (.A1(W4031), .A2(W1318), .ZN(W5870));
  NANDX1 G29545 (.A1(W1135), .A2(W1450), .ZN(W5861));
  NANDX1 G29546 (.A1(W3927), .A2(W5327), .ZN(W5862));
  NANDX1 G29547 (.A1(W2680), .A2(W86), .ZN(W5863));
  NANDX1 G29548 (.A1(W11803), .A2(W10793), .ZN(W16759));
  NANDX1 G29549 (.A1(W698), .A2(W9138), .ZN(W16755));
  NANDX1 G29550 (.A1(W185), .A2(W12418), .ZN(O836));
  NANDX1 G29551 (.A1(W2255), .A2(W5849), .ZN(W5869));
  NANDX1 G29552 (.A1(W7249), .A2(W7687), .ZN(O1250));
  NANDX1 G29553 (.A1(W10367), .A2(W11020), .ZN(W16764));
  NANDX1 G29554 (.A1(W11837), .A2(W14178), .ZN(O1249));
  NANDX1 G29555 (.A1(I1072), .A2(W14808), .ZN(O1248));
  NANDX1 G29556 (.A1(W12612), .A2(W11979), .ZN(W16746));
  NANDX1 G29557 (.A1(W7102), .A2(W1613), .ZN(W14184));
  NANDX1 G29558 (.A1(W6784), .A2(W10738), .ZN(O837));
  NANDX1 G29559 (.A1(W6929), .A2(W12441), .ZN(W14186));
  NANDX1 G29560 (.A1(I1372), .A2(W11387), .ZN(W14187));
  NANDX1 G29561 (.A1(W5709), .A2(W2428), .ZN(W14196));
  NANDX1 G29562 (.A1(I95), .A2(I1918), .ZN(W7485));
  NANDX1 G29563 (.A1(W2357), .A2(W5003), .ZN(W5851));
  NANDX1 G29564 (.A1(I1773), .A2(W7969), .ZN(W16792));
  NANDX1 G29565 (.A1(W4268), .A2(W1649), .ZN(W5852));
  NANDX1 G29566 (.A1(W8177), .A2(W11028), .ZN(W16791));
  NANDX1 G29567 (.A1(W6115), .A2(W5632), .ZN(W16783));
  NANDX1 G29568 (.A1(W1968), .A2(W4908), .ZN(W7488));
  NANDX1 G29569 (.A1(W5293), .A2(W3382), .ZN(W5856));
  NANDX1 G29570 (.A1(W1985), .A2(I441), .ZN(W7487));
  NANDX1 G29571 (.A1(W5751), .A2(W1026), .ZN(W5935));
  NANDX1 G29572 (.A1(W5505), .A2(W4784), .ZN(W5858));
  NANDX1 G29573 (.A1(W8191), .A2(W15166), .ZN(W16776));
  NANDX1 G29574 (.A1(W367), .A2(W9637), .ZN(W16775));
  NANDX1 G29575 (.A1(W12940), .A2(W11952), .ZN(O835));
  NANDX1 G29576 (.A1(W10339), .A2(W7485), .ZN(O1257));
  NANDX1 G29577 (.A1(W16186), .A2(W12282), .ZN(W16770));
  NANDX1 G29578 (.A1(W15588), .A2(W9447), .ZN(W16766));
  NANDX1 G29579 (.A1(W4737), .A2(W12762), .ZN(O1255));
  NANDX1 G29580 (.A1(W1156), .A2(W1763), .ZN(W6022));
  NANDX1 G29581 (.A1(W7320), .A2(W15116), .ZN(W16526));
  NANDX1 G29582 (.A1(W12247), .A2(W11437), .ZN(O1192));
  NANDX1 G29583 (.A1(W7179), .A2(W13426), .ZN(W14288));
  NANDX1 G29584 (.A1(I858), .A2(W11178), .ZN(O851));
  NANDX1 G29585 (.A1(W5029), .A2(W4607), .ZN(W6019));
  NANDX1 G29586 (.A1(W15550), .A2(I1637), .ZN(W16520));
  NANDX1 G29587 (.A1(I1431), .A2(I1532), .ZN(W7414));
  NANDX1 G29588 (.A1(W8748), .A2(W12637), .ZN(W16516));
  NANDX1 G29589 (.A1(I1105), .A2(W1226), .ZN(W6021));
  NANDX1 G29590 (.A1(W14711), .A2(W14876), .ZN(W16528));
  NANDX1 G29591 (.A1(W2017), .A2(W4375), .ZN(W6023));
  NANDX1 G29592 (.A1(W12029), .A2(W4755), .ZN(W16512));
  NANDX1 G29593 (.A1(W3925), .A2(W11774), .ZN(W14291));
  NANDX1 G29594 (.A1(W6029), .A2(W13983), .ZN(W14294));
  NANDX1 G29595 (.A1(W4750), .A2(I1788), .ZN(O1189));
  NANDX1 G29596 (.A1(I1050), .A2(W11763), .ZN(O1188));
  NANDX1 G29597 (.A1(W96), .A2(I460), .ZN(W6026));
  NANDX1 G29598 (.A1(I9), .A2(I547), .ZN(W6028));
  NANDX1 G29599 (.A1(W13690), .A2(W10858), .ZN(O849));
  NANDX1 G29600 (.A1(W2035), .A2(I31), .ZN(O1202));
  NANDX1 G29601 (.A1(W8554), .A2(W733), .ZN(W16555));
  NANDX1 G29602 (.A1(W15821), .A2(W16183), .ZN(O1200));
  NANDX1 G29603 (.A1(I1524), .A2(W2076), .ZN(W6006));
  NANDX1 G29604 (.A1(W5115), .A2(W1838), .ZN(W16549));
  NANDX1 G29605 (.A1(W3946), .A2(W5857), .ZN(W6010));
  NANDX1 G29606 (.A1(W1093), .A2(W3833), .ZN(W6011));
  NANDX1 G29607 (.A1(W6305), .A2(W4436), .ZN(W16545));
  NANDX1 G29608 (.A1(I1120), .A2(I626), .ZN(W6029));
  NANDX1 G29609 (.A1(W14398), .A2(W4325), .ZN(O1197));
  NANDX1 G29610 (.A1(W3508), .A2(I138), .ZN(W6012));
  NANDX1 G29611 (.A1(W3236), .A2(W2001), .ZN(W6013));
  NANDX1 G29612 (.A1(W2791), .A2(W6351), .ZN(O1195));
  NANDX1 G29613 (.A1(W15564), .A2(W2705), .ZN(O1194));
  NANDX1 G29614 (.A1(W1542), .A2(W8429), .ZN(W16532));
  NANDX1 G29615 (.A1(W54), .A2(W5196), .ZN(W6015));
  NANDX1 G29616 (.A1(I1535), .A2(W4662), .ZN(O181));
  NANDX1 G29617 (.A1(W8892), .A2(I660), .ZN(W16469));
  NANDX1 G29618 (.A1(I1472), .A2(W6625), .ZN(W14299));
  NANDX1 G29619 (.A1(W11105), .A2(W6517), .ZN(O1183));
  NANDX1 G29620 (.A1(W15078), .A2(W7880), .ZN(W16479));
  NANDX1 G29621 (.A1(W5966), .A2(W8541), .ZN(W14300));
  NANDX1 G29622 (.A1(W5100), .A2(I1133), .ZN(W7403));
  NANDX1 G29623 (.A1(W11903), .A2(W6563), .ZN(W16473));
  NANDX1 G29624 (.A1(W5159), .A2(W1650), .ZN(W6045));
  NANDX1 G29625 (.A1(W2652), .A2(W9953), .ZN(W16470));
  NANDX1 G29626 (.A1(W5404), .A2(W821), .ZN(W7404));
  NANDX1 G29627 (.A1(W13854), .A2(W5970), .ZN(W16468));
  NANDX1 G29628 (.A1(W8763), .A2(W9897), .ZN(W16463));
  NANDX1 G29629 (.A1(W8196), .A2(W1125), .ZN(W16461));
  NANDX1 G29630 (.A1(W12680), .A2(W6458), .ZN(W14302));
  NANDX1 G29631 (.A1(W14641), .A2(W9869), .ZN(W16458));
  NANDX1 G29632 (.A1(W12187), .A2(W4915), .ZN(W16454));
  NANDX1 G29633 (.A1(W3444), .A2(W3663), .ZN(W6048));
  NANDX1 G29634 (.A1(I638), .A2(W3913), .ZN(W6049));
  NANDX1 G29635 (.A1(W350), .A2(I920), .ZN(W6036));
  NANDX1 G29636 (.A1(W5263), .A2(W7316), .ZN(W7410));
  NANDX1 G29637 (.A1(W16127), .A2(W6946), .ZN(W16503));
  NANDX1 G29638 (.A1(W13719), .A2(W13834), .ZN(W16502));
  NANDX1 G29639 (.A1(W3873), .A2(W5266), .ZN(W7409));
  NANDX1 G29640 (.A1(W14962), .A2(W12802), .ZN(W16500));
  NANDX1 G29641 (.A1(W13546), .A2(W10976), .ZN(W14297));
  NANDX1 G29642 (.A1(W742), .A2(W4451), .ZN(W6035));
  NANDX1 G29643 (.A1(W6324), .A2(W3768), .ZN(W16497));
  NANDX1 G29644 (.A1(W7325), .A2(W15623), .ZN(O1203));
  NANDX1 G29645 (.A1(W6136), .A2(W5826), .ZN(W7406));
  NANDX1 G29646 (.A1(W3271), .A2(W565), .ZN(W16496));
  NANDX1 G29647 (.A1(I17), .A2(W1255), .ZN(W6039));
  NANDX1 G29648 (.A1(W4550), .A2(W7291), .ZN(W16489));
  NANDX1 G29649 (.A1(W3654), .A2(W5880), .ZN(W16488));
  NANDX1 G29650 (.A1(W2786), .A2(W627), .ZN(W6040));
  NANDX1 G29651 (.A1(W5573), .A2(W1021), .ZN(W6041));
  NANDX1 G29652 (.A1(W11403), .A2(W10648), .ZN(W16484));
  NANDX1 G29653 (.A1(W11290), .A2(I1846), .ZN(W16609));
  NANDX1 G29654 (.A1(I1350), .A2(W3248), .ZN(W5954));
  NANDX1 G29655 (.A1(W5526), .A2(W13633), .ZN(W16619));
  NANDX1 G29656 (.A1(W4669), .A2(W2171), .ZN(W5955));
  NANDX1 G29657 (.A1(W10627), .A2(W10741), .ZN(W16617));
  NANDX1 G29658 (.A1(W7961), .A2(W10579), .ZN(W16616));
  NANDX1 G29659 (.A1(W1341), .A2(W2196), .ZN(W5956));
  NANDX1 G29660 (.A1(W3007), .A2(W10797), .ZN(O848));
  NANDX1 G29661 (.A1(W14830), .A2(W9836), .ZN(W16611));
  NANDX1 G29662 (.A1(W16232), .A2(W11655), .ZN(W16610));
  NANDX1 G29663 (.A1(W7049), .A2(W7054), .ZN(W7438));
  NANDX1 G29664 (.A1(W3989), .A2(W2391), .ZN(W5957));
  NANDX1 G29665 (.A1(W1136), .A2(W6640), .ZN(W7436));
  NANDX1 G29666 (.A1(W6227), .A2(W2205), .ZN(W14256));
  NANDX1 G29667 (.A1(I946), .A2(W2904), .ZN(W7433));
  NANDX1 G29668 (.A1(W7915), .A2(W6380), .ZN(W14258));
  NANDX1 G29669 (.A1(W9633), .A2(W9260), .ZN(W14259));
  NANDX1 G29670 (.A1(W5960), .A2(W3319), .ZN(O109));
  NANDX1 G29671 (.A1(W6278), .A2(W12046), .ZN(W14261));
  NANDX1 G29672 (.A1(W6232), .A2(W770), .ZN(O1218));
  NANDX1 G29673 (.A1(W4024), .A2(W5430), .ZN(W5937));
  NANDX1 G29674 (.A1(W9736), .A2(W7315), .ZN(W14239));
  NANDX1 G29675 (.A1(W13885), .A2(W9946), .ZN(W16642));
  NANDX1 G29676 (.A1(W5378), .A2(W2930), .ZN(W7445));
  NANDX1 G29677 (.A1(I909), .A2(W13202), .ZN(W16640));
  NANDX1 G29678 (.A1(W435), .A2(W482), .ZN(W14244));
  NANDX1 G29679 (.A1(W1552), .A2(W541), .ZN(W5944));
  NANDX1 G29680 (.A1(W10583), .A2(W9630), .ZN(W16638));
  NANDX1 G29681 (.A1(W13882), .A2(I1706), .ZN(W16604));
  NANDX1 G29682 (.A1(W7279), .A2(W3386), .ZN(W14246));
  NANDX1 G29683 (.A1(W1061), .A2(W4080), .ZN(W5946));
  NANDX1 G29684 (.A1(W292), .A2(I468), .ZN(W5948));
  NANDX1 G29685 (.A1(W7265), .A2(I1177), .ZN(W14247));
  NANDX1 G29686 (.A1(W8510), .A2(W1791), .ZN(W16631));
  NANDX1 G29687 (.A1(W11279), .A2(W6844), .ZN(W16628));
  NANDX1 G29688 (.A1(W14830), .A2(W5354), .ZN(W16627));
  NANDX1 G29689 (.A1(I1301), .A2(W359), .ZN(W14249));
  NANDX1 G29690 (.A1(W3900), .A2(W143), .ZN(W16570));
  NANDX1 G29691 (.A1(W7379), .A2(W3544), .ZN(O182));
  NANDX1 G29692 (.A1(W11725), .A2(I1922), .ZN(W14269));
  NANDX1 G29693 (.A1(W9520), .A2(W4557), .ZN(W14270));
  NANDX1 G29694 (.A1(W460), .A2(W553), .ZN(W5983));
  NANDX1 G29695 (.A1(W15546), .A2(W2304), .ZN(W16573));
  NANDX1 G29696 (.A1(W2427), .A2(W5593), .ZN(W5986));
  NANDX1 G29697 (.A1(W6645), .A2(I1640), .ZN(W16571));
  NANDX1 G29698 (.A1(W3193), .A2(I145), .ZN(W5987));
  NANDX1 G29699 (.A1(W530), .A2(W275), .ZN(W16579));
  NANDX1 G29700 (.A1(W7312), .A2(W10422), .ZN(W16568));
  NANDX1 G29701 (.A1(W5078), .A2(W4662), .ZN(W5994));
  NANDX1 G29702 (.A1(W185), .A2(W11274), .ZN(W14273));
  NANDX1 G29703 (.A1(I1339), .A2(W5150), .ZN(W7424));
  NANDX1 G29704 (.A1(W5598), .A2(W108), .ZN(W5996));
  NANDX1 G29705 (.A1(W7486), .A2(W9064), .ZN(W16565));
  NANDX1 G29706 (.A1(W1389), .A2(I346), .ZN(W5997));
  NANDX1 G29707 (.A1(W4469), .A2(W12852), .ZN(W14276));
  NANDX1 G29708 (.A1(W14666), .A2(W7931), .ZN(W16594));
  NANDX1 G29709 (.A1(W9286), .A2(W10892), .ZN(W16603));
  NANDX1 G29710 (.A1(I1299), .A2(W12442), .ZN(W14263));
  NANDX1 G29711 (.A1(W2304), .A2(W709), .ZN(W5963));
  NANDX1 G29712 (.A1(W5088), .A2(W1651), .ZN(O110));
  NANDX1 G29713 (.A1(W1556), .A2(W8473), .ZN(W14264));
  NANDX1 G29714 (.A1(W5058), .A2(W14475), .ZN(W16597));
  NANDX1 G29715 (.A1(W13808), .A2(W11491), .ZN(O1210));
  NANDX1 G29716 (.A1(W2626), .A2(W6747), .ZN(W14265));
  NANDX1 G29717 (.A1(W5762), .A2(W2232), .ZN(W7509));
  NANDX1 G29718 (.A1(W452), .A2(W6193), .ZN(W16592));
  NANDX1 G29719 (.A1(I957), .A2(W11708), .ZN(O1208));
  NANDX1 G29720 (.A1(W4278), .A2(W5018), .ZN(O112));
  NANDX1 G29721 (.A1(I1294), .A2(W6340), .ZN(W7428));
  NANDX1 G29722 (.A1(W2209), .A2(W15081), .ZN(W16587));
  NANDX1 G29723 (.A1(W15602), .A2(W14322), .ZN(W16586));
  NANDX1 G29724 (.A1(I1441), .A2(W9480), .ZN(W16584));
  NANDX1 G29725 (.A1(I1054), .A2(W2620), .ZN(W5973));
  NANDX1 G29726 (.A1(W657), .A2(W5562), .ZN(W14048));
  NANDX1 G29727 (.A1(W5508), .A2(W5096), .ZN(W17106));
  NANDX1 G29728 (.A1(W9784), .A2(W1981), .ZN(W14044));
  NANDX1 G29729 (.A1(W633), .A2(W4410), .ZN(W14045));
  NANDX1 G29730 (.A1(I54), .A2(W352), .ZN(W5630));
  NANDX1 G29731 (.A1(W11285), .A2(W13927), .ZN(W17101));
  NANDX1 G29732 (.A1(W4740), .A2(W5117), .ZN(W17100));
  NANDX1 G29733 (.A1(W11289), .A2(W7174), .ZN(W14046));
  NANDX1 G29734 (.A1(W2252), .A2(W899), .ZN(W17097));
  NANDX1 G29735 (.A1(W71), .A2(W4430), .ZN(W5632));
  NANDX1 G29736 (.A1(W12384), .A2(W10672), .ZN(W14040));
  NANDX1 G29737 (.A1(W601), .A2(W2749), .ZN(W7568));
  NANDX1 G29738 (.A1(W10445), .A2(W12839), .ZN(W17092));
  NANDX1 G29739 (.A1(I163), .A2(W2788), .ZN(W5635));
  NANDX1 G29740 (.A1(W4625), .A2(I1562), .ZN(W5638));
  NANDX1 G29741 (.A1(W157), .A2(W5275), .ZN(O821));
  NANDX1 G29742 (.A1(W1283), .A2(W5913), .ZN(W14056));
  NANDX1 G29743 (.A1(I1536), .A2(I344), .ZN(W17089));
  NANDX1 G29744 (.A1(W10901), .A2(W13943), .ZN(W17088));
  NANDX1 G29745 (.A1(W3212), .A2(W6253), .ZN(O1322));
  NANDX1 G29746 (.A1(W7103), .A2(W10287), .ZN(W14034));
  NANDX1 G29747 (.A1(W8816), .A2(W1121), .ZN(W17122));
  NANDX1 G29748 (.A1(W113), .A2(I681), .ZN(W17121));
  NANDX1 G29749 (.A1(W1292), .A2(W1842), .ZN(W5618));
  NANDX1 G29750 (.A1(W4760), .A2(W3125), .ZN(W14035));
  NANDX1 G29751 (.A1(W6183), .A2(W3809), .ZN(O1324));
  NANDX1 G29752 (.A1(W5191), .A2(W5675), .ZN(O1323));
  NANDX1 G29753 (.A1(W14986), .A2(W13811), .ZN(W17117));
  NANDX1 G29754 (.A1(W1362), .A2(I1381), .ZN(W5647));
  NANDX1 G29755 (.A1(W3678), .A2(W2939), .ZN(W5619));
  NANDX1 G29756 (.A1(W1722), .A2(W1112), .ZN(W5621));
  NANDX1 G29757 (.A1(W5834), .A2(W10755), .ZN(O818));
  NANDX1 G29758 (.A1(W1890), .A2(I1639), .ZN(W7577));
  NANDX1 G29759 (.A1(W15294), .A2(W17038), .ZN(W17112));
  NANDX1 G29760 (.A1(W8161), .A2(W15956), .ZN(O1321));
  NANDX1 G29761 (.A1(W4734), .A2(I1541), .ZN(W5623));
  NANDX1 G29762 (.A1(I1736), .A2(W6617), .ZN(W7573));
  NANDX1 G29763 (.A1(W4425), .A2(W3145), .ZN(W5674));
  NANDX1 G29764 (.A1(W2690), .A2(W4660), .ZN(W5668));
  NANDX1 G29765 (.A1(W12976), .A2(W14835), .ZN(W17059));
  NANDX1 G29766 (.A1(W1379), .A2(W2921), .ZN(W5670));
  NANDX1 G29767 (.A1(W10990), .A2(W11605), .ZN(W17056));
  NANDX1 G29768 (.A1(W14264), .A2(W7887), .ZN(W17055));
  NANDX1 G29769 (.A1(W8461), .A2(W818), .ZN(W17054));
  NANDX1 G29770 (.A1(W3781), .A2(I660), .ZN(W5671));
  NANDX1 G29771 (.A1(W1655), .A2(I514), .ZN(W5673));
  NANDX1 G29772 (.A1(W692), .A2(W2604), .ZN(W5663));
  NANDX1 G29773 (.A1(I636), .A2(W2043), .ZN(W5675));
  NANDX1 G29774 (.A1(W2700), .A2(W1952), .ZN(W5677));
  NANDX1 G29775 (.A1(W228), .A2(I223), .ZN(W5678));
  NANDX1 G29776 (.A1(W13949), .A2(W1128), .ZN(W17047));
  NANDX1 G29777 (.A1(W10793), .A2(W12137), .ZN(W17046));
  NANDX1 G29778 (.A1(W3167), .A2(W9237), .ZN(W14074));
  NANDX1 G29779 (.A1(W1887), .A2(W4640), .ZN(W5681));
  NANDX1 G29780 (.A1(W7052), .A2(W11645), .ZN(W17044));
  NANDX1 G29781 (.A1(W16690), .A2(W14973), .ZN(W17079));
  NANDX1 G29782 (.A1(W5081), .A2(I1293), .ZN(W7566));
  NANDX1 G29783 (.A1(I1045), .A2(W4033), .ZN(W14060));
  NANDX1 G29784 (.A1(I824), .A2(I198), .ZN(W5652));
  NANDX1 G29785 (.A1(I118), .A2(W2811), .ZN(W14061));
  NANDX1 G29786 (.A1(W2136), .A2(W1281), .ZN(W5653));
  NANDX1 G29787 (.A1(W1775), .A2(W8338), .ZN(O1314));
  NANDX1 G29788 (.A1(W1397), .A2(W342), .ZN(W17081));
  NANDX1 G29789 (.A1(W15299), .A2(W9631), .ZN(W17080));
  NANDX1 G29790 (.A1(W653), .A2(I530), .ZN(W5612));
  NANDX1 G29791 (.A1(I1306), .A2(I435), .ZN(W5655));
  NANDX1 G29792 (.A1(W16949), .A2(W8077), .ZN(W17077));
  NANDX1 G29793 (.A1(W2827), .A2(W606), .ZN(W5656));
  NANDX1 G29794 (.A1(W12099), .A2(W2264), .ZN(W14067));
  NANDX1 G29795 (.A1(I351), .A2(I752), .ZN(W5661));
  NANDX1 G29796 (.A1(I1792), .A2(W13706), .ZN(W14068));
  NANDX1 G29797 (.A1(W4475), .A2(W4525), .ZN(W14069));
  NANDX1 G29798 (.A1(W13312), .A2(W9848), .ZN(W17065));
  NANDX1 G29799 (.A1(I537), .A2(W8253), .ZN(O1340));
  NANDX1 G29800 (.A1(W689), .A2(W3644), .ZN(W17193));
  NANDX1 G29801 (.A1(W9832), .A2(W10380), .ZN(W17191));
  NANDX1 G29802 (.A1(W4076), .A2(W14904), .ZN(W17188));
  NANDX1 G29803 (.A1(W3812), .A2(I1911), .ZN(W7601));
  NANDX1 G29804 (.A1(I1925), .A2(W13245), .ZN(W14002));
  NANDX1 G29805 (.A1(W951), .A2(W7290), .ZN(O190));
  NANDX1 G29806 (.A1(I1582), .A2(W5261), .ZN(W7599));
  NANDX1 G29807 (.A1(W4297), .A2(W377), .ZN(W17179));
  NANDX1 G29808 (.A1(W1067), .A2(W1862), .ZN(W5568));
  NANDX1 G29809 (.A1(W5958), .A2(W4194), .ZN(W7602));
  NANDX1 G29810 (.A1(W1218), .A2(I792), .ZN(W5570));
  NANDX1 G29811 (.A1(W5726), .A2(W5344), .ZN(W7597));
  NANDX1 G29812 (.A1(W372), .A2(I521), .ZN(W5575));
  NANDX1 G29813 (.A1(W16342), .A2(W11077), .ZN(W17165));
  NANDX1 G29814 (.A1(W4812), .A2(W3663), .ZN(W17163));
  NANDX1 G29815 (.A1(W3877), .A2(W5182), .ZN(W7592));
  NANDX1 G29816 (.A1(W11699), .A2(W14999), .ZN(W17161));
  NANDX1 G29817 (.A1(W888), .A2(W3609), .ZN(W5578));
  NANDX1 G29818 (.A1(I1702), .A2(W14866), .ZN(O1346));
  NANDX1 G29819 (.A1(W2817), .A2(W7542), .ZN(W7610));
  NANDX1 G29820 (.A1(W10875), .A2(W632), .ZN(W17222));
  NANDX1 G29821 (.A1(W11021), .A2(W8516), .ZN(W17220));
  NANDX1 G29822 (.A1(W2120), .A2(W3707), .ZN(W7607));
  NANDX1 G29823 (.A1(W409), .A2(I169), .ZN(W5559));
  NANDX1 G29824 (.A1(I694), .A2(W538), .ZN(W5561));
  NANDX1 G29825 (.A1(W16345), .A2(W15368), .ZN(O1348));
  NANDX1 G29826 (.A1(W16066), .A2(W9942), .ZN(O1347));
  NANDX1 G29827 (.A1(W7298), .A2(I1439), .ZN(W14008));
  NANDX1 G29828 (.A1(I1533), .A2(I1054), .ZN(W5562));
  NANDX1 G29829 (.A1(W4268), .A2(W12669), .ZN(W13996));
  NANDX1 G29830 (.A1(W13498), .A2(W7246), .ZN(W17203));
  NANDX1 G29831 (.A1(I634), .A2(W15057), .ZN(W17202));
  NANDX1 G29832 (.A1(W16876), .A2(W14756), .ZN(O1344));
  NANDX1 G29833 (.A1(W14359), .A2(W10346), .ZN(O1342));
  NANDX1 G29834 (.A1(W1532), .A2(W976), .ZN(W7603));
  NANDX1 G29835 (.A1(W4858), .A2(W13324), .ZN(W17194));
  NANDX1 G29836 (.A1(W1980), .A2(W4295), .ZN(W5608));
  NANDX1 G29837 (.A1(W4115), .A2(I1029), .ZN(W5602));
  NANDX1 G29838 (.A1(W13539), .A2(W11264), .ZN(W14023));
  NANDX1 G29839 (.A1(W5567), .A2(W2725), .ZN(W7582));
  NANDX1 G29840 (.A1(W10941), .A2(W10410), .ZN(W17140));
  NANDX1 G29841 (.A1(W3750), .A2(W8529), .ZN(W17139));
  NANDX1 G29842 (.A1(W1880), .A2(W9076), .ZN(W17138));
  NANDX1 G29843 (.A1(W1079), .A2(W1276), .ZN(O95));
  NANDX1 G29844 (.A1(W3734), .A2(W612), .ZN(W5607));
  NANDX1 G29845 (.A1(I1204), .A2(W2895), .ZN(W5601));
  NANDX1 G29846 (.A1(W1200), .A2(W3435), .ZN(W17136));
  NANDX1 G29847 (.A1(W424), .A2(W13965), .ZN(W17135));
  NANDX1 G29848 (.A1(W9421), .A2(W8278), .ZN(W14025));
  NANDX1 G29849 (.A1(W17063), .A2(W5535), .ZN(O1329));
  NANDX1 G29850 (.A1(W15047), .A2(I234), .ZN(W17130));
  NANDX1 G29851 (.A1(W2280), .A2(W13432), .ZN(W17129));
  NANDX1 G29852 (.A1(W6259), .A2(W10855), .ZN(O1327));
  NANDX1 G29853 (.A1(W985), .A2(W4705), .ZN(W14033));
  NANDX1 G29854 (.A1(W16197), .A2(W5093), .ZN(W17151));
  NANDX1 G29855 (.A1(W12376), .A2(W12878), .ZN(W14010));
  NANDX1 G29856 (.A1(W1317), .A2(W8298), .ZN(O817));
  NANDX1 G29857 (.A1(W5351), .A2(W228), .ZN(W17158));
  NANDX1 G29858 (.A1(W5405), .A2(W3685), .ZN(W5587));
  NANDX1 G29859 (.A1(W8866), .A2(W9572), .ZN(O1336));
  NANDX1 G29860 (.A1(W1532), .A2(W1939), .ZN(W7590));
  NANDX1 G29861 (.A1(W12539), .A2(W12225), .ZN(W17152));
  NANDX1 G29862 (.A1(W8320), .A2(W8361), .ZN(W14017));
  NANDX1 G29863 (.A1(W3809), .A2(W5109), .ZN(W5682));
  NANDX1 G29864 (.A1(W4945), .A2(W5547), .ZN(W5589));
  NANDX1 G29865 (.A1(W1305), .A2(W4038), .ZN(W5591));
  NANDX1 G29866 (.A1(W13067), .A2(W6254), .ZN(W14018));
  NANDX1 G29867 (.A1(W5495), .A2(W2789), .ZN(W5595));
  NANDX1 G29868 (.A1(W3361), .A2(W1273), .ZN(W7585));
  NANDX1 G29869 (.A1(I184), .A2(W3475), .ZN(W5598));
  NANDX1 G29870 (.A1(W1990), .A2(W3480), .ZN(W5599));
  NANDX1 G29871 (.A1(W5024), .A2(W13819), .ZN(W14022));
  NANDX1 G29872 (.A1(W16250), .A2(I116), .ZN(W16901));
  NANDX1 G29873 (.A1(W5506), .A2(W3464), .ZN(W5758));
  NANDX1 G29874 (.A1(W1600), .A2(W2035), .ZN(W16911));
  NANDX1 G29875 (.A1(W4651), .A2(W1659), .ZN(W5761));
  NANDX1 G29876 (.A1(W1217), .A2(W457), .ZN(W5762));
  NANDX1 G29877 (.A1(W1162), .A2(W14340), .ZN(W16906));
  NANDX1 G29878 (.A1(I1054), .A2(W1092), .ZN(W7518));
  NANDX1 G29879 (.A1(W4938), .A2(W747), .ZN(W14137));
  NANDX1 G29880 (.A1(W3248), .A2(W3107), .ZN(W5769));
  NANDX1 G29881 (.A1(W7143), .A2(W4295), .ZN(W16902));
  NANDX1 G29882 (.A1(W3079), .A2(I1651), .ZN(W5757));
  NANDX1 G29883 (.A1(W4037), .A2(W3496), .ZN(W5773));
  NANDX1 G29884 (.A1(W11941), .A2(W1882), .ZN(O1276));
  NANDX1 G29885 (.A1(W14444), .A2(W7004), .ZN(W16894));
  NANDX1 G29886 (.A1(W5773), .A2(W322), .ZN(W16893));
  NANDX1 G29887 (.A1(W6329), .A2(W10988), .ZN(O829));
  NANDX1 G29888 (.A1(W14582), .A2(I1932), .ZN(W16889));
  NANDX1 G29889 (.A1(W8112), .A2(W9550), .ZN(W16887));
  NANDX1 G29890 (.A1(W59), .A2(W808), .ZN(W7513));
  NANDX1 G29891 (.A1(W1144), .A2(W7197), .ZN(W14125));
  NANDX1 G29892 (.A1(W3542), .A2(W276), .ZN(W5743));
  NANDX1 G29893 (.A1(W5441), .A2(I4), .ZN(W5745));
  NANDX1 G29894 (.A1(W8501), .A2(W12417), .ZN(W14123));
  NANDX1 G29895 (.A1(W11877), .A2(W6366), .ZN(W16932));
  NANDX1 G29896 (.A1(W16095), .A2(W8234), .ZN(W16930));
  NANDX1 G29897 (.A1(W15017), .A2(W3152), .ZN(W16929));
  NANDX1 G29898 (.A1(W2255), .A2(I70), .ZN(W5752));
  NANDX1 G29899 (.A1(W8662), .A2(W16527), .ZN(W16928));
  NANDX1 G29900 (.A1(W4496), .A2(W1801), .ZN(W5778));
  NANDX1 G29901 (.A1(W6340), .A2(I1167), .ZN(W16926));
  NANDX1 G29902 (.A1(W9463), .A2(I863), .ZN(W16925));
  NANDX1 G29903 (.A1(W3624), .A2(W6801), .ZN(W7523));
  NANDX1 G29904 (.A1(W856), .A2(W11264), .ZN(O1280));
  NANDX1 G29905 (.A1(W5090), .A2(W2504), .ZN(W16914));
  NANDX1 G29906 (.A1(W3780), .A2(W1032), .ZN(W14127));
  NANDX1 G29907 (.A1(W6607), .A2(W13344), .ZN(W14128));
  NANDX1 G29908 (.A1(W1354), .A2(W2029), .ZN(W7522));
  NANDX1 G29909 (.A1(W2542), .A2(W823), .ZN(W5806));
  NANDX1 G29910 (.A1(W16391), .A2(W4592), .ZN(W16867));
  NANDX1 G29911 (.A1(W3642), .A2(W11377), .ZN(O831));
  NANDX1 G29912 (.A1(W6288), .A2(W111), .ZN(W7511));
  NANDX1 G29913 (.A1(W12636), .A2(I1650), .ZN(W16865));
  NANDX1 G29914 (.A1(W4891), .A2(W2711), .ZN(W5800));
  NANDX1 G29915 (.A1(W3102), .A2(I191), .ZN(O102));
  NANDX1 G29916 (.A1(W12533), .A2(I356), .ZN(W16861));
  NANDX1 G29917 (.A1(W6757), .A2(W9427), .ZN(O1274));
  NANDX1 G29918 (.A1(W4579), .A2(W5457), .ZN(W5797));
  NANDX1 G29919 (.A1(W13122), .A2(W13956), .ZN(W16858));
  NANDX1 G29920 (.A1(W5417), .A2(I24), .ZN(W5807));
  NANDX1 G29921 (.A1(W13355), .A2(W9638), .ZN(W16856));
  NANDX1 G29922 (.A1(W16061), .A2(W12251), .ZN(W16855));
  NANDX1 G29923 (.A1(W2025), .A2(W2810), .ZN(W5808));
  NANDX1 G29924 (.A1(W6757), .A2(W10308), .ZN(W16851));
  NANDX1 G29925 (.A1(W5142), .A2(W208), .ZN(W16850));
  NANDX1 G29926 (.A1(W8736), .A2(W136), .ZN(W16849));
  NANDX1 G29927 (.A1(W5609), .A2(W9591), .ZN(W16876));
  NANDX1 G29928 (.A1(W10558), .A2(W5743), .ZN(W16883));
  NANDX1 G29929 (.A1(W4284), .A2(W2781), .ZN(W7512));
  NANDX1 G29930 (.A1(W445), .A2(W3917), .ZN(O830));
  NANDX1 G29931 (.A1(W2828), .A2(W987), .ZN(W5781));
  NANDX1 G29932 (.A1(W9384), .A2(W7228), .ZN(W14146));
  NANDX1 G29933 (.A1(W4058), .A2(W4198), .ZN(W5784));
  NANDX1 G29934 (.A1(W9122), .A2(I458), .ZN(W14147));
  NANDX1 G29935 (.A1(W2190), .A2(W2892), .ZN(W16880));
  NANDX1 G29936 (.A1(W4161), .A2(W3118), .ZN(O1285));
  NANDX1 G29937 (.A1(W7766), .A2(I49), .ZN(W16875));
  NANDX1 G29938 (.A1(W6873), .A2(W408), .ZN(W14148));
  NANDX1 G29939 (.A1(W13931), .A2(W7623), .ZN(W16874));
  NANDX1 G29940 (.A1(W6073), .A2(W10595), .ZN(W14149));
  NANDX1 G29941 (.A1(W3067), .A2(W4694), .ZN(W5792));
  NANDX1 G29942 (.A1(W2), .A2(W3985), .ZN(W5793));
  NANDX1 G29943 (.A1(W629), .A2(W5772), .ZN(W5794));
  NANDX1 G29944 (.A1(I20), .A2(W2600), .ZN(W14150));
  NANDX1 G29945 (.A1(W4892), .A2(W4712), .ZN(W5702));
  NANDX1 G29946 (.A1(W8433), .A2(W16273), .ZN(W17015));
  NANDX1 G29947 (.A1(I1212), .A2(W2437), .ZN(W5697));
  NANDX1 G29948 (.A1(W13633), .A2(W13568), .ZN(W14089));
  NANDX1 G29949 (.A1(W9383), .A2(W8133), .ZN(W14090));
  NANDX1 G29950 (.A1(W547), .A2(W15150), .ZN(W17012));
  NANDX1 G29951 (.A1(I206), .A2(W11864), .ZN(W14091));
  NANDX1 G29952 (.A1(W12762), .A2(W4806), .ZN(W17009));
  NANDX1 G29953 (.A1(W4288), .A2(W2835), .ZN(W17008));
  NANDX1 G29954 (.A1(W792), .A2(I1138), .ZN(W5701));
  NANDX1 G29955 (.A1(W13725), .A2(W7395), .ZN(O823));
  NANDX1 G29956 (.A1(I1094), .A2(W5022), .ZN(W5704));
  NANDX1 G29957 (.A1(I691), .A2(W5339), .ZN(W5708));
  NANDX1 G29958 (.A1(W7128), .A2(W2549), .ZN(O1298));
  NANDX1 G29959 (.A1(W549), .A2(W1438), .ZN(W5709));
  NANDX1 G29960 (.A1(W5912), .A2(W6011), .ZN(W7541));
  NANDX1 G29961 (.A1(I1497), .A2(I1301), .ZN(W5711));
  NANDX1 G29962 (.A1(W957), .A2(W7197), .ZN(W17000));
  NANDX1 G29963 (.A1(W5263), .A2(W4199), .ZN(W7540));
  NANDX1 G29964 (.A1(W5624), .A2(W11132), .ZN(W17031));
  NANDX1 G29965 (.A1(W13059), .A2(W1521), .ZN(W14075));
  NANDX1 G29966 (.A1(I672), .A2(W5920), .ZN(W7551));
  NANDX1 G29967 (.A1(I1290), .A2(I542), .ZN(W5684));
  NANDX1 G29968 (.A1(W9995), .A2(W5711), .ZN(W17037));
  NANDX1 G29969 (.A1(W4722), .A2(W3302), .ZN(W7549));
  NANDX1 G29970 (.A1(W4002), .A2(W809), .ZN(W14081));
  NANDX1 G29971 (.A1(W5702), .A2(W8458), .ZN(W17034));
  NANDX1 G29972 (.A1(W16947), .A2(W11553), .ZN(O1304));
  NANDX1 G29973 (.A1(I1578), .A2(W292), .ZN(W16995));
  NANDX1 G29974 (.A1(W16277), .A2(W7417), .ZN(W17030));
  NANDX1 G29975 (.A1(W5535), .A2(W4189), .ZN(W5691));
  NANDX1 G29976 (.A1(I1480), .A2(W269), .ZN(W5693));
  NANDX1 G29977 (.A1(W2351), .A2(W6927), .ZN(W17026));
  NANDX1 G29978 (.A1(W7512), .A2(W14449), .ZN(W17022));
  NANDX1 G29979 (.A1(I1596), .A2(W7500), .ZN(W17020));
  NANDX1 G29980 (.A1(W1663), .A2(W6228), .ZN(W7545));
  NANDX1 G29981 (.A1(W9210), .A2(W5256), .ZN(O1300));
  NANDX1 G29982 (.A1(W9304), .A2(W13547), .ZN(W16949));
  NANDX1 G29983 (.A1(W1205), .A2(W11276), .ZN(W14108));
  NANDX1 G29984 (.A1(W7645), .A2(W11055), .ZN(W14110));
  NANDX1 G29985 (.A1(W2024), .A2(W10869), .ZN(W14114));
  NANDX1 G29986 (.A1(W11851), .A2(W3266), .ZN(W16956));
  NANDX1 G29987 (.A1(I1201), .A2(W1326), .ZN(W5730));
  NANDX1 G29988 (.A1(I1058), .A2(W16946), .ZN(W16953));
  NANDX1 G29989 (.A1(W4336), .A2(W623), .ZN(W5731));
  NANDX1 G29990 (.A1(W10978), .A2(W8625), .ZN(W16951));
  NANDX1 G29991 (.A1(W15936), .A2(W14427), .ZN(O1288));
  NANDX1 G29992 (.A1(I1189), .A2(W10333), .ZN(W14117));
  NANDX1 G29993 (.A1(W641), .A2(W5422), .ZN(W16945));
  NANDX1 G29994 (.A1(W2131), .A2(W1474), .ZN(O188));
  NANDX1 G29995 (.A1(W15011), .A2(I1409), .ZN(W16940));
  NANDX1 G29996 (.A1(W2702), .A2(W5406), .ZN(W5735));
  NANDX1 G29997 (.A1(W7912), .A2(W4661), .ZN(W16936));
  NANDX1 G29998 (.A1(I1824), .A2(W4348), .ZN(W5740));
  NANDX1 G29999 (.A1(W537), .A2(W5314), .ZN(W5742));
  NANDX1 G30000 (.A1(W14529), .A2(W15582), .ZN(W16981));
  NANDX1 G30001 (.A1(W1438), .A2(W1087), .ZN(W16994));
  NANDX1 G30002 (.A1(W11693), .A2(W15352), .ZN(W16993));
  NANDX1 G30003 (.A1(W16696), .A2(W11180), .ZN(W16991));
  NANDX1 G30004 (.A1(W9451), .A2(W14057), .ZN(O824));
  NANDX1 G30005 (.A1(W9694), .A2(W448), .ZN(W16988));
  NANDX1 G30006 (.A1(W6190), .A2(W5213), .ZN(W7538));
  NANDX1 G30007 (.A1(I206), .A2(W2652), .ZN(W5716));
  NANDX1 G30008 (.A1(W1473), .A2(W2220), .ZN(W5717));
  NANDX1 G30009 (.A1(W484), .A2(W16188), .ZN(W20185));
  NANDX1 G30010 (.A1(W1444), .A2(W8653), .ZN(W14102));
  NANDX1 G30011 (.A1(W11287), .A2(W16068), .ZN(W16979));
  NANDX1 G30012 (.A1(W7998), .A2(W12419), .ZN(W16971));
  NANDX1 G30013 (.A1(I686), .A2(W4707), .ZN(W7534));
  NANDX1 G30014 (.A1(W11266), .A2(W3546), .ZN(W16967));
  NANDX1 G30015 (.A1(W573), .A2(W4471), .ZN(W5720));
  NANDX1 G30016 (.A1(W1632), .A2(W10241), .ZN(W16966));
  NANDX1 G30017 (.A1(W3111), .A2(W8862), .ZN(W14105));
  NANDX1 G30018 (.A1(W4857), .A2(W17183), .ZN(W22911));
  NANDX1 G30019 (.A1(W10118), .A2(W21905), .ZN(W22902));
  NANDX1 G30020 (.A1(W814), .A2(I1593), .ZN(W9466));
  NANDX1 G30021 (.A1(I360), .A2(W367), .ZN(W1669));
  NANDX1 G30022 (.A1(W1373), .A2(W970), .ZN(W1668));
  NANDX1 G30023 (.A1(I1398), .A2(W1478), .ZN(W1666));
  NANDX1 G30024 (.A1(W5632), .A2(W10705), .ZN(W22904));
  NANDX1 G30025 (.A1(I1688), .A2(I71), .ZN(W1665));
  NANDX1 G30026 (.A1(W420), .A2(W3650), .ZN(W10552));
  NANDX1 G30027 (.A1(W18504), .A2(W6043), .ZN(O2634));
  NANDX1 G30028 (.A1(W13514), .A2(W12904), .ZN(W24576));
  NANDX1 G30029 (.A1(W1548), .A2(W1290), .ZN(W1663));
  NANDX1 G30030 (.A1(W9455), .A2(I1809), .ZN(O498));
  NANDX1 G30031 (.A1(W4847), .A2(W4734), .ZN(O2635));
  NANDX1 G30032 (.A1(W1412), .A2(W8416), .ZN(W9963));
  NANDX1 G30033 (.A1(W1334), .A2(W3247), .ZN(W11306));
  NANDX1 G30034 (.A1(I1088), .A2(I1089), .ZN(W544));
  NANDX1 G30035 (.A1(W22589), .A2(W17359), .ZN(O3123));
  NANDX1 G30036 (.A1(I968), .A2(W787), .ZN(W1658));
  NANDX1 G30037 (.A1(W15399), .A2(W22035), .ZN(W24572));
  NANDX1 G30038 (.A1(W16313), .A2(W4421), .ZN(W22918));
  NANDX1 G30039 (.A1(W8027), .A2(W4525), .ZN(W10553));
  NANDX1 G30040 (.A1(W5905), .A2(W6125), .ZN(W10554));
  NANDX1 G30041 (.A1(W6114), .A2(I1447), .ZN(W9471));
  NANDX1 G30042 (.A1(W8430), .A2(W171), .ZN(O404));
  NANDX1 G30043 (.A1(W7272), .A2(W7817), .ZN(W9473));
  NANDX1 G30044 (.A1(W896), .A2(W8276), .ZN(W22921));
  NANDX1 G30045 (.A1(W7692), .A2(W20724), .ZN(W22922));
  NANDX1 G30046 (.A1(I1102), .A2(I1103), .ZN(W551));
  NANDX1 G30047 (.A1(I498), .A2(I1119), .ZN(W1651));
  NANDX1 G30048 (.A1(W300), .A2(I158), .ZN(W1650));
  NANDX1 G30049 (.A1(W3101), .A2(I1864), .ZN(W22890));
  NANDX1 G30050 (.A1(W121), .A2(W2868), .ZN(W9451));
  NANDX1 G30051 (.A1(W4032), .A2(W6700), .ZN(W9454));
  NANDX1 G30052 (.A1(W14086), .A2(W16394), .ZN(W24590));
  NANDX1 G30053 (.A1(W3834), .A2(W8070), .ZN(W9455));
  NANDX1 G30054 (.A1(W893), .A2(W718), .ZN(W11322));
  NANDX1 G30055 (.A1(I1074), .A2(I1075), .ZN(W537));
  NANDX1 G30056 (.A1(W19195), .A2(W5199), .ZN(W24585));
  NANDX1 G30057 (.A1(W643), .A2(W762), .ZN(W1692));
  NANDX1 G30058 (.A1(W947), .A2(W1543), .ZN(W10547));
  NANDX1 G30059 (.A1(W290), .A2(W7233), .ZN(W9460));
  NANDX1 G30060 (.A1(W5), .A2(W1025), .ZN(O346));
  NANDX1 G30061 (.A1(W5026), .A2(W3817), .ZN(W22884));
  NANDX1 G30062 (.A1(I989), .A2(I1123), .ZN(W1685));
  NANDX1 G30063 (.A1(W5245), .A2(W7708), .ZN(W22888));
  NANDX1 G30064 (.A1(W91), .A2(W408), .ZN(W1684));
  NANDX1 G30065 (.A1(W13629), .A2(W16302), .ZN(O2638));
  NANDX1 G30066 (.A1(W1356), .A2(W20690), .ZN(O2628));
  NANDX1 G30067 (.A1(W584), .A2(I1908), .ZN(W1679));
  NANDX1 G30068 (.A1(I496), .A2(W1265), .ZN(W1678));
  NANDX1 G30069 (.A1(W6921), .A2(I272), .ZN(W11317));
  NANDX1 G30070 (.A1(W6110), .A2(W3079), .ZN(W10549));
  NANDX1 G30071 (.A1(W8796), .A2(W1194), .ZN(O2631));
  NANDX1 G30072 (.A1(W17437), .A2(W4582), .ZN(W22897));
  NANDX1 G30073 (.A1(W3397), .A2(W5812), .ZN(W9463));
  NANDX1 G30074 (.A1(W5519), .A2(W8828), .ZN(W11313));
  NANDX1 G30075 (.A1(I1086), .A2(I1087), .ZN(W543));
  NANDX1 G30076 (.A1(W8744), .A2(I1686), .ZN(W10551));
  NANDX1 G30077 (.A1(W20319), .A2(W6972), .ZN(W22900));
  NANDX1 G30078 (.A1(W10621), .A2(W1331), .ZN(O2632));
  NANDX1 G30079 (.A1(I1254), .A2(W8321), .ZN(W9465));
  NANDX1 G30080 (.A1(W19496), .A2(W3778), .ZN(O2647));
  NANDX1 G30081 (.A1(W1740), .A2(W19262), .ZN(O2645));
  NANDX1 G30082 (.A1(I1730), .A2(W1350), .ZN(W1634));
  NANDX1 G30083 (.A1(W458), .A2(I1846), .ZN(W1633));
  NANDX1 G30084 (.A1(I1132), .A2(I1133), .ZN(W566));
  NANDX1 G30085 (.A1(W2996), .A2(W5221), .ZN(W9480));
  NANDX1 G30086 (.A1(I1134), .A2(I1135), .ZN(W567));
  NANDX1 G30087 (.A1(I50), .A2(W1613), .ZN(W1630));
  NANDX1 G30088 (.A1(W22915), .A2(W15556), .ZN(W24554));
  NANDX1 G30089 (.A1(W817), .A2(W6859), .ZN(W10561));
  NANDX1 G30090 (.A1(W8053), .A2(W8944), .ZN(O496));
  NANDX1 G30091 (.A1(I600), .A2(W10368), .ZN(W11281));
  NANDX1 G30092 (.A1(W18712), .A2(W13496), .ZN(W24552));
  NANDX1 G30093 (.A1(W8169), .A2(I1934), .ZN(W11280));
  NANDX1 G30094 (.A1(W2562), .A2(W5988), .ZN(W9481));
  NANDX1 G30095 (.A1(I1051), .A2(I75), .ZN(W1615));
  NANDX1 G30096 (.A1(I1130), .A2(I1131), .ZN(W565));
  NANDX1 G30097 (.A1(W13429), .A2(W8206), .ZN(W22972));
  NANDX1 G30098 (.A1(I1865), .A2(I1798), .ZN(W1614));
  NANDX1 G30099 (.A1(W10259), .A2(W5622), .ZN(W11275));
  NANDX1 G30100 (.A1(W4808), .A2(W8312), .ZN(W11274));
  NANDX1 G30101 (.A1(I713), .A2(I154), .ZN(W1610));
  NANDX1 G30102 (.A1(W1338), .A2(W38), .ZN(W1607));
  NANDX1 G30103 (.A1(W826), .A2(W16403), .ZN(O2649));
  NANDX1 G30104 (.A1(W2285), .A2(W5837), .ZN(W9482));
  NANDX1 G30105 (.A1(W19503), .A2(W5392), .ZN(W22983));
  NANDX1 G30106 (.A1(W501), .A2(W1668), .ZN(O294));
  NANDX1 G30107 (.A1(W131), .A2(W4850), .ZN(W9484));
  NANDX1 G30108 (.A1(W1571), .A2(I1939), .ZN(W1603));
  NANDX1 G30109 (.A1(W21618), .A2(W799), .ZN(W24550));
  NANDX1 G30110 (.A1(I1614), .A2(W8105), .ZN(W11266));
  NANDX1 G30111 (.A1(W17490), .A2(W10530), .ZN(W22943));
  NANDX1 G30112 (.A1(I1112), .A2(I1113), .ZN(W556));
  NANDX1 G30113 (.A1(I1382), .A2(I10), .ZN(W1649));
  NANDX1 G30114 (.A1(W6710), .A2(W7547), .ZN(W11299));
  NANDX1 G30115 (.A1(I162), .A2(I535), .ZN(W1648));
  NANDX1 G30116 (.A1(W11008), .A2(W8768), .ZN(W22931));
  NANDX1 G30117 (.A1(I1372), .A2(W2913), .ZN(W22932));
  NANDX1 G30118 (.A1(W9649), .A2(W9822), .ZN(W11297));
  NANDX1 G30119 (.A1(W8552), .A2(W13564), .ZN(W24566));
  NANDX1 G30120 (.A1(W7815), .A2(W17770), .ZN(O3119));
  NANDX1 G30121 (.A1(I1114), .A2(I1115), .ZN(W557));
  NANDX1 G30122 (.A1(W14071), .A2(W4483), .ZN(O2641));
  NANDX1 G30123 (.A1(W20923), .A2(W17592), .ZN(W22936));
  NANDX1 G30124 (.A1(I1116), .A2(I1117), .ZN(W558));
  NANDX1 G30125 (.A1(I1166), .A2(W11034), .ZN(O3118));
  NANDX1 G30126 (.A1(W7209), .A2(W245), .ZN(W9478));
  NANDX1 G30127 (.A1(W13276), .A2(W9696), .ZN(W22865));
  NANDX1 G30128 (.A1(W7523), .A2(I597), .ZN(W22944));
  NANDX1 G30129 (.A1(W9270), .A2(W8461), .ZN(W9479));
  NANDX1 G30130 (.A1(W12615), .A2(W12498), .ZN(W22946));
  NANDX1 G30131 (.A1(W1575), .A2(I468), .ZN(W1643));
  NANDX1 G30132 (.A1(W287), .A2(I1080), .ZN(W1641));
  NANDX1 G30133 (.A1(W11016), .A2(W1056), .ZN(W11293));
  NANDX1 G30134 (.A1(W11539), .A2(W9943), .ZN(W22950));
  NANDX1 G30135 (.A1(W19922), .A2(W17750), .ZN(O2643));
  NANDX1 G30136 (.A1(W15313), .A2(W18188), .ZN(O3117));
  NANDX1 G30137 (.A1(I1128), .A2(I1129), .ZN(W564));
  NANDX1 G30138 (.A1(W19213), .A2(W2659), .ZN(W22954));
  NANDX1 G30139 (.A1(I1171), .A2(I501), .ZN(W1635));
  NANDX1 G30140 (.A1(W3206), .A2(W16477), .ZN(W22956));
  NANDX1 G30141 (.A1(W10101), .A2(W4140), .ZN(W11292));
  NANDX1 G30142 (.A1(W21863), .A2(W4978), .ZN(W24620));
  NANDX1 G30143 (.A1(W983), .A2(W4876), .ZN(W22792));
  NANDX1 G30144 (.A1(W11894), .A2(W4718), .ZN(O3149));
  NANDX1 G30145 (.A1(W1466), .A2(I629), .ZN(W1749));
  NANDX1 G30146 (.A1(W10442), .A2(W2623), .ZN(W22793));
  NANDX1 G30147 (.A1(I683), .A2(W8506), .ZN(W10533));
  NANDX1 G30148 (.A1(W15371), .A2(I496), .ZN(W22794));
  NANDX1 G30149 (.A1(W824), .A2(W768), .ZN(W10535));
  NANDX1 G30150 (.A1(W1122), .A2(I1684), .ZN(W1748));
  NANDX1 G30151 (.A1(W2587), .A2(W3125), .ZN(W11363));
  NANDX1 G30152 (.A1(I1040), .A2(I1041), .ZN(W520));
  NANDX1 G30153 (.A1(I854), .A2(W5642), .ZN(W22796));
  NANDX1 G30154 (.A1(W12157), .A2(I705), .ZN(W22797));
  NANDX1 G30155 (.A1(W4487), .A2(W11096), .ZN(W24622));
  NANDX1 G30156 (.A1(W20092), .A2(W10977), .ZN(W24621));
  NANDX1 G30157 (.A1(W515), .A2(I1449), .ZN(W11362));
  NANDX1 G30158 (.A1(I223), .A2(W3725), .ZN(W9419));
  NANDX1 G30159 (.A1(W8371), .A2(W84), .ZN(W9426));
  NANDX1 G30160 (.A1(W6728), .A2(W12438), .ZN(W22801));
  NANDX1 G30161 (.A1(W17464), .A2(W14653), .ZN(W22803));
  NANDX1 G30162 (.A1(W4314), .A2(W21003), .ZN(W22808));
  NANDX1 G30163 (.A1(I415), .A2(I78), .ZN(W1746));
  NANDX1 G30164 (.A1(W17592), .A2(W3201), .ZN(W22811));
  NANDX1 G30165 (.A1(W1541), .A2(I1350), .ZN(W1744));
  NANDX1 G30166 (.A1(W1019), .A2(W588), .ZN(W1743));
  NANDX1 G30167 (.A1(W17354), .A2(W12047), .ZN(O3144));
  NANDX1 G30168 (.A1(W1574), .A2(W1481), .ZN(W1742));
  NANDX1 G30169 (.A1(W7281), .A2(I685), .ZN(W11360));
  NANDX1 G30170 (.A1(W5680), .A2(W1312), .ZN(W9429));
  NANDX1 G30171 (.A1(W11206), .A2(W1690), .ZN(W22814));
  NANDX1 G30172 (.A1(W7259), .A2(W9250), .ZN(W22815));
  NANDX1 G30173 (.A1(I454), .A2(I289), .ZN(W1763));
  NANDX1 G30174 (.A1(I1018), .A2(I1019), .ZN(W509));
  NANDX1 G30175 (.A1(W10412), .A2(W17596), .ZN(O2604));
  NANDX1 G30176 (.A1(W4520), .A2(I1562), .ZN(W11377));
  NANDX1 G30177 (.A1(W8718), .A2(W1658), .ZN(W11375));
  NANDX1 G30178 (.A1(I781), .A2(I1480), .ZN(W1774));
  NANDX1 G30179 (.A1(W5979), .A2(W7493), .ZN(W9410));
  NANDX1 G30180 (.A1(W21391), .A2(W8884), .ZN(O2607));
  NANDX1 G30181 (.A1(W4612), .A2(W123), .ZN(W9412));
  NANDX1 G30182 (.A1(W19413), .A2(W6346), .ZN(W22769));
  NANDX1 G30183 (.A1(I1308), .A2(W1752), .ZN(W9414));
  NANDX1 G30184 (.A1(W3993), .A2(W2471), .ZN(O288));
  NANDX1 G30185 (.A1(I1563), .A2(W126), .ZN(W1768));
  NANDX1 G30186 (.A1(W3306), .A2(W2969), .ZN(W9973));
  NANDX1 G30187 (.A1(W7862), .A2(W6411), .ZN(O289));
  NANDX1 G30188 (.A1(I1026), .A2(I1027), .ZN(W513));
  NANDX1 G30189 (.A1(I1042), .A2(I1043), .ZN(W521));
  NANDX1 G30190 (.A1(I1802), .A2(W564), .ZN(W1762));
  NANDX1 G30191 (.A1(W1524), .A2(I1813), .ZN(W1761));
  NANDX1 G30192 (.A1(W19195), .A2(W4592), .ZN(W22776));
  NANDX1 G30193 (.A1(W1045), .A2(W1652), .ZN(W1760));
  NANDX1 G30194 (.A1(W512), .A2(I833), .ZN(W1758));
  NANDX1 G30195 (.A1(W4979), .A2(W3730), .ZN(W22778));
  NANDX1 G30196 (.A1(I1668), .A2(W5143), .ZN(W9417));
  NANDX1 G30197 (.A1(W4590), .A2(W8592), .ZN(W11367));
  NANDX1 G30198 (.A1(W5245), .A2(W7342), .ZN(W22781));
  NANDX1 G30199 (.A1(W11254), .A2(W15039), .ZN(W22783));
  NANDX1 G30200 (.A1(W7541), .A2(W8160), .ZN(W22786));
  NANDX1 G30201 (.A1(I1115), .A2(W1640), .ZN(W1754));
  NANDX1 G30202 (.A1(W9096), .A2(W9178), .ZN(W9418));
  NANDX1 G30203 (.A1(W10685), .A2(W21617), .ZN(W24633));
  NANDX1 G30204 (.A1(W1204), .A2(W8597), .ZN(W9447));
  NANDX1 G30205 (.A1(I1058), .A2(I1059), .ZN(W529));
  NANDX1 G30206 (.A1(W10319), .A2(W2917), .ZN(W22840));
  NANDX1 G30207 (.A1(W7935), .A2(W5776), .ZN(W22841));
  NANDX1 G30208 (.A1(W2263), .A2(I1156), .ZN(W11340));
  NANDX1 G30209 (.A1(I1680), .A2(I787), .ZN(W1718));
  NANDX1 G30210 (.A1(W2374), .A2(W775), .ZN(W10545));
  NANDX1 G30211 (.A1(W6311), .A2(W8650), .ZN(W9441));
  NANDX1 G30212 (.A1(W6837), .A2(W1039), .ZN(W9445));
  NANDX1 G30213 (.A1(I1518), .A2(I1556), .ZN(W1714));
  NANDX1 G30214 (.A1(W1510), .A2(W582), .ZN(W1712));
  NANDX1 G30215 (.A1(W9306), .A2(W8622), .ZN(W11337));
  NANDX1 G30216 (.A1(W8753), .A2(W4620), .ZN(O500));
  NANDX1 G30217 (.A1(W5858), .A2(W9271), .ZN(W9446));
  NANDX1 G30218 (.A1(W2439), .A2(W5954), .ZN(W11334));
  NANDX1 G30219 (.A1(W10789), .A2(W18008), .ZN(W24596));
  NANDX1 G30220 (.A1(I793), .A2(I1139), .ZN(W22838));
  NANDX1 G30221 (.A1(I1068), .A2(I1069), .ZN(W534));
  NANDX1 G30222 (.A1(W7347), .A2(W7431), .ZN(W24593));
  NANDX1 G30223 (.A1(W2695), .A2(I433), .ZN(W11329));
  NANDX1 G30224 (.A1(W2674), .A2(W5774), .ZN(W11328));
  NANDX1 G30225 (.A1(I360), .A2(W408), .ZN(W1702));
  NANDX1 G30226 (.A1(W19216), .A2(W8742), .ZN(O3131));
  NANDX1 G30227 (.A1(W4098), .A2(W1388), .ZN(W9449));
  NANDX1 G30228 (.A1(W7548), .A2(W9198), .ZN(W11327));
  NANDX1 G30229 (.A1(W1257), .A2(W1025), .ZN(W1699));
  NANDX1 G30230 (.A1(W5576), .A2(W10944), .ZN(W22856));
  NANDX1 G30231 (.A1(W9639), .A2(W22645), .ZN(W22858));
  NANDX1 G30232 (.A1(W5027), .A2(W8759), .ZN(W11326));
  NANDX1 G30233 (.A1(W815), .A2(I637), .ZN(W11324));
  NANDX1 G30234 (.A1(W11476), .A2(I999), .ZN(O2622));
  NANDX1 G30235 (.A1(W9023), .A2(W2190), .ZN(W9435));
  NANDX1 G30236 (.A1(W2013), .A2(W8925), .ZN(O2618));
  NANDX1 G30237 (.A1(W17181), .A2(W11372), .ZN(W24616));
  NANDX1 G30238 (.A1(I1884), .A2(W53), .ZN(W1735));
  NANDX1 G30239 (.A1(W8169), .A2(W13536), .ZN(O3141));
  NANDX1 G30240 (.A1(W19789), .A2(I1980), .ZN(W22822));
  NANDX1 G30241 (.A1(W296), .A2(W1947), .ZN(W9430));
  NANDX1 G30242 (.A1(W8426), .A2(W9312), .ZN(W22826));
  NANDX1 G30243 (.A1(W550), .A2(W1032), .ZN(W1734));
  NANDX1 G30244 (.A1(W2481), .A2(W11044), .ZN(W22827));
  NANDX1 G30245 (.A1(W8337), .A2(W4597), .ZN(W10536));
  NANDX1 G30246 (.A1(W15797), .A2(W20146), .ZN(W22828));
  NANDX1 G30247 (.A1(W58), .A2(I1960), .ZN(O15));
  NANDX1 G30248 (.A1(W6702), .A2(I1453), .ZN(W11351));
  NANDX1 G30249 (.A1(W1265), .A2(W6792), .ZN(W10537));
  NANDX1 G30250 (.A1(I1044), .A2(I1045), .ZN(W522));
  NANDX1 G30251 (.A1(I1853), .A2(I1863), .ZN(W1599));
  NANDX1 G30252 (.A1(W809), .A2(I488), .ZN(W10538));
  NANDX1 G30253 (.A1(W6620), .A2(W7667), .ZN(W11346));
  NANDX1 G30254 (.A1(I1046), .A2(I1047), .ZN(W523));
  NANDX1 G30255 (.A1(W14574), .A2(W18216), .ZN(W22833));
  NANDX1 G30256 (.A1(W17608), .A2(W17789), .ZN(W24606));
  NANDX1 G30257 (.A1(W6799), .A2(W166), .ZN(W11345));
  NANDX1 G30258 (.A1(I1107), .A2(I1339), .ZN(W22834));
  NANDX1 G30259 (.A1(I1050), .A2(I1051), .ZN(W525));
  NANDX1 G30260 (.A1(I1052), .A2(I1053), .ZN(W526));
  NANDX1 G30261 (.A1(W1694), .A2(W1199), .ZN(W1725));
  NANDX1 G30262 (.A1(W14358), .A2(W22326), .ZN(W22837));
  NANDX1 G30263 (.A1(I1054), .A2(I1055), .ZN(W527));
  NANDX1 G30264 (.A1(W3817), .A2(W8981), .ZN(W11341));
  NANDX1 G30265 (.A1(W6516), .A2(W1671), .ZN(W9970));
  NANDX1 G30266 (.A1(W9069), .A2(W2525), .ZN(W9553));
  NANDX1 G30267 (.A1(W2731), .A2(W5425), .ZN(W9550));
  NANDX1 G30268 (.A1(W12543), .A2(W23127), .ZN(W23130));
  NANDX1 G30269 (.A1(W15928), .A2(W9456), .ZN(W23132));
  NANDX1 G30270 (.A1(W15450), .A2(I1044), .ZN(W23134));
  NANDX1 G30271 (.A1(I1216), .A2(I1217), .ZN(W608));
  NANDX1 G30272 (.A1(W14430), .A2(W20716), .ZN(O2684));
  NANDX1 G30273 (.A1(W3566), .A2(W5938), .ZN(W10580));
  NANDX1 G30274 (.A1(W20203), .A2(W18004), .ZN(W23136));
  NANDX1 G30275 (.A1(W750), .A2(W22871), .ZN(O2687));
  NANDX1 G30276 (.A1(W226), .A2(W8687), .ZN(W11202));
  NANDX1 G30277 (.A1(W3519), .A2(W832), .ZN(W9552));
  NANDX1 G30278 (.A1(W90), .A2(W6882), .ZN(W11200));
  NANDX1 G30279 (.A1(I1218), .A2(I1219), .ZN(W609));
  NANDX1 G30280 (.A1(W13092), .A2(W22257), .ZN(O2689));
  NANDX1 G30281 (.A1(W10018), .A2(W8590), .ZN(W24494));
  NANDX1 G30282 (.A1(W12749), .A2(W12254), .ZN(O3100));
  NANDX1 G30283 (.A1(W5785), .A2(W3941), .ZN(O2692));
  NANDX1 G30284 (.A1(W1494), .A2(W14834), .ZN(W23149));
  NANDX1 G30285 (.A1(I164), .A2(I400), .ZN(W11196));
  NANDX1 G30286 (.A1(W16806), .A2(W18502), .ZN(W23151));
  NANDX1 G30287 (.A1(W8955), .A2(W20513), .ZN(W23155));
  NANDX1 G30288 (.A1(W803), .A2(I832), .ZN(W1508));
  NANDX1 G30289 (.A1(W5392), .A2(W17775), .ZN(W23156));
  NANDX1 G30290 (.A1(W1105), .A2(I1965), .ZN(W1507));
  NANDX1 G30291 (.A1(W5716), .A2(W3859), .ZN(W9557));
  NANDX1 G30292 (.A1(I469), .A2(W10145), .ZN(W11189));
  NANDX1 G30293 (.A1(I1231), .A2(I681), .ZN(W1504));
  NANDX1 G30294 (.A1(W3701), .A2(W1388), .ZN(W9558));
  NANDX1 G30295 (.A1(W8900), .A2(W6336), .ZN(O3099));
  NANDX1 G30296 (.A1(W7747), .A2(W19110), .ZN(W23164));
  NANDX1 G30297 (.A1(I1208), .A2(I1209), .ZN(W604));
  NANDX1 G30298 (.A1(W5150), .A2(W14564), .ZN(W23098));
  NANDX1 G30299 (.A1(W325), .A2(I1442), .ZN(W1531));
  NANDX1 G30300 (.A1(I1272), .A2(W7335), .ZN(W9532));
  NANDX1 G30301 (.A1(W14210), .A2(W2013), .ZN(O3105));
  NANDX1 G30302 (.A1(W47), .A2(W697), .ZN(W1525));
  NANDX1 G30303 (.A1(W2140), .A2(W4858), .ZN(W9534));
  NANDX1 G30304 (.A1(I1476), .A2(I1414), .ZN(W9537));
  NANDX1 G30305 (.A1(I376), .A2(W4212), .ZN(W9539));
  NANDX1 G30306 (.A1(W12212), .A2(W15408), .ZN(O2678));
  NANDX1 G30307 (.A1(W275), .A2(W932), .ZN(W1520));
  NANDX1 G30308 (.A1(I506), .A2(I31), .ZN(W1519));
  NANDX1 G30309 (.A1(I409), .A2(W1411), .ZN(W23110));
  NANDX1 G30310 (.A1(W14241), .A2(W2179), .ZN(W23111));
  NANDX1 G30311 (.A1(W1416), .A2(I680), .ZN(W1518));
  NANDX1 G30312 (.A1(W15590), .A2(W5306), .ZN(O3104));
  NANDX1 G30313 (.A1(I1928), .A2(W622), .ZN(W1503));
  NANDX1 G30314 (.A1(W586), .A2(W19358), .ZN(O2679));
  NANDX1 G30315 (.A1(W1300), .A2(W21281), .ZN(W24502));
  NANDX1 G30316 (.A1(W14291), .A2(W10552), .ZN(W23114));
  NANDX1 G30317 (.A1(W1729), .A2(W19814), .ZN(W23117));
  NANDX1 G30318 (.A1(I1214), .A2(I1215), .ZN(W607));
  NANDX1 G30319 (.A1(W4295), .A2(W7612), .ZN(W9548));
  NANDX1 G30320 (.A1(W22522), .A2(W21990), .ZN(O2681));
  NANDX1 G30321 (.A1(I915), .A2(I1865), .ZN(W1515));
  NANDX1 G30322 (.A1(W14850), .A2(W6235), .ZN(W24500));
  NANDX1 G30323 (.A1(W15228), .A2(W5489), .ZN(O3101));
  NANDX1 G30324 (.A1(W22922), .A2(W21763), .ZN(W23119));
  NANDX1 G30325 (.A1(W10014), .A2(I945), .ZN(W23121));
  NANDX1 G30326 (.A1(W9569), .A2(W86), .ZN(W23122));
  NANDX1 G30327 (.A1(W19351), .A2(W11589), .ZN(W23123));
  NANDX1 G30328 (.A1(W10855), .A2(W5642), .ZN(O486));
  NANDX1 G30329 (.A1(W22634), .A2(W15156), .ZN(O2701));
  NANDX1 G30330 (.A1(W2425), .A2(W8133), .ZN(W10588));
  NANDX1 G30331 (.A1(W8911), .A2(I1222), .ZN(W11154));
  NANDX1 G30332 (.A1(W13037), .A2(W15862), .ZN(O2702));
  NANDX1 G30333 (.A1(I1260), .A2(I1261), .ZN(W630));
  NANDX1 G30334 (.A1(W12385), .A2(I1644), .ZN(W23191));
  NANDX1 G30335 (.A1(I1392), .A2(W490), .ZN(W1477));
  NANDX1 G30336 (.A1(W18244), .A2(W13537), .ZN(W23194));
  NANDX1 G30337 (.A1(W11763), .A2(W11863), .ZN(W24483));
  NANDX1 G30338 (.A1(I956), .A2(W7065), .ZN(W10590));
  NANDX1 G30339 (.A1(W3786), .A2(W23111), .ZN(O2704));
  NANDX1 G30340 (.A1(I1262), .A2(I1263), .ZN(W631));
  NANDX1 G30341 (.A1(W833), .A2(W188), .ZN(W1476));
  NANDX1 G30342 (.A1(W22962), .A2(W14833), .ZN(W23199));
  NANDX1 G30343 (.A1(W12129), .A2(W266), .ZN(W24479));
  NANDX1 G30344 (.A1(W7311), .A2(W2206), .ZN(W11155));
  NANDX1 G30345 (.A1(W1904), .A2(W3093), .ZN(W9567));
  NANDX1 G30346 (.A1(W9337), .A2(W4475), .ZN(W11148));
  NANDX1 G30347 (.A1(W5857), .A2(W129), .ZN(O2708));
  NANDX1 G30348 (.A1(I1793), .A2(W18274), .ZN(W23208));
  NANDX1 G30349 (.A1(I241), .A2(W1273), .ZN(W1470));
  NANDX1 G30350 (.A1(I1006), .A2(I1988), .ZN(W1468));
  NANDX1 G30351 (.A1(W16438), .A2(W9025), .ZN(W23211));
  NANDX1 G30352 (.A1(W2752), .A2(W5223), .ZN(O341));
  NANDX1 G30353 (.A1(W918), .A2(W471), .ZN(W1466));
  NANDX1 G30354 (.A1(W13428), .A2(W17596), .ZN(W23218));
  NANDX1 G30355 (.A1(W6359), .A2(W5499), .ZN(W9569));
  NANDX1 G30356 (.A1(W266), .A2(I1582), .ZN(W1463));
  NANDX1 G30357 (.A1(W7638), .A2(W20700), .ZN(W23224));
  NANDX1 G30358 (.A1(I1446), .A2(I1782), .ZN(W9570));
  NANDX1 G30359 (.A1(I1260), .A2(W4060), .ZN(W11171));
  NANDX1 G30360 (.A1(W2291), .A2(W3170), .ZN(W11186));
  NANDX1 G30361 (.A1(W4293), .A2(W15263), .ZN(W23165));
  NANDX1 G30362 (.A1(W1211), .A2(I567), .ZN(W10583));
  NANDX1 G30363 (.A1(I991), .A2(I1426), .ZN(W1497));
  NANDX1 G30364 (.A1(W1317), .A2(W320), .ZN(W1495));
  NANDX1 G30365 (.A1(W4995), .A2(W6668), .ZN(W9937));
  NANDX1 G30366 (.A1(W10345), .A2(I200), .ZN(W10585));
  NANDX1 G30367 (.A1(W8934), .A2(W22994), .ZN(O3098));
  NANDX1 G30368 (.A1(I624), .A2(I61), .ZN(W1493));
  NANDX1 G30369 (.A1(W4361), .A2(W7724), .ZN(W9559));
  NANDX1 G30370 (.A1(W3568), .A2(W13443), .ZN(W23169));
  NANDX1 G30371 (.A1(I1250), .A2(I1251), .ZN(W625));
  NANDX1 G30372 (.A1(W8222), .A2(W1599), .ZN(W11183));
  NANDX1 G30373 (.A1(W2407), .A2(W2478), .ZN(W9561));
  NANDX1 G30374 (.A1(W8429), .A2(I1604), .ZN(W11172));
  NANDX1 G30375 (.A1(I1640), .A2(I174), .ZN(W1532));
  NANDX1 G30376 (.A1(W17), .A2(I1854), .ZN(W1488));
  NANDX1 G30377 (.A1(I1590), .A2(I1536), .ZN(W1486));
  NANDX1 G30378 (.A1(W424), .A2(I1912), .ZN(W1485));
  NANDX1 G30379 (.A1(W19745), .A2(W20415), .ZN(W23176));
  NANDX1 G30380 (.A1(W2834), .A2(W4395), .ZN(W9562));
  NANDX1 G30381 (.A1(W12365), .A2(W4603), .ZN(W23177));
  NANDX1 G30382 (.A1(I1258), .A2(I1259), .ZN(W629));
  NANDX1 G30383 (.A1(I1175), .A2(W9432), .ZN(O299));
  NANDX1 G30384 (.A1(W137), .A2(W713), .ZN(W1480));
  NANDX1 G30385 (.A1(W676), .A2(W4572), .ZN(W9564));
  NANDX1 G30386 (.A1(W9547), .A2(W5821), .ZN(W23184));
  NANDX1 G30387 (.A1(W5667), .A2(W10345), .ZN(W10586));
  NANDX1 G30388 (.A1(W19954), .A2(W20072), .ZN(W23185));
  NANDX1 G30389 (.A1(W7523), .A2(W6912), .ZN(W9936));
  NANDX1 G30390 (.A1(W5829), .A2(W6014), .ZN(O492));
  NANDX1 G30391 (.A1(W4593), .A2(W18750), .ZN(O2661));
  NANDX1 G30392 (.A1(I1156), .A2(I1157), .ZN(W578));
  NANDX1 G30393 (.A1(W4523), .A2(W13664), .ZN(W24537));
  NANDX1 G30394 (.A1(W17563), .A2(W18634), .ZN(W24536));
  NANDX1 G30395 (.A1(W7500), .A2(W7939), .ZN(W9498));
  NANDX1 G30396 (.A1(W20995), .A2(W9446), .ZN(O2663));
  NANDX1 G30397 (.A1(W6061), .A2(W8189), .ZN(W9500));
  NANDX1 G30398 (.A1(I692), .A2(W4296), .ZN(W23026));
  NANDX1 G30399 (.A1(W1352), .A2(W40), .ZN(W1582));
  NANDX1 G30400 (.A1(W275), .A2(I210), .ZN(W1581));
  NANDX1 G30401 (.A1(W10889), .A2(W13380), .ZN(W23027));
  NANDX1 G30402 (.A1(W6019), .A2(I1841), .ZN(W9501));
  NANDX1 G30403 (.A1(I1004), .A2(I463), .ZN(W1578));
  NANDX1 G30404 (.A1(W9955), .A2(W14183), .ZN(W23029));
  NANDX1 G30405 (.A1(W8148), .A2(W9264), .ZN(W23030));
  NANDX1 G30406 (.A1(I932), .A2(I637), .ZN(W1586));
  NANDX1 G30407 (.A1(I1158), .A2(I1159), .ZN(W579));
  NANDX1 G30408 (.A1(W5528), .A2(W10588), .ZN(W11246));
  NANDX1 G30409 (.A1(W1691), .A2(W11436), .ZN(W23031));
  NANDX1 G30410 (.A1(W5386), .A2(W23034), .ZN(W24535));
  NANDX1 G30411 (.A1(I510), .A2(W3383), .ZN(W11245));
  NANDX1 G30412 (.A1(W1672), .A2(W5784), .ZN(W11244));
  NANDX1 G30413 (.A1(W4360), .A2(W1490), .ZN(O343));
  NANDX1 G30414 (.A1(W10940), .A2(W21317), .ZN(W24533));
  NANDX1 G30415 (.A1(W8971), .A2(W19511), .ZN(W23034));
  NANDX1 G30416 (.A1(W6951), .A2(W7551), .ZN(O2665));
  NANDX1 G30417 (.A1(I1174), .A2(I1175), .ZN(W587));
  NANDX1 G30418 (.A1(W14638), .A2(W20283), .ZN(O2667));
  NANDX1 G30419 (.A1(I1176), .A2(I1177), .ZN(W588));
  NANDX1 G30420 (.A1(I1178), .A2(I1179), .ZN(W589));
  NANDX1 G30421 (.A1(I1146), .A2(I1147), .ZN(W573));
  NANDX1 G30422 (.A1(W4275), .A2(W4219), .ZN(W9960));
  NANDX1 G30423 (.A1(W10850), .A2(W10013), .ZN(W11265));
  NANDX1 G30424 (.A1(W1429), .A2(I698), .ZN(W1596));
  NANDX1 G30425 (.A1(W744), .A2(W20624), .ZN(W22996));
  NANDX1 G30426 (.A1(I1051), .A2(I163), .ZN(W9488));
  NANDX1 G30427 (.A1(W4849), .A2(W5965), .ZN(W11263));
  NANDX1 G30428 (.A1(W5379), .A2(I1844), .ZN(W9489));
  NANDX1 G30429 (.A1(W18526), .A2(W4526), .ZN(W23002));
  NANDX1 G30430 (.A1(W7318), .A2(W3105), .ZN(W9490));
  NANDX1 G30431 (.A1(W15222), .A2(W436), .ZN(W23006));
  NANDX1 G30432 (.A1(W22037), .A2(W5457), .ZN(W23007));
  NANDX1 G30433 (.A1(I1140), .A2(I1141), .ZN(W570));
  NANDX1 G30434 (.A1(I1142), .A2(I1143), .ZN(W571));
  NANDX1 G30435 (.A1(W219), .A2(W5170), .ZN(W11258));
  NANDX1 G30436 (.A1(I339), .A2(W1539), .ZN(W1593));
  NANDX1 G30437 (.A1(W2356), .A2(W5420), .ZN(W9504));
  NANDX1 G30438 (.A1(W8409), .A2(W22964), .ZN(W23014));
  NANDX1 G30439 (.A1(I1152), .A2(I1153), .ZN(W576));
  NANDX1 G30440 (.A1(W6638), .A2(W6583), .ZN(W11255));
  NANDX1 G30441 (.A1(W5049), .A2(W8892), .ZN(W9494));
  NANDX1 G30442 (.A1(I808), .A2(W6187), .ZN(W10564));
  NANDX1 G30443 (.A1(W6478), .A2(W5984), .ZN(W23017));
  NANDX1 G30444 (.A1(W3386), .A2(W3266), .ZN(W11253));
  NANDX1 G30445 (.A1(W49), .A2(I1312), .ZN(W1591));
  NANDX1 G30446 (.A1(I1429), .A2(W8241), .ZN(W11251));
  NANDX1 G30447 (.A1(W24251), .A2(W23752), .ZN(W24544));
  NANDX1 G30448 (.A1(W8987), .A2(W5038), .ZN(W9956));
  NANDX1 G30449 (.A1(W6823), .A2(W8496), .ZN(W9495));
  NANDX1 G30450 (.A1(W15604), .A2(W18712), .ZN(W23021));
  NANDX1 G30451 (.A1(W16364), .A2(W13329), .ZN(W24542));
  NANDX1 G30452 (.A1(I1192), .A2(I1193), .ZN(W596));
  NANDX1 G30453 (.A1(W3772), .A2(W11574), .ZN(W23068));
  NANDX1 G30454 (.A1(I1834), .A2(W9340), .ZN(W9516));
  NANDX1 G30455 (.A1(W8545), .A2(I1702), .ZN(W11226));
  NANDX1 G30456 (.A1(I811), .A2(W9000), .ZN(W9517));
  NANDX1 G30457 (.A1(I817), .A2(W609), .ZN(W1549));
  NANDX1 G30458 (.A1(I1188), .A2(I1189), .ZN(W594));
  NANDX1 G30459 (.A1(W7977), .A2(W1689), .ZN(W9518));
  NANDX1 G30460 (.A1(I760), .A2(I771), .ZN(W1543));
  NANDX1 G30461 (.A1(W9095), .A2(W3159), .ZN(W9520));
  NANDX1 G30462 (.A1(W6538), .A2(W17690), .ZN(W23078));
  NANDX1 G30463 (.A1(W14651), .A2(W1042), .ZN(W23079));
  NANDX1 G30464 (.A1(W23185), .A2(W7500), .ZN(W24514));
  NANDX1 G30465 (.A1(W472), .A2(W481), .ZN(W1541));
  NANDX1 G30466 (.A1(W8250), .A2(W6374), .ZN(W23081));
  NANDX1 G30467 (.A1(W631), .A2(W695), .ZN(W1539));
  NANDX1 G30468 (.A1(I1186), .A2(I1187), .ZN(W593));
  NANDX1 G30469 (.A1(W4874), .A2(W2162), .ZN(W23083));
  NANDX1 G30470 (.A1(W12022), .A2(W10904), .ZN(O2674));
  NANDX1 G30471 (.A1(W6429), .A2(W6960), .ZN(W9524));
  NANDX1 G30472 (.A1(W7314), .A2(W398), .ZN(W9525));
  NANDX1 G30473 (.A1(I1196), .A2(I1197), .ZN(W598));
  NANDX1 G30474 (.A1(W17957), .A2(W19964), .ZN(W23087));
  NANDX1 G30475 (.A1(W20572), .A2(W12618), .ZN(W23089));
  NANDX1 G30476 (.A1(W6118), .A2(W6036), .ZN(W10574));
  NANDX1 G30477 (.A1(I1198), .A2(I1199), .ZN(W599));
  NANDX1 G30478 (.A1(W13437), .A2(W21400), .ZN(W23091));
  NANDX1 G30479 (.A1(W9486), .A2(W499), .ZN(W23094));
  NANDX1 G30480 (.A1(W595), .A2(I142), .ZN(W1534));
  NANDX1 G30481 (.A1(I1200), .A2(I1201), .ZN(W600));
  NANDX1 G30482 (.A1(W4502), .A2(W4392), .ZN(W24511));
  NANDX1 G30483 (.A1(W228), .A2(W19828), .ZN(W23056));
  NANDX1 G30484 (.A1(W15734), .A2(W14384), .ZN(W23042));
  NANDX1 G30485 (.A1(W10023), .A2(W6181), .ZN(W23045));
  NANDX1 G30486 (.A1(I1180), .A2(I1181), .ZN(W590));
  NANDX1 G30487 (.A1(W6248), .A2(W3832), .ZN(W9508));
  NANDX1 G30488 (.A1(W7924), .A2(W14553), .ZN(O2669));
  NANDX1 G30489 (.A1(W10822), .A2(W19967), .ZN(W23048));
  NANDX1 G30490 (.A1(W8385), .A2(W1164), .ZN(W23051));
  NANDX1 G30491 (.A1(I1024), .A2(I1653), .ZN(W1565));
  NANDX1 G30492 (.A1(W7300), .A2(I1381), .ZN(W11237));
  NANDX1 G30493 (.A1(I1157), .A2(W8363), .ZN(W23053));
  NANDX1 G30494 (.A1(W1801), .A2(W8430), .ZN(W9509));
  NANDX1 G30495 (.A1(I441), .A2(I1103), .ZN(W1564));
  NANDX1 G30496 (.A1(W4521), .A2(W1397), .ZN(O3109));
  NANDX1 G30497 (.A1(W1490), .A2(W2395), .ZN(W24527));
  NANDX1 G30498 (.A1(W631), .A2(W1699), .ZN(W1775));
  NANDX1 G30499 (.A1(W7815), .A2(W943), .ZN(W9512));
  NANDX1 G30500 (.A1(W1544), .A2(W279), .ZN(W1562));
  NANDX1 G30501 (.A1(W5433), .A2(W13773), .ZN(W23058));
  NANDX1 G30502 (.A1(W7340), .A2(W7955), .ZN(W10571));
  NANDX1 G30503 (.A1(W6441), .A2(W498), .ZN(W9514));
  NANDX1 G30504 (.A1(W1418), .A2(I874), .ZN(W1557));
  NANDX1 G30505 (.A1(I371), .A2(I1795), .ZN(W1556));
  NANDX1 G30506 (.A1(W5945), .A2(W6899), .ZN(W11232));
  NANDX1 G30507 (.A1(W15564), .A2(W6265), .ZN(W24522));
  NANDX1 G30508 (.A1(W17024), .A2(I1158), .ZN(O2672));
  NANDX1 G30509 (.A1(I1819), .A2(I1944), .ZN(W1554));
  NANDX1 G30510 (.A1(W993), .A2(I539), .ZN(W1552));
  NANDX1 G30511 (.A1(W6431), .A2(W1581), .ZN(W9515));
  NANDX1 G30512 (.A1(W21831), .A2(W11763), .ZN(O3107));
  NANDX1 G30513 (.A1(W5357), .A2(W15404), .ZN(O2517));
  NANDX1 G30514 (.A1(W5917), .A2(W7533), .ZN(W9318));
  NANDX1 G30515 (.A1(W7247), .A2(W5626), .ZN(W10481));
  NANDX1 G30516 (.A1(I820), .A2(I821), .ZN(W410));
  NANDX1 G30517 (.A1(W8443), .A2(W992), .ZN(W10483));
  NANDX1 G30518 (.A1(I565), .A2(W1493), .ZN(W1983));
  NANDX1 G30519 (.A1(W4219), .A2(I1884), .ZN(W10007));
  NANDX1 G30520 (.A1(W10852), .A2(W22620), .ZN(O3181));
  NANDX1 G30521 (.A1(W23017), .A2(W5350), .ZN(O3179));
  NANDX1 G30522 (.A1(I826), .A2(I827), .ZN(W413));
  NANDX1 G30523 (.A1(W10905), .A2(W3177), .ZN(O3178));
  NANDX1 G30524 (.A1(I828), .A2(I829), .ZN(W414));
  NANDX1 G30525 (.A1(I884), .A2(I1914), .ZN(W1978));
  NANDX1 G30526 (.A1(W11019), .A2(W7905), .ZN(W11505));
  NANDX1 G30527 (.A1(I1943), .A2(W5871), .ZN(W9325));
  NANDX1 G30528 (.A1(I1957), .A2(I1956), .ZN(W1977));
  NANDX1 G30529 (.A1(I812), .A2(I813), .ZN(W406));
  NANDX1 G30530 (.A1(W6322), .A2(W7455), .ZN(W22448));
  NANDX1 G30531 (.A1(I713), .A2(W9116), .ZN(O283));
  NANDX1 G30532 (.A1(W1634), .A2(I580), .ZN(W1975));
  NANDX1 G30533 (.A1(W1595), .A2(W1849), .ZN(W11503));
  NANDX1 G30534 (.A1(W2290), .A2(W4824), .ZN(W9327));
  NANDX1 G30535 (.A1(W2648), .A2(I1373), .ZN(W9328));
  NANDX1 G30536 (.A1(W1388), .A2(W654), .ZN(W1969));
  NANDX1 G30537 (.A1(W9587), .A2(W14130), .ZN(O2520));
  NANDX1 G30538 (.A1(W5517), .A2(W4112), .ZN(W10004));
  NANDX1 G30539 (.A1(I558), .A2(W12594), .ZN(W22462));
  NANDX1 G30540 (.A1(W8576), .A2(W20894), .ZN(W22465));
  NANDX1 G30541 (.A1(W22184), .A2(W5183), .ZN(O2521));
  NANDX1 G30542 (.A1(W6944), .A2(W6295), .ZN(W11502));
  NANDX1 G30543 (.A1(W3319), .A2(W21108), .ZN(W22469));
  NANDX1 G30544 (.A1(W20434), .A2(W11479), .ZN(W22430));
  NANDX1 G30545 (.A1(W2309), .A2(W21313), .ZN(O2505));
  NANDX1 G30546 (.A1(W159), .A2(W2866), .ZN(W9303));
  NANDX1 G30547 (.A1(W2318), .A2(W1311), .ZN(W9304));
  NANDX1 G30548 (.A1(W15124), .A2(W12354), .ZN(O2507));
  NANDX1 G30549 (.A1(W12594), .A2(W8570), .ZN(O2508));
  NANDX1 G30550 (.A1(W3845), .A2(W1535), .ZN(O2509));
  NANDX1 G30551 (.A1(W2014), .A2(W6970), .ZN(W9306));
  NANDX1 G30552 (.A1(W4426), .A2(I906), .ZN(W10476));
  NANDX1 G30553 (.A1(W2028), .A2(I1672), .ZN(W11515));
  NANDX1 G30554 (.A1(W5430), .A2(W3400), .ZN(W9308));
  NANDX1 G30555 (.A1(W3075), .A2(I1912), .ZN(W10477));
  NANDX1 G30556 (.A1(W14221), .A2(W1282), .ZN(W22425));
  NANDX1 G30557 (.A1(I1718), .A2(W1249), .ZN(O16));
  NANDX1 G30558 (.A1(W7417), .A2(W2999), .ZN(W22427));
  NANDX1 G30559 (.A1(W16018), .A2(W14549), .ZN(W22428));
  NANDX1 G30560 (.A1(W11976), .A2(W15049), .ZN(W22470));
  NANDX1 G30561 (.A1(W2622), .A2(W20872), .ZN(W22431));
  NANDX1 G30562 (.A1(W2430), .A2(W10713), .ZN(W11514));
  NANDX1 G30563 (.A1(W17739), .A2(I1300), .ZN(O2512));
  NANDX1 G30564 (.A1(W8947), .A2(W9561), .ZN(W10478));
  NANDX1 G30565 (.A1(W1785), .A2(I659), .ZN(W1992));
  NANDX1 G30566 (.A1(W770), .A2(W1460), .ZN(W1991));
  NANDX1 G30567 (.A1(W870), .A2(W7901), .ZN(W9313));
  NANDX1 G30568 (.A1(W1534), .A2(W439), .ZN(W1990));
  NANDX1 G30569 (.A1(W11639), .A2(W8398), .ZN(W22434));
  NANDX1 G30570 (.A1(W9900), .A2(W7907), .ZN(W22435));
  NANDX1 G30571 (.A1(W9088), .A2(W2520), .ZN(W10479));
  NANDX1 G30572 (.A1(W1760), .A2(I111), .ZN(W1987));
  NANDX1 G30573 (.A1(I810), .A2(I811), .ZN(W405));
  NANDX1 G30574 (.A1(I1832), .A2(W8163), .ZN(W11511));
  NANDX1 G30575 (.A1(W282), .A2(I366), .ZN(W1935));
  NANDX1 G30576 (.A1(W7860), .A2(I450), .ZN(W10488));
  NANDX1 G30577 (.A1(W5010), .A2(W9271), .ZN(O514));
  NANDX1 G30578 (.A1(W4347), .A2(W16236), .ZN(O3174));
  NANDX1 G30579 (.A1(W3262), .A2(W3054), .ZN(W9337));
  NANDX1 G30580 (.A1(I416), .A2(W1451), .ZN(W9338));
  NANDX1 G30581 (.A1(W16514), .A2(W18210), .ZN(W22512));
  NANDX1 G30582 (.A1(W1348), .A2(W284), .ZN(W1941));
  NANDX1 G30583 (.A1(W8747), .A2(W10134), .ZN(W10489));
  NANDX1 G30584 (.A1(W6868), .A2(W4786), .ZN(W11475));
  NANDX1 G30585 (.A1(W4350), .A2(W15814), .ZN(W24729));
  NANDX1 G30586 (.A1(W1565), .A2(W1216), .ZN(O2540));
  NANDX1 G30587 (.A1(W5059), .A2(I498), .ZN(O2541));
  NANDX1 G30588 (.A1(I200), .A2(W5377), .ZN(W9341));
  NANDX1 G30589 (.A1(W1248), .A2(W2494), .ZN(W22522));
  NANDX1 G30590 (.A1(I115), .A2(I538), .ZN(W1936));
  NANDX1 G30591 (.A1(W9738), .A2(W13174), .ZN(O2535));
  NANDX1 G30592 (.A1(W11981), .A2(W2326), .ZN(W22531));
  NANDX1 G30593 (.A1(W1236), .A2(W3229), .ZN(W11470));
  NANDX1 G30594 (.A1(W5010), .A2(W5623), .ZN(W11469));
  NANDX1 G30595 (.A1(W10355), .A2(W3286), .ZN(W11466));
  NANDX1 G30596 (.A1(W20277), .A2(W10200), .ZN(W22535));
  NANDX1 G30597 (.A1(W14358), .A2(W17622), .ZN(W22536));
  NANDX1 G30598 (.A1(W6527), .A2(W9776), .ZN(W22537));
  NANDX1 G30599 (.A1(I1464), .A2(W1851), .ZN(W11465));
  NANDX1 G30600 (.A1(I1168), .A2(W1056), .ZN(W1929));
  NANDX1 G30601 (.A1(W5029), .A2(W14863), .ZN(W22542));
  NANDX1 G30602 (.A1(W5790), .A2(W16181), .ZN(W22543));
  NANDX1 G30603 (.A1(W2315), .A2(W14527), .ZN(O3173));
  NANDX1 G30604 (.A1(W748), .A2(W1509), .ZN(W1928));
  NANDX1 G30605 (.A1(W3700), .A2(W10116), .ZN(W11464));
  NANDX1 G30606 (.A1(I1346), .A2(I316), .ZN(W1954));
  NANDX1 G30607 (.A1(W46), .A2(W1085), .ZN(W1966));
  NANDX1 G30608 (.A1(W14), .A2(I1214), .ZN(W1964));
  NANDX1 G30609 (.A1(W12634), .A2(W4087), .ZN(O2527));
  NANDX1 G30610 (.A1(W7483), .A2(W20671), .ZN(O3177));
  NANDX1 G30611 (.A1(W1507), .A2(W3879), .ZN(W10002));
  NANDX1 G30612 (.A1(I842), .A2(I843), .ZN(W421));
  NANDX1 G30613 (.A1(W9928), .A2(I991), .ZN(W11497));
  NANDX1 G30614 (.A1(I1022), .A2(W45), .ZN(O515));
  NANDX1 G30615 (.A1(W7223), .A2(W10480), .ZN(W11495));
  NANDX1 G30616 (.A1(W17161), .A2(W3758), .ZN(O2529));
  NANDX1 G30617 (.A1(W5791), .A2(W9447), .ZN(W10485));
  NANDX1 G30618 (.A1(I1167), .A2(W4048), .ZN(W11492));
  NANDX1 G30619 (.A1(W601), .A2(W3207), .ZN(W11490));
  NANDX1 G30620 (.A1(I1261), .A2(I1442), .ZN(W1956));
  NANDX1 G30621 (.A1(I42), .A2(W6616), .ZN(W24738));
  NANDX1 G30622 (.A1(W730), .A2(I850), .ZN(W1996));
  NANDX1 G30623 (.A1(W8036), .A2(W2809), .ZN(W22486));
  NANDX1 G30624 (.A1(I1232), .A2(W8554), .ZN(W11487));
  NANDX1 G30625 (.A1(W1565), .A2(W3716), .ZN(W11486));
  NANDX1 G30626 (.A1(W12543), .A2(W10528), .ZN(W22491));
  NANDX1 G30627 (.A1(W3074), .A2(W8001), .ZN(W10486));
  NANDX1 G30628 (.A1(W164), .A2(W1415), .ZN(W1949));
  NANDX1 G30629 (.A1(W793), .A2(W1890), .ZN(W22494));
  NANDX1 G30630 (.A1(I848), .A2(I849), .ZN(W424));
  NANDX1 G30631 (.A1(W24279), .A2(W12581), .ZN(W24733));
  NANDX1 G30632 (.A1(W19071), .A2(W17700), .ZN(W24731));
  NANDX1 G30633 (.A1(W1313), .A2(W727), .ZN(W10487));
  NANDX1 G30634 (.A1(W825), .A2(W329), .ZN(W1948));
  NANDX1 G30635 (.A1(I1439), .A2(I400), .ZN(W11484));
  NANDX1 G30636 (.A1(W13021), .A2(W12042), .ZN(W22500));
  NANDX1 G30637 (.A1(W5997), .A2(W5693), .ZN(W11560));
  NANDX1 G30638 (.A1(W5458), .A2(W2410), .ZN(W11569));
  NANDX1 G30639 (.A1(I758), .A2(I759), .ZN(W379));
  NANDX1 G30640 (.A1(W470), .A2(W111), .ZN(W9270));
  NANDX1 G30641 (.A1(I75), .A2(W12742), .ZN(O2485));
  NANDX1 G30642 (.A1(W11182), .A2(W12444), .ZN(W22345));
  NANDX1 G30643 (.A1(W1825), .A2(W4967), .ZN(W10018));
  NANDX1 G30644 (.A1(W17896), .A2(W942), .ZN(O2486));
  NANDX1 G30645 (.A1(W928), .A2(W2514), .ZN(W22349));
  NANDX1 G30646 (.A1(W12075), .A2(W1987), .ZN(O2487));
  NANDX1 G30647 (.A1(W12599), .A2(I117), .ZN(W22351));
  NANDX1 G30648 (.A1(W9308), .A2(W5083), .ZN(W11564));
  NANDX1 G30649 (.A1(W327), .A2(I1725), .ZN(W2061));
  NANDX1 G30650 (.A1(I1919), .A2(I995), .ZN(W2060));
  NANDX1 G30651 (.A1(I296), .A2(W7982), .ZN(W10456));
  NANDX1 G30652 (.A1(W3804), .A2(W8614), .ZN(W24780));
  NANDX1 G30653 (.A1(W6350), .A2(W20372), .ZN(O3192));
  NANDX1 G30654 (.A1(W10634), .A2(W9083), .ZN(W11558));
  NANDX1 G30655 (.A1(W4819), .A2(W17416), .ZN(W22357));
  NANDX1 G30656 (.A1(W3621), .A2(I1264), .ZN(W11557));
  NANDX1 G30657 (.A1(W2047), .A2(W14912), .ZN(W22358));
  NANDX1 G30658 (.A1(W12497), .A2(W6405), .ZN(O3191));
  NANDX1 G30659 (.A1(W6668), .A2(W3873), .ZN(O394));
  NANDX1 G30660 (.A1(W11248), .A2(W1363), .ZN(O520));
  NANDX1 G30661 (.A1(W1256), .A2(I1921), .ZN(W2055));
  NANDX1 G30662 (.A1(W9615), .A2(W4488), .ZN(W22362));
  NANDX1 G30663 (.A1(W10450), .A2(W8253), .ZN(W24776));
  NANDX1 G30664 (.A1(I770), .A2(I771), .ZN(W385));
  NANDX1 G30665 (.A1(W81), .A2(I980), .ZN(W2053));
  NANDX1 G30666 (.A1(W7901), .A2(W7013), .ZN(W11551));
  NANDX1 G30667 (.A1(I772), .A2(I773), .ZN(W386));
  NANDX1 G30668 (.A1(I1182), .A2(W6491), .ZN(W22328));
  NANDX1 G30669 (.A1(I1656), .A2(I319), .ZN(W2077));
  NANDX1 G30670 (.A1(W13102), .A2(W13070), .ZN(W22316));
  NANDX1 G30671 (.A1(W6723), .A2(W5578), .ZN(W22318));
  NANDX1 G30672 (.A1(I1538), .A2(I40), .ZN(W2075));
  NANDX1 G30673 (.A1(W1010), .A2(W1082), .ZN(W2074));
  NANDX1 G30674 (.A1(I1240), .A2(W724), .ZN(W11580));
  NANDX1 G30675 (.A1(W10), .A2(W9929), .ZN(W24788));
  NANDX1 G30676 (.A1(I5), .A2(W1581), .ZN(W11578));
  NANDX1 G30677 (.A1(W18575), .A2(W21652), .ZN(W22320));
  NANDX1 G30678 (.A1(I915), .A2(W1087), .ZN(W11577));
  NANDX1 G30679 (.A1(I432), .A2(I0), .ZN(O2482));
  NANDX1 G30680 (.A1(W135), .A2(W18898), .ZN(W22324));
  NANDX1 G30681 (.A1(W21083), .A2(W14578), .ZN(W22326));
  NANDX1 G30682 (.A1(W8821), .A2(W16549), .ZN(W24787));
  NANDX1 G30683 (.A1(W15078), .A2(W20441), .ZN(W22327));
  NANDX1 G30684 (.A1(W14766), .A2(W22329), .ZN(W24772));
  NANDX1 G30685 (.A1(W4910), .A2(W7365), .ZN(W9264));
  NANDX1 G30686 (.A1(W21276), .A2(W8824), .ZN(W22330));
  NANDX1 G30687 (.A1(I1703), .A2(W10860), .ZN(W11572));
  NANDX1 G30688 (.A1(W842), .A2(W11380), .ZN(W22333));
  NANDX1 G30689 (.A1(W16697), .A2(W7410), .ZN(W22335));
  NANDX1 G30690 (.A1(W4450), .A2(W13718), .ZN(W22336));
  NANDX1 G30691 (.A1(I754), .A2(I755), .ZN(W377));
  NANDX1 G30692 (.A1(W9370), .A2(W3774), .ZN(W10449));
  NANDX1 G30693 (.A1(W5228), .A2(W13339), .ZN(W22337));
  NANDX1 G30694 (.A1(W9963), .A2(W3246), .ZN(W10450));
  NANDX1 G30695 (.A1(W21817), .A2(W5360), .ZN(W22339));
  NANDX1 G30696 (.A1(W1293), .A2(W2115), .ZN(W9267));
  NANDX1 G30697 (.A1(W21792), .A2(W23423), .ZN(O3193));
  NANDX1 G30698 (.A1(W10012), .A2(I1165), .ZN(W22340));
  NANDX1 G30699 (.A1(W1709), .A2(W8718), .ZN(O2499));
  NANDX1 G30700 (.A1(W11324), .A2(W9479), .ZN(W24763));
  NANDX1 G30701 (.A1(I980), .A2(W15632), .ZN(O2497));
  NANDX1 G30702 (.A1(W55), .A2(W15048), .ZN(W22393));
  NANDX1 G30703 (.A1(W1998), .A2(W1930), .ZN(W2020));
  NANDX1 G30704 (.A1(W4713), .A2(I1708), .ZN(W11527));
  NANDX1 G30705 (.A1(I913), .A2(W1888), .ZN(W2018));
  NANDX1 G30706 (.A1(W4751), .A2(W13155), .ZN(W22395));
  NANDX1 G30707 (.A1(W421), .A2(I400), .ZN(W2017));
  NANDX1 G30708 (.A1(I214), .A2(W284), .ZN(W2015));
  NANDX1 G30709 (.A1(W1271), .A2(W463), .ZN(W9294));
  NANDX1 G30710 (.A1(I796), .A2(I797), .ZN(W398));
  NANDX1 G30711 (.A1(W16499), .A2(W16979), .ZN(W22398));
  NANDX1 G30712 (.A1(I284), .A2(W389), .ZN(W2013));
  NANDX1 G30713 (.A1(W922), .A2(W1370), .ZN(W2012));
  NANDX1 G30714 (.A1(W6917), .A2(W20986), .ZN(O3187));
  NANDX1 G30715 (.A1(W8924), .A2(W11547), .ZN(W22391));
  NANDX1 G30716 (.A1(W14298), .A2(W4066), .ZN(O2500));
  NANDX1 G30717 (.A1(W1284), .A2(I558), .ZN(W2010));
  NANDX1 G30718 (.A1(I798), .A2(I799), .ZN(W399));
  NANDX1 G30719 (.A1(W8355), .A2(W4372), .ZN(O352));
  NANDX1 G30720 (.A1(W6663), .A2(W6632), .ZN(W22404));
  NANDX1 G30721 (.A1(I290), .A2(I1730), .ZN(W2007));
  NANDX1 G30722 (.A1(W9887), .A2(W15084), .ZN(W22405));
  NANDX1 G30723 (.A1(W1386), .A2(W1616), .ZN(W2005));
  NANDX1 G30724 (.A1(W6376), .A2(W9116), .ZN(W11522));
  NANDX1 G30725 (.A1(W9712), .A2(W289), .ZN(W11519));
  NANDX1 G30726 (.A1(W1366), .A2(I250), .ZN(W1999));
  NANDX1 G30727 (.A1(W7058), .A2(W7658), .ZN(W10475));
  NANDX1 G30728 (.A1(W22154), .A2(I839), .ZN(W22412));
  NANDX1 G30729 (.A1(I887), .A2(I914), .ZN(W1997));
  NANDX1 G30730 (.A1(W22052), .A2(W13107), .ZN(O2494));
  NANDX1 G30731 (.A1(W10949), .A2(W9362), .ZN(W22368));
  NANDX1 G30732 (.A1(W1475), .A2(W3305), .ZN(W11546));
  NANDX1 G30733 (.A1(W3417), .A2(W1296), .ZN(W22371));
  NANDX1 G30734 (.A1(W734), .A2(W1419), .ZN(W2047));
  NANDX1 G30735 (.A1(W2336), .A2(W5952), .ZN(O517));
  NANDX1 G30736 (.A1(I1942), .A2(W2954), .ZN(W10016));
  NANDX1 G30737 (.A1(W125), .A2(W11457), .ZN(W11542));
  NANDX1 G30738 (.A1(I1008), .A2(W64), .ZN(W22373));
  NANDX1 G30739 (.A1(W8629), .A2(W11383), .ZN(W11541));
  NANDX1 G30740 (.A1(W10198), .A2(W7152), .ZN(W10465));
  NANDX1 G30741 (.A1(W6957), .A2(W2460), .ZN(W9286));
  NANDX1 G30742 (.A1(W3493), .A2(I1143), .ZN(W10013));
  NANDX1 G30743 (.A1(I564), .A2(W642), .ZN(W2034));
  NANDX1 G30744 (.A1(W1273), .A2(W17377), .ZN(O2492));
  NANDX1 G30745 (.A1(W23328), .A2(W8735), .ZN(O3188));
  NANDX1 G30746 (.A1(W1643), .A2(W6255), .ZN(W9343));
  NANDX1 G30747 (.A1(W319), .A2(I490), .ZN(W2032));
  NANDX1 G30748 (.A1(W18505), .A2(W12109), .ZN(W22382));
  NANDX1 G30749 (.A1(W1685), .A2(W5901), .ZN(W11538));
  NANDX1 G30750 (.A1(W6096), .A2(W7901), .ZN(W9287));
  NANDX1 G30751 (.A1(W6269), .A2(W6058), .ZN(W11536));
  NANDX1 G30752 (.A1(W469), .A2(I622), .ZN(W2029));
  NANDX1 G30753 (.A1(W6755), .A2(W4917), .ZN(W9288));
  NANDX1 G30754 (.A1(W5798), .A2(I1554), .ZN(W11531));
  NANDX1 G30755 (.A1(I856), .A2(W760), .ZN(W2027));
  NANDX1 G30756 (.A1(W7344), .A2(W644), .ZN(W10012));
  NANDX1 G30757 (.A1(I1504), .A2(W158), .ZN(W2022));
  NANDX1 G30758 (.A1(W7796), .A2(W668), .ZN(W9291));
  NANDX1 G30759 (.A1(W4256), .A2(W2919), .ZN(W11528));
  NANDX1 G30760 (.A1(W10420), .A2(W19441), .ZN(O2496));
  NANDX1 G30761 (.A1(W8943), .A2(W2116), .ZN(W11409));
  NANDX1 G30762 (.A1(W2097), .A2(W8168), .ZN(W11418));
  NANDX1 G30763 (.A1(I966), .A2(I967), .ZN(W483));
  NANDX1 G30764 (.A1(W1382), .A2(W393), .ZN(W22675));
  NANDX1 G30765 (.A1(I972), .A2(I973), .ZN(W486));
  NANDX1 G30766 (.A1(W9537), .A2(W8560), .ZN(W11417));
  NANDX1 G30767 (.A1(W18824), .A2(W17179), .ZN(W22676));
  NANDX1 G30768 (.A1(W1404), .A2(I1343), .ZN(W1822));
  NANDX1 G30769 (.A1(W982), .A2(W92), .ZN(W1821));
  NANDX1 G30770 (.A1(W3182), .A2(W10161), .ZN(W11416));
  NANDX1 G30771 (.A1(I1396), .A2(W5999), .ZN(W11415));
  NANDX1 G30772 (.A1(I1114), .A2(W294), .ZN(W1817));
  NANDX1 G30773 (.A1(W3465), .A2(I1997), .ZN(W9385));
  NANDX1 G30774 (.A1(W1486), .A2(W1129), .ZN(W1816));
  NANDX1 G30775 (.A1(I1563), .A2(W1769), .ZN(W1815));
  NANDX1 G30776 (.A1(W4997), .A2(W6755), .ZN(W10520));
  NANDX1 G30777 (.A1(I964), .A2(I965), .ZN(W482));
  NANDX1 G30778 (.A1(W8976), .A2(W10346), .ZN(O506));
  NANDX1 G30779 (.A1(W19610), .A2(I1825), .ZN(W22685));
  NANDX1 G30780 (.A1(W11709), .A2(W7325), .ZN(W22688));
  NANDX1 G30781 (.A1(W12637), .A2(W2321), .ZN(W22689));
  NANDX1 G30782 (.A1(W3548), .A2(W17482), .ZN(O2582));
  NANDX1 G30783 (.A1(I1962), .A2(W17515), .ZN(O3158));
  NANDX1 G30784 (.A1(I976), .A2(I977), .ZN(W488));
  NANDX1 G30785 (.A1(W1734), .A2(W6419), .ZN(W24663));
  NANDX1 G30786 (.A1(I980), .A2(I981), .ZN(W490));
  NANDX1 G30787 (.A1(W21249), .A2(W7314), .ZN(O2585));
  NANDX1 G30788 (.A1(I1958), .A2(W2172), .ZN(W9388));
  NANDX1 G30789 (.A1(W8920), .A2(W7443), .ZN(W11406));
  NANDX1 G30790 (.A1(I1098), .A2(W2920), .ZN(W9389));
  NANDX1 G30791 (.A1(I986), .A2(I987), .ZN(W493));
  NANDX1 G30792 (.A1(I1941), .A2(W1553), .ZN(W1836));
  NANDX1 G30793 (.A1(W315), .A2(W2413), .ZN(W22637));
  NANDX1 G30794 (.A1(W847), .A2(W12329), .ZN(O2562));
  NANDX1 G30795 (.A1(I598), .A2(W153), .ZN(W1845));
  NANDX1 G30796 (.A1(W7116), .A2(W640), .ZN(W10513));
  NANDX1 G30797 (.A1(I565), .A2(W1618), .ZN(W1844));
  NANDX1 G30798 (.A1(W711), .A2(I1310), .ZN(W1843));
  NANDX1 G30799 (.A1(W1655), .A2(W18123), .ZN(W22641));
  NANDX1 G30800 (.A1(W10029), .A2(W22579), .ZN(W24679));
  NANDX1 G30801 (.A1(W432), .A2(W14), .ZN(W1840));
  NANDX1 G30802 (.A1(W7930), .A2(W9670), .ZN(W22644));
  NANDX1 G30803 (.A1(W467), .A2(W661), .ZN(W1838));
  NANDX1 G30804 (.A1(I616), .A2(W21652), .ZN(W24677));
  NANDX1 G30805 (.A1(W5932), .A2(W501), .ZN(O403));
  NANDX1 G30806 (.A1(W10185), .A2(W10566), .ZN(W11427));
  NANDX1 G30807 (.A1(I18), .A2(W7158), .ZN(O285));
  NANDX1 G30808 (.A1(W24523), .A2(W18206), .ZN(W24657));
  NANDX1 G30809 (.A1(W17613), .A2(W14504), .ZN(O2569));
  NANDX1 G30810 (.A1(W15117), .A2(W22018), .ZN(O2571));
  NANDX1 G30811 (.A1(I962), .A2(I963), .ZN(W481));
  NANDX1 G30812 (.A1(W7310), .A2(W2479), .ZN(W10516));
  NANDX1 G30813 (.A1(W21158), .A2(I1717), .ZN(W24676));
  NANDX1 G30814 (.A1(W22393), .A2(W11204), .ZN(W22659));
  NANDX1 G30815 (.A1(W1473), .A2(W1469), .ZN(W1834));
  NANDX1 G30816 (.A1(W7197), .A2(W10615), .ZN(W11425));
  NANDX1 G30817 (.A1(W5), .A2(I1534), .ZN(W1831));
  NANDX1 G30818 (.A1(W6674), .A2(I255), .ZN(W9982));
  NANDX1 G30819 (.A1(W3528), .A2(W5877), .ZN(W11424));
  NANDX1 G30820 (.A1(I1755), .A2(I299), .ZN(W1830));
  NANDX1 G30821 (.A1(W21841), .A2(W20696), .ZN(O2579));
  NANDX1 G30822 (.A1(W5289), .A2(W2864), .ZN(W9383));
  NANDX1 G30823 (.A1(W8333), .A2(W11858), .ZN(O2601));
  NANDX1 G30824 (.A1(W8131), .A2(W6984), .ZN(W11395));
  NANDX1 G30825 (.A1(W11530), .A2(W1218), .ZN(O3152));
  NANDX1 G30826 (.A1(W5217), .A2(W2673), .ZN(W9405));
  NANDX1 G30827 (.A1(W869), .A2(W9849), .ZN(W11392));
  NANDX1 G30828 (.A1(W8491), .A2(W9259), .ZN(W11391));
  NANDX1 G30829 (.A1(I1032), .A2(W557), .ZN(O287));
  NANDX1 G30830 (.A1(W2077), .A2(W2206), .ZN(W9976));
  NANDX1 G30831 (.A1(W21145), .A2(W428), .ZN(W22743));
  NANDX1 G30832 (.A1(W4714), .A2(W648), .ZN(W11388));
  NANDX1 G30833 (.A1(I1004), .A2(I1005), .ZN(W502));
  NANDX1 G30834 (.A1(W7254), .A2(W18876), .ZN(W22747));
  NANDX1 G30835 (.A1(W17990), .A2(W10314), .ZN(W22749));
  NANDX1 G30836 (.A1(W496), .A2(W557), .ZN(W11387));
  NANDX1 G30837 (.A1(W13826), .A2(W18460), .ZN(O2600));
  NANDX1 G30838 (.A1(W3514), .A2(W15690), .ZN(W22752));
  NANDX1 G30839 (.A1(W18335), .A2(W17422), .ZN(O2597));
  NANDX1 G30840 (.A1(I538), .A2(I1105), .ZN(W1785));
  NANDX1 G30841 (.A1(W1210), .A2(W8083), .ZN(O504));
  NANDX1 G30842 (.A1(W4931), .A2(W1770), .ZN(W11384));
  NANDX1 G30843 (.A1(W4404), .A2(W5809), .ZN(W9975));
  NANDX1 G30844 (.A1(W187), .A2(W791), .ZN(W1782));
  NANDX1 G30845 (.A1(I1154), .A2(W8643), .ZN(W9409));
  NANDX1 G30846 (.A1(W1653), .A2(W13717), .ZN(O3151));
  NANDX1 G30847 (.A1(W5484), .A2(W9678), .ZN(W10529));
  NANDX1 G30848 (.A1(W6290), .A2(W12739), .ZN(W24635));
  NANDX1 G30849 (.A1(I1012), .A2(I1013), .ZN(W506));
  NANDX1 G30850 (.A1(W3127), .A2(W7338), .ZN(W11381));
  NANDX1 G30851 (.A1(W552), .A2(W10145), .ZN(W22759));
  NANDX1 G30852 (.A1(I898), .A2(I664), .ZN(W1776));
  NANDX1 G30853 (.A1(W109), .A2(W3137), .ZN(W11379));
  NANDX1 G30854 (.A1(W21284), .A2(W16528), .ZN(W22724));
  NANDX1 G30855 (.A1(W15707), .A2(W20391), .ZN(W22702));
  NANDX1 G30856 (.A1(W14896), .A2(W24020), .ZN(W24656));
  NANDX1 G30857 (.A1(W16982), .A2(W8639), .ZN(W22703));
  NANDX1 G30858 (.A1(W9713), .A2(W2269), .ZN(W22706));
  NANDX1 G30859 (.A1(I706), .A2(I1948), .ZN(W1804));
  NANDX1 G30860 (.A1(W10533), .A2(W996), .ZN(W11401));
  NANDX1 G30861 (.A1(W12858), .A2(W2443), .ZN(W22710));
  NANDX1 G30862 (.A1(W14015), .A2(W11638), .ZN(O2589));
  NANDX1 G30863 (.A1(W14252), .A2(W12966), .ZN(O2590));
  NANDX1 G30864 (.A1(W2690), .A2(W16235), .ZN(W22714));
  NANDX1 G30865 (.A1(I1438), .A2(I1424), .ZN(W1802));
  NANDX1 G30866 (.A1(W15957), .A2(W9926), .ZN(W22720));
  NANDX1 G30867 (.A1(I912), .A2(I1503), .ZN(W9395));
  NANDX1 G30868 (.A1(W4029), .A2(I1027), .ZN(W22723));
  NANDX1 G30869 (.A1(I992), .A2(I993), .ZN(W496));
  NANDX1 G30870 (.A1(W8946), .A2(W14852), .ZN(O2561));
  NANDX1 G30871 (.A1(I994), .A2(I995), .ZN(W497));
  NANDX1 G30872 (.A1(W14288), .A2(W9555), .ZN(O2593));
  NANDX1 G30873 (.A1(W10497), .A2(W15593), .ZN(W22729));
  NANDX1 G30874 (.A1(W15073), .A2(W11349), .ZN(W24653));
  NANDX1 G30875 (.A1(W3470), .A2(W6338), .ZN(W9399));
  NANDX1 G30876 (.A1(W4022), .A2(I1460), .ZN(W9400));
  NANDX1 G30877 (.A1(W12973), .A2(W9741), .ZN(W22730));
  NANDX1 G30878 (.A1(W6468), .A2(I1634), .ZN(W9401));
  NANDX1 G30879 (.A1(W1927), .A2(W23218), .ZN(W24649));
  NANDX1 G30880 (.A1(W6130), .A2(W1910), .ZN(W10525));
  NANDX1 G30881 (.A1(W6552), .A2(I1632), .ZN(W11396));
  NANDX1 G30882 (.A1(I1656), .A2(I1329), .ZN(W1795));
  NANDX1 G30883 (.A1(W6663), .A2(W17343), .ZN(O2596));
  NANDX1 G30884 (.A1(I1002), .A2(I1003), .ZN(W501));
  NANDX1 G30885 (.A1(W6892), .A2(W10602), .ZN(W22589));
  NANDX1 G30886 (.A1(W22742), .A2(W7464), .ZN(W24715));
  NANDX1 G30887 (.A1(I1021), .A2(I1330), .ZN(O3170));
  NANDX1 G30888 (.A1(W5510), .A2(W6912), .ZN(O284));
  NANDX1 G30889 (.A1(I316), .A2(I31), .ZN(W1901));
  NANDX1 G30890 (.A1(I876), .A2(I877), .ZN(W438));
  NANDX1 G30891 (.A1(I878), .A2(I879), .ZN(W439));
  NANDX1 G30892 (.A1(W630), .A2(I1969), .ZN(W1896));
  NANDX1 G30893 (.A1(W2075), .A2(W10454), .ZN(W22580));
  NANDX1 G30894 (.A1(W1710), .A2(W7775), .ZN(W22581));
  NANDX1 G30895 (.A1(W14846), .A2(W857), .ZN(W22582));
  NANDX1 G30896 (.A1(W368), .A2(W6675), .ZN(W10497));
  NANDX1 G30897 (.A1(W962), .A2(I609), .ZN(W1894));
  NANDX1 G30898 (.A1(I886), .A2(I887), .ZN(W443));
  NANDX1 G30899 (.A1(W5616), .A2(W2206), .ZN(W24708));
  NANDX1 G30900 (.A1(I738), .A2(I1271), .ZN(W1892));
  NANDX1 G30901 (.A1(W18218), .A2(W18783), .ZN(O2550));
  NANDX1 G30902 (.A1(W7896), .A2(I1636), .ZN(W22590));
  NANDX1 G30903 (.A1(W22515), .A2(W14949), .ZN(O2553));
  NANDX1 G30904 (.A1(I892), .A2(I893), .ZN(W446));
  NANDX1 G30905 (.A1(W487), .A2(W8930), .ZN(W11451));
  NANDX1 G30906 (.A1(W4979), .A2(W8355), .ZN(W10499));
  NANDX1 G30907 (.A1(W19099), .A2(W23640), .ZN(W24705));
  NANDX1 G30908 (.A1(I1786), .A2(W1049), .ZN(W1887));
  NANDX1 G30909 (.A1(W12521), .A2(I375), .ZN(W22595));
  NANDX1 G30910 (.A1(W881), .A2(I175), .ZN(W1886));
  NANDX1 G30911 (.A1(W9952), .A2(W6937), .ZN(W11449));
  NANDX1 G30912 (.A1(W7927), .A2(W2935), .ZN(W10500));
  NANDX1 G30913 (.A1(I691), .A2(W10003), .ZN(W22599));
  NANDX1 G30914 (.A1(I900), .A2(I901), .ZN(W450));
  NANDX1 G30915 (.A1(I1380), .A2(I1598), .ZN(W1884));
  NANDX1 G30916 (.A1(W2751), .A2(W11018), .ZN(W24722));
  NANDX1 G30917 (.A1(W8376), .A2(W21857), .ZN(W22545));
  NANDX1 G30918 (.A1(I1262), .A2(I1524), .ZN(W1926));
  NANDX1 G30919 (.A1(W1140), .A2(I994), .ZN(W1925));
  NANDX1 G30920 (.A1(W1380), .A2(I161), .ZN(W1922));
  NANDX1 G30921 (.A1(W1031), .A2(W602), .ZN(W1921));
  NANDX1 G30922 (.A1(I1141), .A2(W940), .ZN(W1920));
  NANDX1 G30923 (.A1(W13271), .A2(W21354), .ZN(O2545));
  NANDX1 G30924 (.A1(W942), .A2(W1065), .ZN(W1917));
  NANDX1 G30925 (.A1(W13866), .A2(W3843), .ZN(O2546));
  NANDX1 G30926 (.A1(W20112), .A2(W13958), .ZN(W24725));
  NANDX1 G30927 (.A1(W9149), .A2(W4282), .ZN(W11462));
  NANDX1 G30928 (.A1(W17092), .A2(W11918), .ZN(W22555));
  NANDX1 G30929 (.A1(W6413), .A2(W8331), .ZN(O512));
  NANDX1 G30930 (.A1(W15351), .A2(I1220), .ZN(O2548));
  NANDX1 G30931 (.A1(W21349), .A2(W4633), .ZN(W24723));
  NANDX1 G30932 (.A1(W10194), .A2(W10345), .ZN(W11448));
  NANDX1 G30933 (.A1(W810), .A2(W1321), .ZN(W1911));
  NANDX1 G30934 (.A1(I830), .A2(W1205), .ZN(W1910));
  NANDX1 G30935 (.A1(W16790), .A2(W1085), .ZN(W22558));
  NANDX1 G30936 (.A1(W171), .A2(W152), .ZN(W1909));
  NANDX1 G30937 (.A1(I872), .A2(I873), .ZN(W436));
  NANDX1 G30938 (.A1(I1033), .A2(W3833), .ZN(O349));
  NANDX1 G30939 (.A1(W98), .A2(W614), .ZN(W1908));
  NANDX1 G30940 (.A1(W2921), .A2(W3548), .ZN(W9345));
  NANDX1 G30941 (.A1(W8402), .A2(W22074), .ZN(W24719));
  NANDX1 G30942 (.A1(W17740), .A2(W11527), .ZN(W22562));
  NANDX1 G30943 (.A1(I212), .A2(W6678), .ZN(W11456));
  NANDX1 G30944 (.A1(W1615), .A2(I154), .ZN(W1904));
  NANDX1 G30945 (.A1(W6059), .A2(W4952), .ZN(W24716));
  NANDX1 G30946 (.A1(W12828), .A2(W6279), .ZN(O2549));
  NANDX1 G30947 (.A1(W7838), .A2(I1264), .ZN(W9365));
  NANDX1 G30948 (.A1(W22868), .A2(W18800), .ZN(W24687));
  NANDX1 G30949 (.A1(W19563), .A2(W4393), .ZN(W22615));
  NANDX1 G30950 (.A1(I437), .A2(W1687), .ZN(W1863));
  NANDX1 G30951 (.A1(W9788), .A2(W2749), .ZN(W11438));
  NANDX1 G30952 (.A1(I932), .A2(I933), .ZN(W466));
  NANDX1 G30953 (.A1(I1585), .A2(W8348), .ZN(W9989));
  NANDX1 G30954 (.A1(W3667), .A2(W18809), .ZN(O2558));
  NANDX1 G30955 (.A1(W22448), .A2(W9335), .ZN(O3164));
  NANDX1 G30956 (.A1(W1666), .A2(W1246), .ZN(W1861));
  NANDX1 G30957 (.A1(W13320), .A2(W11060), .ZN(W22619));
  NANDX1 G30958 (.A1(I938), .A2(I939), .ZN(W469));
  NANDX1 G30959 (.A1(W20322), .A2(W6256), .ZN(W22620));
  NANDX1 G30960 (.A1(W2568), .A2(I1261), .ZN(W24685));
  NANDX1 G30961 (.A1(W3376), .A2(W22757), .ZN(O3163));
  NANDX1 G30962 (.A1(I940), .A2(I941), .ZN(W470));
  NANDX1 G30963 (.A1(W15234), .A2(W9092), .ZN(W22614));
  NANDX1 G30964 (.A1(I944), .A2(I945), .ZN(W472));
  NANDX1 G30965 (.A1(I207), .A2(I902), .ZN(W1858));
  NANDX1 G30966 (.A1(I1165), .A2(W4203), .ZN(W9366));
  NANDX1 G30967 (.A1(W11182), .A2(W5273), .ZN(W11436));
  NANDX1 G30968 (.A1(I1622), .A2(I1570), .ZN(W1855));
  NANDX1 G30969 (.A1(I946), .A2(I947), .ZN(W473));
  NANDX1 G30970 (.A1(I1933), .A2(W1472), .ZN(W1854));
  NANDX1 G30971 (.A1(W8157), .A2(I622), .ZN(W9367));
  NANDX1 G30972 (.A1(I1274), .A2(I1449), .ZN(W1852));
  NANDX1 G30973 (.A1(I1074), .A2(W15270), .ZN(W22633));
  NANDX1 G30974 (.A1(I952), .A2(I953), .ZN(W476));
  NANDX1 G30975 (.A1(W4118), .A2(W801), .ZN(W11429));
  NANDX1 G30976 (.A1(W410), .A2(W181), .ZN(W1846));
  NANDX1 G30977 (.A1(W5526), .A2(W6059), .ZN(W10512));
  NANDX1 G30978 (.A1(W1956), .A2(W8943), .ZN(O2555));
  NANDX1 G30979 (.A1(W2511), .A2(W9554), .ZN(W11446));
  NANDX1 G30980 (.A1(I902), .A2(I903), .ZN(W451));
  NANDX1 G30981 (.A1(W853), .A2(W20798), .ZN(W22602));
  NANDX1 G30982 (.A1(I904), .A2(I905), .ZN(W452));
  NANDX1 G30983 (.A1(I906), .A2(I907), .ZN(W453));
  NANDX1 G30984 (.A1(W1254), .A2(W1277), .ZN(W1882));
  NANDX1 G30985 (.A1(W996), .A2(W1189), .ZN(W1881));
  NANDX1 G30986 (.A1(W7831), .A2(W1539), .ZN(W9992));
  NANDX1 G30987 (.A1(W1368), .A2(I396), .ZN(W1877));
  NANDX1 G30988 (.A1(W3034), .A2(W12228), .ZN(O2554));
  NANDX1 G30989 (.A1(W3966), .A2(W17603), .ZN(W24699));
  NANDX1 G30990 (.A1(W6889), .A2(W5), .ZN(W9356));
  NANDX1 G30991 (.A1(I918), .A2(I919), .ZN(W459));
  NANDX1 G30992 (.A1(I920), .A2(I921), .ZN(W460));
  NANDX1 G30993 (.A1(W5952), .A2(W19533), .ZN(W23228));
  NANDX1 G30994 (.A1(I1639), .A2(I1698), .ZN(W1873));
  NANDX1 G30995 (.A1(I926), .A2(I927), .ZN(W463));
  NANDX1 G30996 (.A1(W4494), .A2(W2135), .ZN(W10504));
  NANDX1 G30997 (.A1(W9997), .A2(W19110), .ZN(W24691));
  NANDX1 G30998 (.A1(W3451), .A2(W21681), .ZN(W22608));
  NANDX1 G30999 (.A1(W9079), .A2(W5384), .ZN(W9358));
  NANDX1 G31000 (.A1(W16873), .A2(W10979), .ZN(W22609));
  NANDX1 G31001 (.A1(W1705), .A2(I120), .ZN(W1869));
  NANDX1 G31002 (.A1(W598), .A2(W1698), .ZN(W10506));
  NANDX1 G31003 (.A1(W2512), .A2(W9781), .ZN(O401));
  NANDX1 G31004 (.A1(W1696), .A2(W553), .ZN(W1866));
  NANDX1 G31005 (.A1(W402), .A2(W5002), .ZN(W9360));
  NANDX1 G31006 (.A1(W14350), .A2(W61), .ZN(W22613));
  NANDX1 G31007 (.A1(W11563), .A2(W14086), .ZN(O3165));
  NANDX1 G31008 (.A1(W5476), .A2(W4068), .ZN(W9872));
  NANDX1 G31009 (.A1(W7401), .A2(W2694), .ZN(O446));
  NANDX1 G31010 (.A1(W5815), .A2(W8612), .ZN(W9756));
  NANDX1 G31011 (.A1(I1642), .A2(W3624), .ZN(W10873));
  NANDX1 G31012 (.A1(W242), .A2(I704), .ZN(W1066));
  NANDX1 G31013 (.A1(I464), .A2(I1935), .ZN(W1065));
  NANDX1 G31014 (.A1(W1200), .A2(W16), .ZN(W9758));
  NANDX1 G31015 (.A1(I1104), .A2(W1145), .ZN(O445));
  NANDX1 G31016 (.A1(W6966), .A2(W4665), .ZN(W10694));
  NANDX1 G31017 (.A1(W2718), .A2(W23914), .ZN(W24240));
  NANDX1 G31018 (.A1(W18760), .A2(W7454), .ZN(W23790));
  NANDX1 G31019 (.A1(W755), .A2(I104), .ZN(W1063));
  NANDX1 G31020 (.A1(W4801), .A2(W9343), .ZN(O2881));
  NANDX1 G31021 (.A1(W4804), .A2(W2925), .ZN(W10695));
  NANDX1 G31022 (.A1(W411), .A2(W991), .ZN(W10870));
  NANDX1 G31023 (.A1(W2267), .A2(W20705), .ZN(W23793));
  NANDX1 G31024 (.A1(W239), .A2(I1811), .ZN(W1068));
  NANDX1 G31025 (.A1(I1716), .A2(W16741), .ZN(W23796));
  NANDX1 G31026 (.A1(W18550), .A2(W3072), .ZN(O3011));
  NANDX1 G31027 (.A1(W17736), .A2(I1743), .ZN(O2883));
  NANDX1 G31028 (.A1(W2479), .A2(W16847), .ZN(W23798));
  NANDX1 G31029 (.A1(I1546), .A2(I79), .ZN(W1059));
  NANDX1 G31030 (.A1(I1393), .A2(W1195), .ZN(W9760));
  NANDX1 G31031 (.A1(I1552), .A2(I1553), .ZN(W776));
  NANDX1 G31032 (.A1(W10152), .A2(W21055), .ZN(O3010));
  NANDX1 G31033 (.A1(W10375), .A2(W8006), .ZN(W10864));
  NANDX1 G31034 (.A1(W11007), .A2(W18566), .ZN(W23805));
  NANDX1 G31035 (.A1(W6397), .A2(W19039), .ZN(O2885));
  NANDX1 G31036 (.A1(I1911), .A2(W5816), .ZN(W9871));
  NANDX1 G31037 (.A1(W9645), .A2(W2863), .ZN(W10863));
  NANDX1 G31038 (.A1(I1343), .A2(I1432), .ZN(W1056));
  NANDX1 G31039 (.A1(I1534), .A2(I1535), .ZN(W767));
  NANDX1 G31040 (.A1(I1534), .A2(W217), .ZN(W1085));
  NANDX1 G31041 (.A1(W2391), .A2(W7649), .ZN(W9748));
  NANDX1 G31042 (.A1(W6732), .A2(W1776), .ZN(W10889));
  NANDX1 G31043 (.A1(W5775), .A2(W8447), .ZN(W9875));
  NANDX1 G31044 (.A1(W12446), .A2(W908), .ZN(O3019));
  NANDX1 G31045 (.A1(I1530), .A2(I1531), .ZN(W765));
  NANDX1 G31046 (.A1(W13496), .A2(W10054), .ZN(O2872));
  NANDX1 G31047 (.A1(I1098), .A2(W14677), .ZN(W23768));
  NANDX1 G31048 (.A1(W1710), .A2(W5937), .ZN(O449));
  NANDX1 G31049 (.A1(W2056), .A2(W425), .ZN(W10886));
  NANDX1 G31050 (.A1(W2605), .A2(W169), .ZN(O448));
  NANDX1 G31051 (.A1(W11815), .A2(W10297), .ZN(O2873));
  NANDX1 G31052 (.A1(W1407), .A2(W2260), .ZN(W10692));
  NANDX1 G31053 (.A1(I896), .A2(W5860), .ZN(W9750));
  NANDX1 G31054 (.A1(W6432), .A2(W2479), .ZN(W10884));
  NANDX1 G31055 (.A1(W2133), .A2(W23793), .ZN(O3009));
  NANDX1 G31056 (.A1(W2127), .A2(W9394), .ZN(W23775));
  NANDX1 G31057 (.A1(W11225), .A2(W14360), .ZN(W24251));
  NANDX1 G31058 (.A1(I555), .A2(W545), .ZN(W1075));
  NANDX1 G31059 (.A1(W10598), .A2(W2110), .ZN(W23778));
  NANDX1 G31060 (.A1(W16666), .A2(W2752), .ZN(O2877));
  NANDX1 G31061 (.A1(W18589), .A2(W5101), .ZN(W24248));
  NANDX1 G31062 (.A1(W6384), .A2(I1324), .ZN(O3016));
  NANDX1 G31063 (.A1(I1744), .A2(W8012), .ZN(O322));
  NANDX1 G31064 (.A1(W8044), .A2(W19498), .ZN(O3015));
  NANDX1 G31065 (.A1(W1671), .A2(W897), .ZN(W24243));
  NANDX1 G31066 (.A1(W3462), .A2(W9578), .ZN(W10880));
  NANDX1 G31067 (.A1(W4807), .A2(W9665), .ZN(W10878));
  NANDX1 G31068 (.A1(I1544), .A2(I1545), .ZN(W772));
  NANDX1 G31069 (.A1(W11695), .A2(W23179), .ZN(W23785));
  NANDX1 G31070 (.A1(W5512), .A2(W12704), .ZN(O2903));
  NANDX1 G31071 (.A1(I720), .A2(W5594), .ZN(W9859));
  NANDX1 G31072 (.A1(W13921), .A2(W15181), .ZN(W23841));
  NANDX1 G31073 (.A1(W97), .A2(W7656), .ZN(O442));
  NANDX1 G31074 (.A1(I925), .A2(W421), .ZN(W1038));
  NANDX1 G31075 (.A1(W21688), .A2(I1496), .ZN(O2899));
  NANDX1 G31076 (.A1(W4283), .A2(W16215), .ZN(W23847));
  NANDX1 G31077 (.A1(W1766), .A2(W3318), .ZN(W10851));
  NANDX1 G31078 (.A1(W12397), .A2(W23687), .ZN(W23850));
  NANDX1 G31079 (.A1(W1464), .A2(W18420), .ZN(W23852));
  NANDX1 G31080 (.A1(W5738), .A2(W52), .ZN(W9857));
  NANDX1 G31081 (.A1(W2055), .A2(W1863), .ZN(W10850));
  NANDX1 G31082 (.A1(I1782), .A2(I1354), .ZN(W1034));
  NANDX1 G31083 (.A1(W18049), .A2(W11783), .ZN(O2902));
  NANDX1 G31084 (.A1(W8566), .A2(W4658), .ZN(W23856));
  NANDX1 G31085 (.A1(W15486), .A2(W7242), .ZN(W23857));
  NANDX1 G31086 (.A1(I495), .A2(W186), .ZN(W1041));
  NANDX1 G31087 (.A1(I1584), .A2(I1585), .ZN(W792));
  NANDX1 G31088 (.A1(W749), .A2(I429), .ZN(W1031));
  NANDX1 G31089 (.A1(W6604), .A2(W5037), .ZN(W24218));
  NANDX1 G31090 (.A1(W8484), .A2(W6195), .ZN(W9768));
  NANDX1 G31091 (.A1(W274), .A2(W6995), .ZN(W10704));
  NANDX1 G31092 (.A1(W18830), .A2(W16824), .ZN(W24215));
  NANDX1 G31093 (.A1(W13759), .A2(W19641), .ZN(O3003));
  NANDX1 G31094 (.A1(W418), .A2(W214), .ZN(W1029));
  NANDX1 G31095 (.A1(W10449), .A2(W870), .ZN(O2907));
  NANDX1 G31096 (.A1(I1588), .A2(I1589), .ZN(W794));
  NANDX1 G31097 (.A1(W3665), .A2(I370), .ZN(W9771));
  NANDX1 G31098 (.A1(W10298), .A2(W5363), .ZN(W10847));
  NANDX1 G31099 (.A1(I1758), .A2(I534), .ZN(W1027));
  NANDX1 G31100 (.A1(I1590), .A2(I1591), .ZN(W795));
  NANDX1 G31101 (.A1(I1562), .A2(I1563), .ZN(W781));
  NANDX1 G31102 (.A1(W6274), .A2(W13620), .ZN(W23813));
  NANDX1 G31103 (.A1(W14279), .A2(W15284), .ZN(W23816));
  NANDX1 G31104 (.A1(I911), .A2(W17752), .ZN(W23819));
  NANDX1 G31105 (.A1(W8878), .A2(W8401), .ZN(W10862));
  NANDX1 G31106 (.A1(I1146), .A2(I1459), .ZN(W1052));
  NANDX1 G31107 (.A1(I180), .A2(I574), .ZN(W1050));
  NANDX1 G31108 (.A1(W20694), .A2(W20305), .ZN(W24228));
  NANDX1 G31109 (.A1(W950), .A2(W8854), .ZN(W10699));
  NANDX1 G31110 (.A1(W245), .A2(W200), .ZN(W1049));
  NANDX1 G31111 (.A1(W13315), .A2(W4923), .ZN(W23823));
  NANDX1 G31112 (.A1(I1560), .A2(I1561), .ZN(W780));
  NANDX1 G31113 (.A1(W16139), .A2(W14746), .ZN(W23824));
  NANDX1 G31114 (.A1(I633), .A2(W51), .ZN(W1048));
  NANDX1 G31115 (.A1(W13156), .A2(W21431), .ZN(O2891));
  NANDX1 G31116 (.A1(W11449), .A2(W18994), .ZN(W23827));
  NANDX1 G31117 (.A1(W20541), .A2(W65), .ZN(O2870));
  NANDX1 G31118 (.A1(I165), .A2(I736), .ZN(W1047));
  NANDX1 G31119 (.A1(W3551), .A2(I1804), .ZN(W10859));
  NANDX1 G31120 (.A1(W23310), .A2(W9055), .ZN(O2892));
  NANDX1 G31121 (.A1(W21432), .A2(W3531), .ZN(W23829));
  NANDX1 G31122 (.A1(I1564), .A2(I1565), .ZN(W782));
  NANDX1 G31123 (.A1(W9985), .A2(W3146), .ZN(W24225));
  NANDX1 G31124 (.A1(W9683), .A2(W9610), .ZN(W10857));
  NANDX1 G31125 (.A1(W14846), .A2(W9142), .ZN(W23831));
  NANDX1 G31126 (.A1(W71), .A2(I1374), .ZN(W1044));
  NANDX1 G31127 (.A1(I1570), .A2(I1571), .ZN(W785));
  NANDX1 G31128 (.A1(W13436), .A2(W13543), .ZN(W24223));
  NANDX1 G31129 (.A1(W6921), .A2(W15011), .ZN(O2894));
  NANDX1 G31130 (.A1(W6423), .A2(W14118), .ZN(O2895));
  NANDX1 G31131 (.A1(W13775), .A2(W22627), .ZN(O3006));
  NANDX1 G31132 (.A1(W7722), .A2(W8363), .ZN(O3032));
  NANDX1 G31133 (.A1(I384), .A2(I477), .ZN(W1156));
  NANDX1 G31134 (.A1(I1496), .A2(I1497), .ZN(W748));
  NANDX1 G31135 (.A1(W3081), .A2(I1923), .ZN(W23680));
  NANDX1 G31136 (.A1(W2423), .A2(W13317), .ZN(O2849));
  NANDX1 G31137 (.A1(W20856), .A2(W22666), .ZN(W24286));
  NANDX1 G31138 (.A1(W1073), .A2(W6159), .ZN(W10683));
  NANDX1 G31139 (.A1(I376), .A2(W675), .ZN(W1154));
  NANDX1 G31140 (.A1(I1500), .A2(I1501), .ZN(W750));
  NANDX1 G31141 (.A1(I598), .A2(W83), .ZN(W1153));
  NANDX1 G31142 (.A1(I1502), .A2(I1503), .ZN(W751));
  NANDX1 G31143 (.A1(W169), .A2(I1746), .ZN(W1149));
  NANDX1 G31144 (.A1(W17875), .A2(W20701), .ZN(W23688));
  NANDX1 G31145 (.A1(I1467), .A2(W12688), .ZN(O2851));
  NANDX1 G31146 (.A1(W1071), .A2(W670), .ZN(W1148));
  NANDX1 G31147 (.A1(W445), .A2(W3667), .ZN(O454));
  NANDX1 G31148 (.A1(I1488), .A2(I1489), .ZN(W744));
  NANDX1 G31149 (.A1(W8082), .A2(W20716), .ZN(W23692));
  NANDX1 G31150 (.A1(W989), .A2(I998), .ZN(W1146));
  NANDX1 G31151 (.A1(W749), .A2(W253), .ZN(W1145));
  NANDX1 G31152 (.A1(I1799), .A2(W7855), .ZN(W23694));
  NANDX1 G31153 (.A1(W10233), .A2(I921), .ZN(W10920));
  NANDX1 G31154 (.A1(W8422), .A2(W19760), .ZN(W23695));
  NANDX1 G31155 (.A1(W17560), .A2(W51), .ZN(W23698));
  NANDX1 G31156 (.A1(W259), .A2(W4500), .ZN(W10684));
  NANDX1 G31157 (.A1(W18179), .A2(W22976), .ZN(W23702));
  NANDX1 G31158 (.A1(I364), .A2(W650), .ZN(W1140));
  NANDX1 G31159 (.A1(I1504), .A2(I1505), .ZN(W752));
  NANDX1 G31160 (.A1(W16981), .A2(W1556), .ZN(W23704));
  NANDX1 G31161 (.A1(W5894), .A2(W2871), .ZN(W10919));
  NANDX1 G31162 (.A1(I442), .A2(I1593), .ZN(W1139));
  NANDX1 G31163 (.A1(W13765), .A2(W265), .ZN(W23668));
  NANDX1 G31164 (.A1(W4047), .A2(W2629), .ZN(W9727));
  NANDX1 G31165 (.A1(W623), .A2(I848), .ZN(W10934));
  NANDX1 G31166 (.A1(W734), .A2(W207), .ZN(W1168));
  NANDX1 G31167 (.A1(W7406), .A2(W10152), .ZN(O2842));
  NANDX1 G31168 (.A1(W11406), .A2(W23573), .ZN(O2843));
  NANDX1 G31169 (.A1(W4526), .A2(W16627), .ZN(W23662));
  NANDX1 G31170 (.A1(W3385), .A2(W21428), .ZN(W23663));
  NANDX1 G31171 (.A1(W7778), .A2(W1209), .ZN(W10933));
  NANDX1 G31172 (.A1(I122), .A2(W8449), .ZN(W24298));
  NANDX1 G31173 (.A1(W2170), .A2(W1844), .ZN(W10931));
  NANDX1 G31174 (.A1(W652), .A2(I1426), .ZN(W1165));
  NANDX1 G31175 (.A1(W6687), .A2(W9464), .ZN(W9884));
  NANDX1 G31176 (.A1(W16108), .A2(W9372), .ZN(O2844));
  NANDX1 G31177 (.A1(W2989), .A2(I190), .ZN(W9728));
  NANDX1 G31178 (.A1(W17387), .A2(W6120), .ZN(O2845));
  NANDX1 G31179 (.A1(I1506), .A2(I1507), .ZN(W753));
  NANDX1 G31180 (.A1(W931), .A2(I335), .ZN(W1162));
  NANDX1 G31181 (.A1(W9369), .A2(W14646), .ZN(W24296));
  NANDX1 G31182 (.A1(I1972), .A2(W92), .ZN(W1160));
  NANDX1 G31183 (.A1(W18844), .A2(W11064), .ZN(W23670));
  NANDX1 G31184 (.A1(W12633), .A2(W4512), .ZN(W23671));
  NANDX1 G31185 (.A1(I1480), .A2(I678), .ZN(W1159));
  NANDX1 G31186 (.A1(W7345), .A2(W9456), .ZN(W9883));
  NANDX1 G31187 (.A1(W7841), .A2(W6433), .ZN(W23674));
  NANDX1 G31188 (.A1(W7896), .A2(I710), .ZN(W10679));
  NANDX1 G31189 (.A1(I1482), .A2(I1483), .ZN(W741));
  NANDX1 G31190 (.A1(W754), .A2(W57), .ZN(W1158));
  NANDX1 G31191 (.A1(W2923), .A2(I44), .ZN(W23678));
  NANDX1 G31192 (.A1(W6234), .A2(W64), .ZN(O422));
  NANDX1 G31193 (.A1(W5972), .A2(W6206), .ZN(W10681));
  NANDX1 G31194 (.A1(W8164), .A2(W7778), .ZN(W9876));
  NANDX1 G31195 (.A1(W10904), .A2(W8402), .ZN(W10908));
  NANDX1 G31196 (.A1(W8496), .A2(W4937), .ZN(W9877));
  NANDX1 G31197 (.A1(I1612), .A2(W891), .ZN(W1104));
  NANDX1 G31198 (.A1(W6290), .A2(I1352), .ZN(W23741));
  NANDX1 G31199 (.A1(W4586), .A2(W8487), .ZN(W24260));
  NANDX1 G31200 (.A1(W10315), .A2(W10103), .ZN(W10907));
  NANDX1 G31201 (.A1(I210), .A2(W775), .ZN(W1102));
  NANDX1 G31202 (.A1(I1522), .A2(I1523), .ZN(W761));
  NANDX1 G31203 (.A1(W8992), .A2(W5276), .ZN(W10905));
  NANDX1 G31204 (.A1(W5672), .A2(W11016), .ZN(W24259));
  NANDX1 G31205 (.A1(W6678), .A2(W6042), .ZN(W10902));
  NANDX1 G31206 (.A1(W1191), .A2(W19312), .ZN(O2865));
  NANDX1 G31207 (.A1(W5355), .A2(W7575), .ZN(W10901));
  NANDX1 G31208 (.A1(W18119), .A2(W11719), .ZN(O2866));
  NANDX1 G31209 (.A1(W8837), .A2(W4252), .ZN(W10900));
  NANDX1 G31210 (.A1(W5180), .A2(W3725), .ZN(W23739));
  NANDX1 G31211 (.A1(W276), .A2(W30), .ZN(W1093));
  NANDX1 G31212 (.A1(W19103), .A2(W22482), .ZN(W23750));
  NANDX1 G31213 (.A1(W2229), .A2(W7471), .ZN(W10898));
  NANDX1 G31214 (.A1(W11433), .A2(W5280), .ZN(W23752));
  NANDX1 G31215 (.A1(I387), .A2(I831), .ZN(W10689));
  NANDX1 G31216 (.A1(W9591), .A2(W1671), .ZN(W10691));
  NANDX1 G31217 (.A1(I1528), .A2(I1529), .ZN(W764));
  NANDX1 G31218 (.A1(W20400), .A2(W993), .ZN(W23755));
  NANDX1 G31219 (.A1(W1737), .A2(W766), .ZN(W10895));
  NANDX1 G31220 (.A1(W22238), .A2(W15983), .ZN(W23758));
  NANDX1 G31221 (.A1(I55), .A2(W729), .ZN(W1089));
  NANDX1 G31222 (.A1(W935), .A2(W3739), .ZN(W10894));
  NANDX1 G31223 (.A1(W792), .A2(W2469), .ZN(W9747));
  NANDX1 G31224 (.A1(W20895), .A2(W20281), .ZN(W23760));
  NANDX1 G31225 (.A1(W231), .A2(I1161), .ZN(W1129));
  NANDX1 G31226 (.A1(W5776), .A2(W8619), .ZN(W10917));
  NANDX1 G31227 (.A1(W2020), .A2(W8390), .ZN(W10685));
  NANDX1 G31228 (.A1(W21543), .A2(W22496), .ZN(W23709));
  NANDX1 G31229 (.A1(W13960), .A2(W18824), .ZN(W23710));
  NANDX1 G31230 (.A1(W8368), .A2(I999), .ZN(W10686));
  NANDX1 G31231 (.A1(I628), .A2(W16635), .ZN(W24270));
  NANDX1 G31232 (.A1(W771), .A2(I562), .ZN(W1133));
  NANDX1 G31233 (.A1(W774), .A2(I1287), .ZN(O8));
  NANDX1 G31234 (.A1(I673), .A2(W1061), .ZN(W1130));
  NANDX1 G31235 (.A1(I1512), .A2(I1513), .ZN(W756));
  NANDX1 G31236 (.A1(W9157), .A2(W9355), .ZN(W9737));
  NANDX1 G31237 (.A1(W752), .A2(W6494), .ZN(W9738));
  NANDX1 G31238 (.A1(W8497), .A2(W6509), .ZN(W10687));
  NANDX1 G31239 (.A1(W10469), .A2(W5882), .ZN(O424));
  NANDX1 G31240 (.A1(W22676), .A2(I765), .ZN(O2858));
  NANDX1 G31241 (.A1(W11676), .A2(W4752), .ZN(O2909));
  NANDX1 G31242 (.A1(W1731), .A2(W23021), .ZN(W24267));
  NANDX1 G31243 (.A1(I943), .A2(W506), .ZN(W1125));
  NANDX1 G31244 (.A1(W2407), .A2(W19265), .ZN(W23722));
  NANDX1 G31245 (.A1(W19547), .A2(W15338), .ZN(W24265));
  NANDX1 G31246 (.A1(W6269), .A2(W3816), .ZN(W9882));
  NANDX1 G31247 (.A1(I1438), .A2(W346), .ZN(W1121));
  NANDX1 G31248 (.A1(W374), .A2(I1959), .ZN(W1120));
  NANDX1 G31249 (.A1(I1968), .A2(W47), .ZN(W1119));
  NANDX1 G31250 (.A1(I664), .A2(I456), .ZN(W1114));
  NANDX1 G31251 (.A1(W9267), .A2(W1851), .ZN(W9743));
  NANDX1 G31252 (.A1(I1518), .A2(I1519), .ZN(W759));
  NANDX1 G31253 (.A1(W55), .A2(I1642), .ZN(W1108));
  NANDX1 G31254 (.A1(W10299), .A2(I285), .ZN(W10910));
  NANDX1 G31255 (.A1(I414), .A2(I882), .ZN(W1107));
  NANDX1 G31256 (.A1(I1814), .A2(I1815), .ZN(W907));
  NANDX1 G31257 (.A1(W805), .A2(W10370), .ZN(O2954));
  NANDX1 G31258 (.A1(W1810), .A2(I121), .ZN(W10778));
  NANDX1 G31259 (.A1(I200), .A2(W1874), .ZN(W10777));
  NANDX1 G31260 (.A1(I1824), .A2(I1825), .ZN(W912));
  NANDX1 G31261 (.A1(W5816), .A2(W15618), .ZN(W24031));
  NANDX1 G31262 (.A1(W19501), .A2(W9216), .ZN(W24032));
  NANDX1 G31263 (.A1(I1694), .A2(I1695), .ZN(W847));
  NANDX1 G31264 (.A1(I1818), .A2(I1819), .ZN(W909));
  NANDX1 G31265 (.A1(W6632), .A2(W3251), .ZN(W24139));
  NANDX1 G31266 (.A1(W1661), .A2(W3056), .ZN(W10773));
  NANDX1 G31267 (.A1(W12170), .A2(W10597), .ZN(O2956));
  NANDX1 G31268 (.A1(W14686), .A2(W5511), .ZN(O2980));
  NANDX1 G31269 (.A1(W7004), .A2(W5450), .ZN(W24039));
  NANDX1 G31270 (.A1(W9600), .A2(W1502), .ZN(O432));
  NANDX1 G31271 (.A1(W22810), .A2(W21644), .ZN(W24041));
  NANDX1 G31272 (.A1(W20070), .A2(I48), .ZN(W24028));
  NANDX1 G31273 (.A1(I1696), .A2(I1697), .ZN(W848));
  NANDX1 G31274 (.A1(I1812), .A2(I1813), .ZN(W906));
  NANDX1 G31275 (.A1(I1810), .A2(I1811), .ZN(W905));
  NANDX1 G31276 (.A1(W10621), .A2(W15998), .ZN(O2958));
  NANDX1 G31277 (.A1(W15592), .A2(W19130), .ZN(W24047));
  NANDX1 G31278 (.A1(I1808), .A2(I1809), .ZN(W904));
  NANDX1 G31279 (.A1(I1806), .A2(I1807), .ZN(W903));
  NANDX1 G31280 (.A1(W16821), .A2(W7820), .ZN(W24137));
  NANDX1 G31281 (.A1(W7438), .A2(W12779), .ZN(W24136));
  NANDX1 G31282 (.A1(W4648), .A2(W17255), .ZN(W24135));
  NANDX1 G31283 (.A1(W1914), .A2(W14388), .ZN(W24134));
  NANDX1 G31284 (.A1(I1802), .A2(I1803), .ZN(W901));
  NANDX1 G31285 (.A1(I1800), .A2(I1801), .ZN(W900));
  NANDX1 G31286 (.A1(I1952), .A2(W1345), .ZN(W10767));
  NANDX1 G31287 (.A1(W4928), .A2(W2999), .ZN(W10787));
  NANDX1 G31288 (.A1(W8324), .A2(W5002), .ZN(W10794));
  NANDX1 G31289 (.A1(I1874), .A2(I1875), .ZN(W937));
  NANDX1 G31290 (.A1(I1680), .A2(I1681), .ZN(W840));
  NANDX1 G31291 (.A1(W8256), .A2(W2630), .ZN(W24159));
  NANDX1 G31292 (.A1(W2696), .A2(W7291), .ZN(W23999));
  NANDX1 G31293 (.A1(W19567), .A2(W9814), .ZN(W24000));
  NANDX1 G31294 (.A1(W4207), .A2(W6965), .ZN(W24001));
  NANDX1 G31295 (.A1(W18040), .A2(W23286), .ZN(O2946));
  NANDX1 G31296 (.A1(W5551), .A2(W13843), .ZN(W24157));
  NANDX1 G31297 (.A1(W4826), .A2(W6857), .ZN(O2947));
  NANDX1 G31298 (.A1(W5798), .A2(W335), .ZN(W10792));
  NANDX1 G31299 (.A1(W22595), .A2(W505), .ZN(W24006));
  NANDX1 G31300 (.A1(W7248), .A2(W7584), .ZN(W9807));
  NANDX1 G31301 (.A1(I1862), .A2(I1863), .ZN(W931));
  NANDX1 G31302 (.A1(W6689), .A2(W4703), .ZN(W10788));
  NANDX1 G31303 (.A1(W9266), .A2(I398), .ZN(W9827));
  NANDX1 G31304 (.A1(W3180), .A2(W640), .ZN(O434));
  NANDX1 G31305 (.A1(W7900), .A2(W9786), .ZN(W24017));
  NANDX1 G31306 (.A1(I1684), .A2(I1685), .ZN(W842));
  NANDX1 G31307 (.A1(W21169), .A2(W19677), .ZN(W24019));
  NANDX1 G31308 (.A1(W16014), .A2(W21425), .ZN(O2951));
  NANDX1 G31309 (.A1(I1840), .A2(I1841), .ZN(W920));
  NANDX1 G31310 (.A1(I1836), .A2(I1837), .ZN(W918));
  NANDX1 G31311 (.A1(I1688), .A2(I1689), .ZN(W844));
  NANDX1 G31312 (.A1(W7086), .A2(I1940), .ZN(W10783));
  NANDX1 G31313 (.A1(W15228), .A2(W2969), .ZN(W24151));
  NANDX1 G31314 (.A1(W6481), .A2(W499), .ZN(W24146));
  NANDX1 G31315 (.A1(W8650), .A2(W18739), .ZN(W24144));
  NANDX1 G31316 (.A1(W1273), .A2(W4594), .ZN(W9829));
  NANDX1 G31317 (.A1(I1840), .A2(W4072), .ZN(W10779));
  NANDX1 G31318 (.A1(I583), .A2(I1652), .ZN(W10752));
  NANDX1 G31319 (.A1(I1758), .A2(I1759), .ZN(W879));
  NANDX1 G31320 (.A1(W858), .A2(W8789), .ZN(W9824));
  NANDX1 G31321 (.A1(I1714), .A2(I1715), .ZN(W857));
  NANDX1 G31322 (.A1(W8807), .A2(W8731), .ZN(W24088));
  NANDX1 G31323 (.A1(I1754), .A2(I1755), .ZN(W877));
  NANDX1 G31324 (.A1(I1718), .A2(I1719), .ZN(W859));
  NANDX1 G31325 (.A1(I104), .A2(W19913), .ZN(W24089));
  NANDX1 G31326 (.A1(W7272), .A2(W22500), .ZN(W24091));
  NANDX1 G31327 (.A1(I1750), .A2(I1751), .ZN(W875));
  NANDX1 G31328 (.A1(W1600), .A2(W7618), .ZN(W9820));
  NANDX1 G31329 (.A1(W20976), .A2(W3081), .ZN(W24093));
  NANDX1 G31330 (.A1(W7837), .A2(W3829), .ZN(W24094));
  NANDX1 G31331 (.A1(W8113), .A2(I1676), .ZN(W10744));
  NANDX1 G31332 (.A1(W22574), .A2(I1267), .ZN(O2969));
  NANDX1 G31333 (.A1(I1748), .A2(I1749), .ZN(W874));
  NANDX1 G31334 (.A1(I1762), .A2(I1763), .ZN(W881));
  NANDX1 G31335 (.A1(W6548), .A2(W9512), .ZN(W10745));
  NANDX1 G31336 (.A1(W6866), .A2(W1082), .ZN(W9821));
  NANDX1 G31337 (.A1(W9925), .A2(W1685), .ZN(W24099));
  NANDX1 G31338 (.A1(W8005), .A2(W5266), .ZN(O2971));
  NANDX1 G31339 (.A1(I1742), .A2(I1743), .ZN(W871));
  NANDX1 G31340 (.A1(W2479), .A2(W262), .ZN(W10749));
  NANDX1 G31341 (.A1(I1726), .A2(I1727), .ZN(W863));
  NANDX1 G31342 (.A1(W18264), .A2(W7104), .ZN(W24109));
  NANDX1 G31343 (.A1(W6957), .A2(W324), .ZN(W10748));
  NANDX1 G31344 (.A1(W2307), .A2(W16665), .ZN(O2975));
  NANDX1 G31345 (.A1(W18046), .A2(W21283), .ZN(O2976));
  NANDX1 G31346 (.A1(I1736), .A2(I1737), .ZN(W868));
  NANDX1 G31347 (.A1(W5626), .A2(W5905), .ZN(W10747));
  NANDX1 G31348 (.A1(W19700), .A2(W2229), .ZN(W24113));
  NANDX1 G31349 (.A1(W10791), .A2(W1591), .ZN(O2965));
  NANDX1 G31350 (.A1(W5923), .A2(W11288), .ZN(O2960));
  NANDX1 G31351 (.A1(I1794), .A2(I1795), .ZN(W897));
  NANDX1 G31352 (.A1(W16468), .A2(W22496), .ZN(W24059));
  NANDX1 G31353 (.A1(W17004), .A2(W3399), .ZN(W24060));
  NANDX1 G31354 (.A1(W8200), .A2(W11738), .ZN(W24131));
  NANDX1 G31355 (.A1(I1700), .A2(I1701), .ZN(W850));
  NANDX1 G31356 (.A1(W10179), .A2(W3963), .ZN(W10765));
  NANDX1 G31357 (.A1(W4220), .A2(W126), .ZN(W24068));
  NANDX1 G31358 (.A1(W3983), .A2(W9622), .ZN(W10764));
  NANDX1 G31359 (.A1(W14498), .A2(W13542), .ZN(O2964));
  NANDX1 G31360 (.A1(W9028), .A2(W2373), .ZN(W10763));
  NANDX1 G31361 (.A1(I382), .A2(W3177), .ZN(W10759));
  NANDX1 G31362 (.A1(W12686), .A2(W6253), .ZN(W24071));
  NANDX1 G31363 (.A1(I1239), .A2(W7628), .ZN(O2978));
  NANDX1 G31364 (.A1(I1782), .A2(I1783), .ZN(W891));
  NANDX1 G31365 (.A1(W14521), .A2(W12728), .ZN(W23996));
  NANDX1 G31366 (.A1(I1271), .A2(W2290), .ZN(W9826));
  NANDX1 G31367 (.A1(W5612), .A2(W6212), .ZN(W10757));
  NANDX1 G31368 (.A1(I1778), .A2(I1779), .ZN(W889));
  NANDX1 G31369 (.A1(I1776), .A2(I1777), .ZN(W888));
  NANDX1 G31370 (.A1(I1774), .A2(I1775), .ZN(W887));
  NANDX1 G31371 (.A1(I1706), .A2(I1707), .ZN(W853));
  NANDX1 G31372 (.A1(W19511), .A2(W14704), .ZN(W24127));
  NANDX1 G31373 (.A1(I1768), .A2(I1769), .ZN(W884));
  NANDX1 G31374 (.A1(I1708), .A2(I1709), .ZN(W854));
  NANDX1 G31375 (.A1(W8087), .A2(W9942), .ZN(W10753));
  NANDX1 G31376 (.A1(I1571), .A2(W3884), .ZN(W10742));
  NANDX1 G31377 (.A1(W2888), .A2(W2335), .ZN(W10743));
  NANDX1 G31378 (.A1(W11332), .A2(W20315), .ZN(O2967));
  NANDX1 G31379 (.A1(W9690), .A2(W14263), .ZN(W24121));
  NANDX1 G31380 (.A1(W9182), .A2(W2010), .ZN(W10721));
  NANDX1 G31381 (.A1(W4109), .A2(W23884), .ZN(O2918));
  NANDX1 G31382 (.A1(W8932), .A2(W2183), .ZN(W9848));
  NANDX1 G31383 (.A1(W6174), .A2(W22984), .ZN(W23906));
  NANDX1 G31384 (.A1(W203), .A2(W6731), .ZN(W23907));
  NANDX1 G31385 (.A1(W776), .A2(I734), .ZN(W1000));
  NANDX1 G31386 (.A1(W384), .A2(W2546), .ZN(W9786));
  NANDX1 G31387 (.A1(W7224), .A2(W514), .ZN(W10718));
  NANDX1 G31388 (.A1(I1608), .A2(I1609), .ZN(W804));
  NANDX1 G31389 (.A1(I1610), .A2(I1611), .ZN(W805));
  NANDX1 G31390 (.A1(W7759), .A2(W5399), .ZN(W10720));
  NANDX1 G31391 (.A1(W6165), .A2(W17622), .ZN(W23918));
  NANDX1 G31392 (.A1(I1992), .A2(I1993), .ZN(W996));
  NANDX1 G31393 (.A1(W10418), .A2(W7489), .ZN(O2921));
  NANDX1 G31394 (.A1(W17827), .A2(W12423), .ZN(W23921));
  NANDX1 G31395 (.A1(W6795), .A2(W6988), .ZN(O2922));
  NANDX1 G31396 (.A1(W1993), .A2(W241), .ZN(W23903));
  NANDX1 G31397 (.A1(I765), .A2(W20873), .ZN(W24202));
  NANDX1 G31398 (.A1(I1986), .A2(I1987), .ZN(W993));
  NANDX1 G31399 (.A1(W6010), .A2(W417), .ZN(W24201));
  NANDX1 G31400 (.A1(I1618), .A2(I1619), .ZN(W809));
  NANDX1 G31401 (.A1(W8291), .A2(W2246), .ZN(W23927));
  NANDX1 G31402 (.A1(I1620), .A2(I1621), .ZN(W810));
  NANDX1 G31403 (.A1(W19325), .A2(W21356), .ZN(W23928));
  NANDX1 G31404 (.A1(W1983), .A2(W9918), .ZN(W10722));
  NANDX1 G31405 (.A1(W8744), .A2(W6766), .ZN(W10723));
  NANDX1 G31406 (.A1(I943), .A2(W6049), .ZN(W9847));
  NANDX1 G31407 (.A1(I1628), .A2(I1629), .ZN(W814));
  NANDX1 G31408 (.A1(W13561), .A2(W18171), .ZN(W23933));
  NANDX1 G31409 (.A1(W5007), .A2(W1622), .ZN(W10725));
  NANDX1 G31410 (.A1(I1974), .A2(I1975), .ZN(W987));
  NANDX1 G31411 (.A1(W20551), .A2(W22202), .ZN(W24209));
  NANDX1 G31412 (.A1(W19473), .A2(W20625), .ZN(W24212));
  NANDX1 G31413 (.A1(W19935), .A2(W7983), .ZN(O3001));
  NANDX1 G31414 (.A1(W8142), .A2(W4217), .ZN(W9851));
  NANDX1 G31415 (.A1(I977), .A2(I1364), .ZN(W10842));
  NANDX1 G31416 (.A1(W886), .A2(W696), .ZN(O441));
  NANDX1 G31417 (.A1(W7028), .A2(W8525), .ZN(W9775));
  NANDX1 G31418 (.A1(W21569), .A2(W10011), .ZN(W23870));
  NANDX1 G31419 (.A1(I973), .A2(I1917), .ZN(W10838));
  NANDX1 G31420 (.A1(W997), .A2(I952), .ZN(W1015));
  NANDX1 G31421 (.A1(W14442), .A2(W14598), .ZN(W23875));
  NANDX1 G31422 (.A1(W17835), .A2(W18032), .ZN(W23878));
  NANDX1 G31423 (.A1(W415), .A2(W428), .ZN(W1014));
  NANDX1 G31424 (.A1(W14205), .A2(W12867), .ZN(W23881));
  NANDX1 G31425 (.A1(I1466), .A2(W390), .ZN(W1013));
  NANDX1 G31426 (.A1(W2981), .A2(W10468), .ZN(W10707));
  NANDX1 G31427 (.A1(W7530), .A2(I459), .ZN(W9844));
  NANDX1 G31428 (.A1(W11505), .A2(W17005), .ZN(W23883));
  NANDX1 G31429 (.A1(W21832), .A2(W11379), .ZN(W23884));
  NANDX1 G31430 (.A1(W6747), .A2(W5370), .ZN(W10710));
  NANDX1 G31431 (.A1(W15640), .A2(W15862), .ZN(W23887));
  NANDX1 G31432 (.A1(W3949), .A2(W9357), .ZN(W9850));
  NANDX1 G31433 (.A1(W7888), .A2(W7829), .ZN(W10831));
  NANDX1 G31434 (.A1(W12072), .A2(W12324), .ZN(W23890));
  NANDX1 G31435 (.A1(I843), .A2(I387), .ZN(W1003));
  NANDX1 G31436 (.A1(W9143), .A2(W7317), .ZN(W23893));
  NANDX1 G31437 (.A1(W15323), .A2(W13845), .ZN(W23894));
  NANDX1 G31438 (.A1(W6696), .A2(W9062), .ZN(W24207));
  NANDX1 G31439 (.A1(W4446), .A2(W17559), .ZN(W23898));
  NANDX1 G31440 (.A1(W487), .A2(I1690), .ZN(W1002));
  NANDX1 G31441 (.A1(W495), .A2(W8869), .ZN(W23902));
  NANDX1 G31442 (.A1(W9401), .A2(W1562), .ZN(W10804));
  NANDX1 G31443 (.A1(I1948), .A2(I1949), .ZN(W974));
  NANDX1 G31444 (.A1(I1662), .A2(I1663), .ZN(W831));
  NANDX1 G31445 (.A1(I1944), .A2(I1945), .ZN(W972));
  NANDX1 G31446 (.A1(I1938), .A2(I1939), .ZN(W969));
  NANDX1 G31447 (.A1(I1936), .A2(I1937), .ZN(W968));
  NANDX1 G31448 (.A1(W14898), .A2(I1647), .ZN(W24169));
  NANDX1 G31449 (.A1(W19019), .A2(I1843), .ZN(W24168));
  NANDX1 G31450 (.A1(I1928), .A2(W10371), .ZN(W10806));
  NANDX1 G31451 (.A1(I1664), .A2(I1665), .ZN(W832));
  NANDX1 G31452 (.A1(W10058), .A2(W16983), .ZN(W24167));
  NANDX1 G31453 (.A1(I1666), .A2(I1667), .ZN(W833));
  NANDX1 G31454 (.A1(W19865), .A2(W3082), .ZN(W23975));
  NANDX1 G31455 (.A1(I1926), .A2(I1927), .ZN(W963));
  NANDX1 G31456 (.A1(I1670), .A2(I1671), .ZN(W835));
  NANDX1 G31457 (.A1(W2776), .A2(W2615), .ZN(W24164));
  NANDX1 G31458 (.A1(W10142), .A2(W20874), .ZN(W24174));
  NANDX1 G31459 (.A1(I1924), .A2(I1925), .ZN(W962));
  NANDX1 G31460 (.A1(W20766), .A2(W23066), .ZN(O2939));
  NANDX1 G31461 (.A1(I1914), .A2(I1915), .ZN(W957));
  NANDX1 G31462 (.A1(W9640), .A2(I1032), .ZN(W10803));
  NANDX1 G31463 (.A1(W20300), .A2(W235), .ZN(W23985));
  NANDX1 G31464 (.A1(W8163), .A2(W141), .ZN(W10801));
  NANDX1 G31465 (.A1(I1888), .A2(I1889), .ZN(W944));
  NANDX1 G31466 (.A1(W15540), .A2(W23823), .ZN(W24161));
  NANDX1 G31467 (.A1(I1676), .A2(I1677), .ZN(W838));
  NANDX1 G31468 (.A1(I1880), .A2(I1881), .ZN(W940));
  NANDX1 G31469 (.A1(W21517), .A2(W3275), .ZN(W23993));
  NANDX1 G31470 (.A1(W5639), .A2(W2923), .ZN(W10736));
  NANDX1 G31471 (.A1(W4662), .A2(W10396), .ZN(O436));
  NANDX1 G31472 (.A1(W7009), .A2(W6179), .ZN(W10795));
  NANDX1 G31473 (.A1(I134), .A2(W14910), .ZN(O2993));
  NANDX1 G31474 (.A1(W7796), .A2(W7309), .ZN(W10818));
  NANDX1 G31475 (.A1(W5240), .A2(W9579), .ZN(W9839));
  NANDX1 G31476 (.A1(W19389), .A2(W1638), .ZN(O2925));
  NANDX1 G31477 (.A1(W3688), .A2(W2882), .ZN(W23939));
  NANDX1 G31478 (.A1(I1964), .A2(I1965), .ZN(W982));
  NANDX1 G31479 (.A1(W9883), .A2(I1087), .ZN(O439));
  NANDX1 G31480 (.A1(W1690), .A2(W2472), .ZN(W23943));
  NANDX1 G31481 (.A1(W5175), .A2(I710), .ZN(W23944));
  NANDX1 G31482 (.A1(W4781), .A2(W1647), .ZN(O2927));
  NANDX1 G31483 (.A1(W20675), .A2(W10534), .ZN(O2928));
  NANDX1 G31484 (.A1(I1648), .A2(I1649), .ZN(W824));
  NANDX1 G31485 (.A1(I1652), .A2(I1653), .ZN(W826));
  NANDX1 G31486 (.A1(W5254), .A2(W14387), .ZN(W23949));
  NANDX1 G31487 (.A1(W20358), .A2(W8119), .ZN(W23950));
  NANDX1 G31488 (.A1(I1454), .A2(W1376), .ZN(W10935));
  NANDX1 G31489 (.A1(I1962), .A2(I1963), .ZN(W981));
  NANDX1 G31490 (.A1(W10692), .A2(W10583), .ZN(W23953));
  NANDX1 G31491 (.A1(W4422), .A2(I1892), .ZN(W23955));
  NANDX1 G31492 (.A1(W21071), .A2(W12498), .ZN(W23956));
  NANDX1 G31493 (.A1(W4539), .A2(I1816), .ZN(O327));
  NANDX1 G31494 (.A1(W6989), .A2(W4730), .ZN(W10729));
  NANDX1 G31495 (.A1(I1570), .A2(W14139), .ZN(O2931));
  NANDX1 G31496 (.A1(I1958), .A2(I1959), .ZN(W979));
  NANDX1 G31497 (.A1(W9835), .A2(W9773), .ZN(W24178));
  NANDX1 G31498 (.A1(W12108), .A2(W3474), .ZN(W23961));
  NANDX1 G31499 (.A1(W9342), .A2(W19709), .ZN(O2992));
  NANDX1 G31500 (.A1(I1954), .A2(I1955), .ZN(W977));
  NANDX1 G31501 (.A1(I1952), .A2(I1953), .ZN(W976));
  NANDX1 G31502 (.A1(W2680), .A2(W2729), .ZN(W9836));
  NANDX1 G31503 (.A1(W6587), .A2(W2557), .ZN(W9924));
  NANDX1 G31504 (.A1(I1912), .A2(W13489), .ZN(W23364));
  NANDX1 G31505 (.A1(W8978), .A2(W3647), .ZN(W11087));
  NANDX1 G31506 (.A1(W9369), .A2(W3765), .ZN(O2752));
  NANDX1 G31507 (.A1(I1354), .A2(I1355), .ZN(W677));
  NANDX1 G31508 (.A1(W6286), .A2(W4266), .ZN(W9617));
  NANDX1 G31509 (.A1(W1074), .A2(W3302), .ZN(W9618));
  NANDX1 G31510 (.A1(I1356), .A2(I1357), .ZN(W678));
  NANDX1 G31511 (.A1(W6397), .A2(W1940), .ZN(W9619));
  NANDX1 G31512 (.A1(W5002), .A2(W4100), .ZN(W9620));
  NANDX1 G31513 (.A1(W11046), .A2(W2379), .ZN(W23367));
  NANDX1 G31514 (.A1(W3046), .A2(W1504), .ZN(W11079));
  NANDX1 G31515 (.A1(W6677), .A2(W22055), .ZN(W23372));
  NANDX1 G31516 (.A1(I161), .A2(W1211), .ZN(W1370));
  NANDX1 G31517 (.A1(W10540), .A2(W15989), .ZN(O3075));
  NANDX1 G31518 (.A1(W8577), .A2(W17859), .ZN(W23374));
  NANDX1 G31519 (.A1(W1289), .A2(I1422), .ZN(W1375));
  NANDX1 G31520 (.A1(W6018), .A2(W3425), .ZN(W9623));
  NANDX1 G31521 (.A1(W1903), .A2(W22340), .ZN(O2753));
  NANDX1 G31522 (.A1(W187), .A2(I1832), .ZN(W1368));
  NANDX1 G31523 (.A1(W11865), .A2(W13106), .ZN(W23382));
  NANDX1 G31524 (.A1(W4764), .A2(I150), .ZN(W11073));
  NANDX1 G31525 (.A1(I435), .A2(I1814), .ZN(W1367));
  NANDX1 G31526 (.A1(W760), .A2(W1234), .ZN(W1366));
  NANDX1 G31527 (.A1(W18179), .A2(W2998), .ZN(O2759));
  NANDX1 G31528 (.A1(I1968), .A2(W19368), .ZN(W24408));
  NANDX1 G31529 (.A1(W4517), .A2(W8633), .ZN(W23389));
  NANDX1 G31530 (.A1(W6203), .A2(W3864), .ZN(O306));
  NANDX1 G31531 (.A1(W5882), .A2(W4418), .ZN(W10625));
  NANDX1 G31532 (.A1(W5191), .A2(I850), .ZN(O2760));
  NANDX1 G31533 (.A1(I1360), .A2(I1361), .ZN(W680));
  NANDX1 G31534 (.A1(W9021), .A2(I315), .ZN(W11096));
  NANDX1 G31535 (.A1(W7949), .A2(W17582), .ZN(W23330));
  NANDX1 G31536 (.A1(W4572), .A2(W8995), .ZN(W11109));
  NANDX1 G31537 (.A1(I1338), .A2(I1339), .ZN(W669));
  NANDX1 G31538 (.A1(I1340), .A2(I1341), .ZN(W670));
  NANDX1 G31539 (.A1(W12826), .A2(W6992), .ZN(W23331));
  NANDX1 G31540 (.A1(W6346), .A2(W6760), .ZN(W9612));
  NANDX1 G31541 (.A1(W12655), .A2(W3594), .ZN(O2745));
  NANDX1 G31542 (.A1(W10102), .A2(W9420), .ZN(O482));
  NANDX1 G31543 (.A1(W815), .A2(W9896), .ZN(W23334));
  NANDX1 G31544 (.A1(I1095), .A2(W2050), .ZN(O2746));
  NANDX1 G31545 (.A1(W4717), .A2(I701), .ZN(W11102));
  NANDX1 G31546 (.A1(I1342), .A2(I1343), .ZN(W671));
  NANDX1 G31547 (.A1(W23171), .A2(W20764), .ZN(W23337));
  NANDX1 G31548 (.A1(W5377), .A2(W21348), .ZN(W23340));
  NANDX1 G31549 (.A1(I1473), .A2(W1110), .ZN(W1387));
  NANDX1 G31550 (.A1(I616), .A2(I1960), .ZN(W1359));
  NANDX1 G31551 (.A1(W3929), .A2(W9610), .ZN(W9613));
  NANDX1 G31552 (.A1(W5477), .A2(I294), .ZN(W9614));
  NANDX1 G31553 (.A1(W9633), .A2(W13146), .ZN(O2748));
  NANDX1 G31554 (.A1(W2425), .A2(W3346), .ZN(W9616));
  NANDX1 G31555 (.A1(W9781), .A2(W13711), .ZN(W23352));
  NANDX1 G31556 (.A1(W2913), .A2(W24336), .ZN(O3076));
  NANDX1 G31557 (.A1(W8542), .A2(W2647), .ZN(W11091));
  NANDX1 G31558 (.A1(I366), .A2(W298), .ZN(W1378));
  NANDX1 G31559 (.A1(W18467), .A2(W8577), .ZN(W23359));
  NANDX1 G31560 (.A1(W18355), .A2(W10352), .ZN(O2750));
  NANDX1 G31561 (.A1(W22434), .A2(W2543), .ZN(W24413));
  NANDX1 G31562 (.A1(I1337), .A2(W6251), .ZN(W11089));
  NANDX1 G31563 (.A1(I1344), .A2(I1345), .ZN(W672));
  NANDX1 G31564 (.A1(I922), .A2(W3999), .ZN(W9925));
  NANDX1 G31565 (.A1(W89), .A2(W9670), .ZN(W23434));
  NANDX1 G31566 (.A1(I1425), .A2(I146), .ZN(W1320));
  NANDX1 G31567 (.A1(W20654), .A2(W21260), .ZN(W23421));
  NANDX1 G31568 (.A1(I1783), .A2(I27), .ZN(W1319));
  NANDX1 G31569 (.A1(W8680), .A2(W10820), .ZN(W23422));
  NANDX1 G31570 (.A1(W453), .A2(I967), .ZN(W1317));
  NANDX1 G31571 (.A1(W8911), .A2(W14835), .ZN(W23423));
  NANDX1 G31572 (.A1(W4683), .A2(W9635), .ZN(W9639));
  NANDX1 G31573 (.A1(W7789), .A2(W12562), .ZN(O2769));
  NANDX1 G31574 (.A1(I1391), .A2(W13845), .ZN(O3071));
  NANDX1 G31575 (.A1(W9469), .A2(W1702), .ZN(W11043));
  NANDX1 G31576 (.A1(W21883), .A2(W23014), .ZN(O2770));
  NANDX1 G31577 (.A1(W7188), .A2(W274), .ZN(W9917));
  NANDX1 G31578 (.A1(W19191), .A2(W2597), .ZN(O3070));
  NANDX1 G31579 (.A1(I682), .A2(W4775), .ZN(W10633));
  NANDX1 G31580 (.A1(W1650), .A2(W20026), .ZN(W23432));
  NANDX1 G31581 (.A1(W356), .A2(I816), .ZN(W1321));
  NANDX1 G31582 (.A1(I661), .A2(W14124), .ZN(W23436));
  NANDX1 G31583 (.A1(W6053), .A2(W23104), .ZN(O2773));
  NANDX1 G31584 (.A1(W5716), .A2(W22265), .ZN(W23438));
  NANDX1 G31585 (.A1(W1097), .A2(W2178), .ZN(W23439));
  NANDX1 G31586 (.A1(W8063), .A2(I300), .ZN(W23443));
  NANDX1 G31587 (.A1(W6474), .A2(W546), .ZN(W24389));
  NANDX1 G31588 (.A1(W2321), .A2(W4814), .ZN(W9911));
  NANDX1 G31589 (.A1(I1700), .A2(I737), .ZN(W1308));
  NANDX1 G31590 (.A1(W964), .A2(W1045), .ZN(O413));
  NANDX1 G31591 (.A1(I1724), .A2(W912), .ZN(W1305));
  NANDX1 G31592 (.A1(W22098), .A2(W22830), .ZN(O2776));
  NANDX1 G31593 (.A1(W3319), .A2(W9271), .ZN(O472));
  NANDX1 G31594 (.A1(W7161), .A2(W8226), .ZN(W11039));
  NANDX1 G31595 (.A1(W1058), .A2(W800), .ZN(O310));
  NANDX1 G31596 (.A1(I600), .A2(I351), .ZN(W1341));
  NANDX1 G31597 (.A1(W21353), .A2(W10255), .ZN(W23395));
  NANDX1 G31598 (.A1(W953), .A2(W636), .ZN(W1354));
  NANDX1 G31599 (.A1(W24381), .A2(W23261), .ZN(W24406));
  NANDX1 G31600 (.A1(W9027), .A2(W3718), .ZN(W9630));
  NANDX1 G31601 (.A1(W6438), .A2(W16132), .ZN(W24405));
  NANDX1 G31602 (.A1(W13745), .A2(W22415), .ZN(O2764));
  NANDX1 G31603 (.A1(I1496), .A2(W1346), .ZN(W1350));
  NANDX1 G31604 (.A1(I7), .A2(I1742), .ZN(W1349));
  NANDX1 G31605 (.A1(W11245), .A2(W13324), .ZN(W23404));
  NANDX1 G31606 (.A1(W22590), .A2(W22128), .ZN(W24404));
  NANDX1 G31607 (.A1(I1923), .A2(W9711), .ZN(W11063));
  NANDX1 G31608 (.A1(W1023), .A2(I160), .ZN(W1344));
  NANDX1 G31609 (.A1(W1735), .A2(W152), .ZN(O2767));
  NANDX1 G31610 (.A1(W6448), .A2(I601), .ZN(W10626));
  NANDX1 G31611 (.A1(W19714), .A2(W10726), .ZN(W23411));
  NANDX1 G31612 (.A1(W16312), .A2(W20341), .ZN(W24420));
  NANDX1 G31613 (.A1(I563), .A2(W1231), .ZN(W1337));
  NANDX1 G31614 (.A1(W4571), .A2(W5781), .ZN(W23412));
  NANDX1 G31615 (.A1(W1654), .A2(I1486), .ZN(O411));
  NANDX1 G31616 (.A1(W1119), .A2(I1952), .ZN(W1335));
  NANDX1 G31617 (.A1(W2978), .A2(W5448), .ZN(W11058));
  NANDX1 G31618 (.A1(W8732), .A2(W3603), .ZN(O339));
  NANDX1 G31619 (.A1(W7), .A2(I226), .ZN(W1332));
  NANDX1 G31620 (.A1(I956), .A2(W9183), .ZN(W11055));
  NANDX1 G31621 (.A1(W4220), .A2(W4296), .ZN(W10632));
  NANDX1 G31622 (.A1(I1374), .A2(I1375), .ZN(W687));
  NANDX1 G31623 (.A1(W7046), .A2(I168), .ZN(W9637));
  NANDX1 G31624 (.A1(I1376), .A2(I1377), .ZN(W688));
  NANDX1 G31625 (.A1(W6162), .A2(W6411), .ZN(W11052));
  NANDX1 G31626 (.A1(W16696), .A2(W2301), .ZN(W23420));
  NANDX1 G31627 (.A1(W2080), .A2(W11581), .ZN(O3090));
  NANDX1 G31628 (.A1(W2037), .A2(W9078), .ZN(W10598));
  NANDX1 G31629 (.A1(W5435), .A2(W1352), .ZN(W11134));
  NANDX1 G31630 (.A1(W1534), .A2(W7557), .ZN(W11133));
  NANDX1 G31631 (.A1(W11612), .A2(W7115), .ZN(W24464));
  NANDX1 G31632 (.A1(I385), .A2(I1080), .ZN(W1442));
  NANDX1 G31633 (.A1(W3274), .A2(W10518), .ZN(W23253));
  NANDX1 G31634 (.A1(W22608), .A2(W2315), .ZN(O3092));
  NANDX1 G31635 (.A1(I1505), .A2(W5581), .ZN(W11131));
  NANDX1 G31636 (.A1(W1301), .A2(W947), .ZN(W1441));
  NANDX1 G31637 (.A1(I1197), .A2(W909), .ZN(W1440));
  NANDX1 G31638 (.A1(W6492), .A2(W23088), .ZN(O2725));
  NANDX1 G31639 (.A1(I1292), .A2(I1293), .ZN(W646));
  NANDX1 G31640 (.A1(W201), .A2(I1913), .ZN(W1438));
  NANDX1 G31641 (.A1(W22084), .A2(W18212), .ZN(O2727));
  NANDX1 G31642 (.A1(W4768), .A2(W6908), .ZN(W10601));
  NANDX1 G31643 (.A1(W9410), .A2(W5762), .ZN(W9582));
  NANDX1 G31644 (.A1(W8410), .A2(W2878), .ZN(W9931));
  NANDX1 G31645 (.A1(I637), .A2(I1267), .ZN(W1436));
  NANDX1 G31646 (.A1(W12626), .A2(I907), .ZN(O2729));
  NANDX1 G31647 (.A1(W6200), .A2(W22003), .ZN(W23264));
  NANDX1 G31648 (.A1(I1743), .A2(W798), .ZN(W1434));
  NANDX1 G31649 (.A1(W10927), .A2(W2106), .ZN(W11130));
  NANDX1 G31650 (.A1(I1962), .A2(W583), .ZN(W1433));
  NANDX1 G31651 (.A1(I1913), .A2(I1250), .ZN(W10602));
  NANDX1 G31652 (.A1(W3896), .A2(I1200), .ZN(O2730));
  NANDX1 G31653 (.A1(W21419), .A2(I48), .ZN(O2731));
  NANDX1 G31654 (.A1(W13040), .A2(W22872), .ZN(W24456));
  NANDX1 G31655 (.A1(I710), .A2(W4706), .ZN(W10603));
  NANDX1 G31656 (.A1(I1298), .A2(I1299), .ZN(W649));
  NANDX1 G31657 (.A1(I1302), .A2(I1303), .ZN(W651));
  NANDX1 G31658 (.A1(I540), .A2(W5496), .ZN(O301));
  NANDX1 G31659 (.A1(W1252), .A2(I1639), .ZN(W11144));
  NANDX1 G31660 (.A1(W13528), .A2(W12668), .ZN(W24477));
  NANDX1 G31661 (.A1(W23065), .A2(W8713), .ZN(O3095));
  NANDX1 G31662 (.A1(I1544), .A2(W5842), .ZN(O484));
  NANDX1 G31663 (.A1(I144), .A2(W6983), .ZN(O2715));
  NANDX1 G31664 (.A1(W7653), .A2(I1994), .ZN(W9572));
  NANDX1 G31665 (.A1(W10326), .A2(W16825), .ZN(W24474));
  NANDX1 G31666 (.A1(W1507), .A2(W16103), .ZN(W23231));
  NANDX1 G31667 (.A1(I1264), .A2(I1265), .ZN(W632));
  NANDX1 G31668 (.A1(I1266), .A2(I1267), .ZN(W633));
  NANDX1 G31669 (.A1(W3568), .A2(W1234), .ZN(W10592));
  NANDX1 G31670 (.A1(W1261), .A2(W415), .ZN(W1461));
  NANDX1 G31671 (.A1(I1270), .A2(I1271), .ZN(W635));
  NANDX1 G31672 (.A1(W8074), .A2(W9077), .ZN(W10593));
  NANDX1 G31673 (.A1(W22135), .A2(W5744), .ZN(W24471));
  NANDX1 G31674 (.A1(W16449), .A2(W5669), .ZN(O2732));
  NANDX1 G31675 (.A1(W71), .A2(I1072), .ZN(W1458));
  NANDX1 G31676 (.A1(W6638), .A2(W11913), .ZN(W23238));
  NANDX1 G31677 (.A1(W3023), .A2(W19082), .ZN(W24470));
  NANDX1 G31678 (.A1(W3583), .A2(W3016), .ZN(W9933));
  NANDX1 G31679 (.A1(W17368), .A2(W4460), .ZN(O2719));
  NANDX1 G31680 (.A1(I991), .A2(I1435), .ZN(W24467));
  NANDX1 G31681 (.A1(I271), .A2(I1246), .ZN(W1456));
  NANDX1 G31682 (.A1(W679), .A2(W9306), .ZN(W9576));
  NANDX1 G31683 (.A1(W9107), .A2(W18237), .ZN(W23245));
  NANDX1 G31684 (.A1(W8856), .A2(I378), .ZN(W11138));
  NANDX1 G31685 (.A1(W286), .A2(I117), .ZN(W1450));
  NANDX1 G31686 (.A1(I1286), .A2(I1287), .ZN(W643));
  NANDX1 G31687 (.A1(W7811), .A2(W1942), .ZN(W9579));
  NANDX1 G31688 (.A1(W11683), .A2(W1538), .ZN(W24465));
  NANDX1 G31689 (.A1(I915), .A2(I916), .ZN(W1400));
  NANDX1 G31690 (.A1(I1546), .A2(W1193), .ZN(W23294));
  NANDX1 G31691 (.A1(I1322), .A2(I1323), .ZN(W661));
  NANDX1 G31692 (.A1(W21965), .A2(W23016), .ZN(W23298));
  NANDX1 G31693 (.A1(I806), .A2(I1784), .ZN(W1406));
  NANDX1 G31694 (.A1(W13670), .A2(W17576), .ZN(W23301));
  NANDX1 G31695 (.A1(W17286), .A2(W527), .ZN(O3082));
  NANDX1 G31696 (.A1(W5127), .A2(W8628), .ZN(W10609));
  NANDX1 G31697 (.A1(W18204), .A2(W3569), .ZN(W24430));
  NANDX1 G31698 (.A1(W20986), .A2(W21746), .ZN(W24429));
  NANDX1 G31699 (.A1(W5896), .A2(W3438), .ZN(W9606));
  NANDX1 G31700 (.A1(I1324), .A2(I1325), .ZN(W662));
  NANDX1 G31701 (.A1(W2240), .A2(W1462), .ZN(W23306));
  NANDX1 G31702 (.A1(I96), .A2(I565), .ZN(W1402));
  NANDX1 G31703 (.A1(W6866), .A2(W6579), .ZN(W10611));
  NANDX1 G31704 (.A1(W10326), .A2(W10140), .ZN(W11114));
  NANDX1 G31705 (.A1(I1056), .A2(W7062), .ZN(W23293));
  NANDX1 G31706 (.A1(I219), .A2(W8602), .ZN(W23312));
  NANDX1 G31707 (.A1(W21047), .A2(W8090), .ZN(O3080));
  NANDX1 G31708 (.A1(W6455), .A2(W5628), .ZN(W23313));
  NANDX1 G31709 (.A1(W21769), .A2(W12953), .ZN(O2741));
  NANDX1 G31710 (.A1(W17035), .A2(W9052), .ZN(W24425));
  NANDX1 G31711 (.A1(I1328), .A2(I1329), .ZN(W664));
  NANDX1 G31712 (.A1(W10098), .A2(W7182), .ZN(W11111));
  NANDX1 G31713 (.A1(W18669), .A2(W354), .ZN(W23316));
  NANDX1 G31714 (.A1(I1330), .A2(I1331), .ZN(W665));
  NANDX1 G31715 (.A1(I924), .A2(I120), .ZN(W1394));
  NANDX1 G31716 (.A1(W1112), .A2(W10880), .ZN(W24422));
  NANDX1 G31717 (.A1(W9987), .A2(W6297), .ZN(W10619));
  NANDX1 G31718 (.A1(I23), .A2(W10308), .ZN(W10620));
  NANDX1 G31719 (.A1(I1336), .A2(I1337), .ZN(W668));
  NANDX1 G31720 (.A1(W15946), .A2(W13366), .ZN(W24438));
  NANDX1 G31721 (.A1(I1304), .A2(I1305), .ZN(W652));
  NANDX1 G31722 (.A1(W226), .A2(I440), .ZN(W1426));
  NANDX1 G31723 (.A1(I1306), .A2(I1307), .ZN(W653));
  NANDX1 G31724 (.A1(W7784), .A2(W6769), .ZN(W9591));
  NANDX1 G31725 (.A1(W5294), .A2(W4561), .ZN(W9929));
  NANDX1 G31726 (.A1(W15994), .A2(W9683), .ZN(W24450));
  NANDX1 G31727 (.A1(W10142), .A2(W5224), .ZN(W10605));
  NANDX1 G31728 (.A1(W8422), .A2(I1019), .ZN(W10606));
  NANDX1 G31729 (.A1(W21642), .A2(W16887), .ZN(W23273));
  NANDX1 G31730 (.A1(W7103), .A2(W4194), .ZN(W9596));
  NANDX1 G31731 (.A1(W8775), .A2(W20265), .ZN(W24446));
  NANDX1 G31732 (.A1(W1339), .A2(W561), .ZN(W1421));
  NANDX1 G31733 (.A1(W4578), .A2(W23683), .ZN(O3085));
  NANDX1 G31734 (.A1(W9748), .A2(W2012), .ZN(W23276));
  NANDX1 G31735 (.A1(W10269), .A2(W9471), .ZN(W11036));
  NANDX1 G31736 (.A1(W10361), .A2(W19769), .ZN(W24434));
  NANDX1 G31737 (.A1(I1786), .A2(I1064), .ZN(W1413));
  NANDX1 G31738 (.A1(W6246), .A2(I861), .ZN(O304));
  NANDX1 G31739 (.A1(I1427), .A2(I690), .ZN(W1412));
  NANDX1 G31740 (.A1(W9291), .A2(W9879), .ZN(W9928));
  NANDX1 G31741 (.A1(W10127), .A2(W20466), .ZN(W23279));
  NANDX1 G31742 (.A1(W5696), .A2(W5940), .ZN(W9600));
  NANDX1 G31743 (.A1(I1802), .A2(W2777), .ZN(W9601));
  NANDX1 G31744 (.A1(I1318), .A2(I1319), .ZN(O5));
  NANDX1 G31745 (.A1(W2516), .A2(W4810), .ZN(W10608));
  NANDX1 G31746 (.A1(I1701), .A2(W1032), .ZN(W1410));
  NANDX1 G31747 (.A1(W3310), .A2(I1287), .ZN(W9603));
  NANDX1 G31748 (.A1(W230), .A2(I1325), .ZN(W1407));
  NANDX1 G31749 (.A1(W2536), .A2(W2513), .ZN(W23292));
  NANDX1 G31750 (.A1(W63), .A2(I516), .ZN(W1209));
  NANDX1 G31751 (.A1(I1519), .A2(W1020), .ZN(W9699));
  NANDX1 G31752 (.A1(W6286), .A2(W8015), .ZN(W10663));
  NANDX1 G31753 (.A1(W6780), .A2(W5198), .ZN(W10973));
  NANDX1 G31754 (.A1(W20225), .A2(W1946), .ZN(W23577));
  NANDX1 G31755 (.A1(W7232), .A2(I1758), .ZN(O459));
  NANDX1 G31756 (.A1(W152), .A2(W895), .ZN(W1211));
  NANDX1 G31757 (.A1(W6487), .A2(W598), .ZN(W9702));
  NANDX1 G31758 (.A1(I1440), .A2(I1441), .ZN(W720));
  NANDX1 G31759 (.A1(I812), .A2(I1589), .ZN(W10665));
  NANDX1 G31760 (.A1(I1305), .A2(W1858), .ZN(W10666));
  NANDX1 G31761 (.A1(W13733), .A2(W22503), .ZN(W23580));
  NANDX1 G31762 (.A1(W21203), .A2(W1987), .ZN(O3044));
  NANDX1 G31763 (.A1(W10510), .A2(W16955), .ZN(W24324));
  NANDX1 G31764 (.A1(W14007), .A2(W17755), .ZN(W24323));
  NANDX1 G31765 (.A1(W8503), .A2(W8904), .ZN(O457));
  NANDX1 G31766 (.A1(W7894), .A2(I1591), .ZN(W9697));
  NANDX1 G31767 (.A1(W7326), .A2(W6882), .ZN(W10962));
  NANDX1 G31768 (.A1(W18136), .A2(W4527), .ZN(W23585));
  NANDX1 G31769 (.A1(W1254), .A2(W8110), .ZN(W9707));
  NANDX1 G31770 (.A1(W9660), .A2(W9679), .ZN(W9709));
  NANDX1 G31771 (.A1(W5644), .A2(W9381), .ZN(W10960));
  NANDX1 G31772 (.A1(W143), .A2(W421), .ZN(O317));
  NANDX1 G31773 (.A1(W6130), .A2(W5265), .ZN(W10956));
  NANDX1 G31774 (.A1(I1446), .A2(I1447), .ZN(W723));
  NANDX1 G31775 (.A1(W3521), .A2(W4372), .ZN(W9711));
  NANDX1 G31776 (.A1(W19005), .A2(W5683), .ZN(W23594));
  NANDX1 G31777 (.A1(W594), .A2(W6234), .ZN(W10952));
  NANDX1 G31778 (.A1(W4151), .A2(W8742), .ZN(W23596));
  NANDX1 G31779 (.A1(I197), .A2(I1250), .ZN(W1201));
  NANDX1 G31780 (.A1(W3832), .A2(W3882), .ZN(W10951));
  NANDX1 G31781 (.A1(W20713), .A2(W10844), .ZN(O2817));
  NANDX1 G31782 (.A1(I1418), .A2(I1419), .ZN(W709));
  NANDX1 G31783 (.A1(W21012), .A2(W9980), .ZN(W23548));
  NANDX1 G31784 (.A1(W11429), .A2(W12659), .ZN(O2813));
  NANDX1 G31785 (.A1(W19413), .A2(W9073), .ZN(W23550));
  NANDX1 G31786 (.A1(W900), .A2(I106), .ZN(W1229));
  NANDX1 G31787 (.A1(W859), .A2(I1055), .ZN(W10997));
  NANDX1 G31788 (.A1(W7243), .A2(W3720), .ZN(W10995));
  NANDX1 G31789 (.A1(W11658), .A2(W13997), .ZN(W24343));
  NANDX1 G31790 (.A1(W4493), .A2(W304), .ZN(W9690));
  NANDX1 G31791 (.A1(W7424), .A2(W14481), .ZN(W24341));
  NANDX1 G31792 (.A1(W10098), .A2(W19312), .ZN(O3048));
  NANDX1 G31793 (.A1(W543), .A2(W889), .ZN(W1227));
  NANDX1 G31794 (.A1(W17203), .A2(I210), .ZN(O2815));
  NANDX1 G31795 (.A1(W1154), .A2(I1935), .ZN(W1226));
  NANDX1 G31796 (.A1(I1422), .A2(I1423), .ZN(W711));
  NANDX1 G31797 (.A1(W20954), .A2(W265), .ZN(O2824));
  NANDX1 G31798 (.A1(I1844), .A2(W802), .ZN(W1221));
  NANDX1 G31799 (.A1(W20315), .A2(W15185), .ZN(W23567));
  NANDX1 G31800 (.A1(W23406), .A2(W1022), .ZN(W24335));
  NANDX1 G31801 (.A1(W5771), .A2(W2767), .ZN(W10658));
  NANDX1 G31802 (.A1(W3295), .A2(W16704), .ZN(W24329));
  NANDX1 G31803 (.A1(W3903), .A2(W9717), .ZN(W10988));
  NANDX1 G31804 (.A1(I1434), .A2(I1435), .ZN(W717));
  NANDX1 G31805 (.A1(I1436), .A2(I1437), .ZN(W718));
  NANDX1 G31806 (.A1(W10555), .A2(W10388), .ZN(W10987));
  NANDX1 G31807 (.A1(W356), .A2(W6081), .ZN(W24328));
  NANDX1 G31808 (.A1(W3250), .A2(W10362), .ZN(W10982));
  NANDX1 G31809 (.A1(W22707), .A2(W11631), .ZN(W23569));
  NANDX1 G31810 (.A1(W16575), .A2(W16242), .ZN(W24327));
  NANDX1 G31811 (.A1(W5573), .A2(W196), .ZN(W9694));
  NANDX1 G31812 (.A1(W1848), .A2(W18236), .ZN(O2840));
  NANDX1 G31813 (.A1(W1109), .A2(I243), .ZN(W1182));
  NANDX1 G31814 (.A1(I1193), .A2(W8381), .ZN(O318));
  NANDX1 G31815 (.A1(W17644), .A2(W13213), .ZN(W24309));
  NANDX1 G31816 (.A1(W9582), .A2(W2361), .ZN(W9721));
  NANDX1 G31817 (.A1(W5051), .A2(W4969), .ZN(W10670));
  NANDX1 G31818 (.A1(I1460), .A2(I1461), .ZN(W730));
  NANDX1 G31819 (.A1(W4007), .A2(W1011), .ZN(W23640));
  NANDX1 G31820 (.A1(W10055), .A2(W606), .ZN(O2836));
  NANDX1 G31821 (.A1(W9689), .A2(W6146), .ZN(O333));
  NANDX1 G31822 (.A1(W16774), .A2(W12198), .ZN(O3040));
  NANDX1 G31823 (.A1(I1470), .A2(I1471), .ZN(W735));
  NANDX1 G31824 (.A1(W21747), .A2(W2446), .ZN(O2838));
  NANDX1 G31825 (.A1(W20177), .A2(W8639), .ZN(W23644));
  NANDX1 G31826 (.A1(W685), .A2(I1518), .ZN(W1174));
  NANDX1 G31827 (.A1(W10818), .A2(W18682), .ZN(W23646));
  NANDX1 G31828 (.A1(W21770), .A2(W7519), .ZN(O2835));
  NANDX1 G31829 (.A1(I1435), .A2(W22943), .ZN(W23648));
  NANDX1 G31830 (.A1(W12587), .A2(W10337), .ZN(W23649));
  NANDX1 G31831 (.A1(I1474), .A2(I1475), .ZN(W737));
  NANDX1 G31832 (.A1(W2425), .A2(I960), .ZN(W10940));
  NANDX1 G31833 (.A1(W5358), .A2(W3645), .ZN(W10672));
  NANDX1 G31834 (.A1(W10622), .A2(W11353), .ZN(W24299));
  NANDX1 G31835 (.A1(W8812), .A2(W6792), .ZN(W10938));
  NANDX1 G31836 (.A1(W17903), .A2(W9419), .ZN(W23651));
  NANDX1 G31837 (.A1(W6474), .A2(W21647), .ZN(W23652));
  NANDX1 G31838 (.A1(I351), .A2(W3067), .ZN(W23654));
  NANDX1 G31839 (.A1(W4943), .A2(W18680), .ZN(W23655));
  NANDX1 G31840 (.A1(I1476), .A2(I1477), .ZN(W738));
  NANDX1 G31841 (.A1(I1866), .A2(W21338), .ZN(W23656));
  NANDX1 G31842 (.A1(I1692), .A2(I1993), .ZN(W1170));
  NANDX1 G31843 (.A1(I347), .A2(I1444), .ZN(W1189));
  NANDX1 G31844 (.A1(W2237), .A2(W7469), .ZN(W9713));
  NANDX1 G31845 (.A1(W7842), .A2(W10173), .ZN(W23600));
  NANDX1 G31846 (.A1(W5683), .A2(I1034), .ZN(W9890));
  NANDX1 G31847 (.A1(I481), .A2(W1132), .ZN(W1198));
  NANDX1 G31848 (.A1(W21646), .A2(W5525), .ZN(W24319));
  NANDX1 G31849 (.A1(I896), .A2(W842), .ZN(O2826));
  NANDX1 G31850 (.A1(I489), .A2(I1281), .ZN(W1195));
  NANDX1 G31851 (.A1(W5279), .A2(I1454), .ZN(W10667));
  NANDX1 G31852 (.A1(W2875), .A2(W5806), .ZN(W24318));
  NANDX1 G31853 (.A1(W4994), .A2(W18487), .ZN(O2827));
  NANDX1 G31854 (.A1(W5603), .A2(W8416), .ZN(W10947));
  NANDX1 G31855 (.A1(I1634), .A2(I218), .ZN(W1192));
  NANDX1 G31856 (.A1(I626), .A2(W14174), .ZN(W24317));
  NANDX1 G31857 (.A1(W60), .A2(I398), .ZN(W1191));
  NANDX1 G31858 (.A1(W13892), .A2(W18213), .ZN(W23612));
  NANDX1 G31859 (.A1(I1042), .A2(W774), .ZN(W1230));
  NANDX1 G31860 (.A1(W22400), .A2(W137), .ZN(W23616));
  NANDX1 G31861 (.A1(W816), .A2(W7525), .ZN(W10946));
  NANDX1 G31862 (.A1(W17435), .A2(W14780), .ZN(O2830));
  NANDX1 G31863 (.A1(W9335), .A2(W9880), .ZN(W10944));
  NANDX1 G31864 (.A1(W16931), .A2(W15636), .ZN(W23619));
  NANDX1 G31865 (.A1(W530), .A2(W22292), .ZN(W23620));
  NANDX1 G31866 (.A1(I1452), .A2(I1453), .ZN(W726));
  NANDX1 G31867 (.A1(I564), .A2(I1513), .ZN(W1186));
  NANDX1 G31868 (.A1(I1454), .A2(I1455), .ZN(W727));
  NANDX1 G31869 (.A1(I1456), .A2(I1457), .ZN(W728));
  NANDX1 G31870 (.A1(W10225), .A2(W3644), .ZN(W23630));
  NANDX1 G31871 (.A1(W4955), .A2(W2145), .ZN(W23631));
  NANDX1 G31872 (.A1(I1927), .A2(I1535), .ZN(W1184));
  NANDX1 G31873 (.A1(I764), .A2(W1016), .ZN(W1183));
  NANDX1 G31874 (.A1(W4607), .A2(W7080), .ZN(W10644));
  NANDX1 G31875 (.A1(W5736), .A2(W12682), .ZN(W23471));
  NANDX1 G31876 (.A1(W4625), .A2(W8991), .ZN(W11015));
  NANDX1 G31877 (.A1(I1780), .A2(W7776), .ZN(W23474));
  NANDX1 G31878 (.A1(W200), .A2(I1599), .ZN(W1288));
  NANDX1 G31879 (.A1(I1163), .A2(I1452), .ZN(W1287));
  NANDX1 G31880 (.A1(W8815), .A2(W5273), .ZN(O415));
  NANDX1 G31881 (.A1(I23), .A2(I624), .ZN(W1283));
  NANDX1 G31882 (.A1(I1148), .A2(I478), .ZN(W1281));
  NANDX1 G31883 (.A1(I1166), .A2(I1536), .ZN(W1279));
  NANDX1 G31884 (.A1(W17365), .A2(W157), .ZN(W23483));
  NANDX1 G31885 (.A1(W3661), .A2(W7000), .ZN(W9664));
  NANDX1 G31886 (.A1(W5528), .A2(W6588), .ZN(W9665));
  NANDX1 G31887 (.A1(W15783), .A2(W8469), .ZN(W24367));
  NANDX1 G31888 (.A1(W2489), .A2(W9663), .ZN(O335));
  NANDX1 G31889 (.A1(W10470), .A2(W3411), .ZN(W10643));
  NANDX1 G31890 (.A1(W5996), .A2(W6255), .ZN(W11019));
  NANDX1 G31891 (.A1(I1406), .A2(I1407), .ZN(W703));
  NANDX1 G31892 (.A1(W6362), .A2(W3665), .ZN(W23488));
  NANDX1 G31893 (.A1(I315), .A2(I762), .ZN(W1274));
  NANDX1 G31894 (.A1(W9190), .A2(W2637), .ZN(O2794));
  NANDX1 G31895 (.A1(W2532), .A2(I874), .ZN(W9668));
  NANDX1 G31896 (.A1(I169), .A2(I1347), .ZN(W1273));
  NANDX1 G31897 (.A1(W2764), .A2(W13192), .ZN(W23493));
  NANDX1 G31898 (.A1(I1408), .A2(I1409), .ZN(W704));
  NANDX1 G31899 (.A1(W16777), .A2(W9826), .ZN(O2795));
  NANDX1 G31900 (.A1(W7538), .A2(W4927), .ZN(O464));
  NANDX1 G31901 (.A1(I813), .A2(W818), .ZN(W1268));
  NANDX1 G31902 (.A1(W7754), .A2(W2761), .ZN(W9669));
  NANDX1 G31903 (.A1(W16000), .A2(W12886), .ZN(O2799));
  NANDX1 G31904 (.A1(W16397), .A2(W2494), .ZN(W23502));
  NANDX1 G31905 (.A1(W8777), .A2(W4041), .ZN(O2784));
  NANDX1 G31906 (.A1(I659), .A2(W12912), .ZN(W23450));
  NANDX1 G31907 (.A1(I491), .A2(W8033), .ZN(W11033));
  NANDX1 G31908 (.A1(W8152), .A2(W3646), .ZN(W11032));
  NANDX1 G31909 (.A1(W4644), .A2(W1925), .ZN(O337));
  NANDX1 G31910 (.A1(W344), .A2(W7095), .ZN(W24387));
  NANDX1 G31911 (.A1(W2574), .A2(W7775), .ZN(W9648));
  NANDX1 G31912 (.A1(W6203), .A2(W12564), .ZN(W24384));
  NANDX1 G31913 (.A1(I1384), .A2(I1385), .ZN(W692));
  NANDX1 G31914 (.A1(W3015), .A2(W22585), .ZN(W23455));
  NANDX1 G31915 (.A1(W22321), .A2(W17949), .ZN(W24380));
  NANDX1 G31916 (.A1(W1737), .A2(I1210), .ZN(O2781));
  NANDX1 G31917 (.A1(W6797), .A2(W4427), .ZN(W11028));
  NANDX1 G31918 (.A1(W1231), .A2(I1966), .ZN(W1297));
  NANDX1 G31919 (.A1(W9163), .A2(W6435), .ZN(O312));
  NANDX1 G31920 (.A1(W307), .A2(W7710), .ZN(W9908));
  NANDX1 G31921 (.A1(W8894), .A2(W20767), .ZN(O3056));
  NANDX1 G31922 (.A1(I1388), .A2(I1389), .ZN(W694));
  NANDX1 G31923 (.A1(I518), .A2(I1251), .ZN(W1295));
  NANDX1 G31924 (.A1(W20562), .A2(W17978), .ZN(W23465));
  NANDX1 G31925 (.A1(I82), .A2(I950), .ZN(W1294));
  NANDX1 G31926 (.A1(I1190), .A2(W9333), .ZN(W11026));
  NANDX1 G31927 (.A1(W1124), .A2(W200), .ZN(O3064));
  NANDX1 G31928 (.A1(I1394), .A2(I1395), .ZN(W697));
  NANDX1 G31929 (.A1(I1777), .A2(W5119), .ZN(O469));
  NANDX1 G31930 (.A1(W19044), .A2(W7514), .ZN(W23467));
  NANDX1 G31931 (.A1(W7972), .A2(W17145), .ZN(O3062));
  NANDX1 G31932 (.A1(W6635), .A2(W8691), .ZN(W9659));
  NANDX1 G31933 (.A1(I1918), .A2(W4169), .ZN(W11021));
  NANDX1 G31934 (.A1(W7789), .A2(W3531), .ZN(O336));
  NANDX1 G31935 (.A1(W14234), .A2(W8580), .ZN(W23470));
  NANDX1 G31936 (.A1(W10981), .A2(W129), .ZN(O2809));
  NANDX1 G31937 (.A1(W254), .A2(W17876), .ZN(O2806));
  NANDX1 G31938 (.A1(W783), .A2(I863), .ZN(W1248));
  NANDX1 G31939 (.A1(I1743), .A2(W861), .ZN(W1246));
  NANDX1 G31940 (.A1(W13151), .A2(W13227), .ZN(W23527));
  NANDX1 G31941 (.A1(W18429), .A2(W15090), .ZN(W23528));
  NANDX1 G31942 (.A1(W2581), .A2(W10519), .ZN(W10651));
  NANDX1 G31943 (.A1(W3021), .A2(W13517), .ZN(W23529));
  NANDX1 G31944 (.A1(I1066), .A2(I876), .ZN(W1242));
  NANDX1 G31945 (.A1(W15194), .A2(W14000), .ZN(O2807));
  NANDX1 G31946 (.A1(W8134), .A2(I652), .ZN(W9681));
  NANDX1 G31947 (.A1(W10716), .A2(W18706), .ZN(O2808));
  NANDX1 G31948 (.A1(I91), .A2(W7852), .ZN(W11004));
  NANDX1 G31949 (.A1(W9453), .A2(I196), .ZN(W10653));
  NANDX1 G31950 (.A1(W192), .A2(W739), .ZN(W1237));
  NANDX1 G31951 (.A1(I1566), .A2(W6353), .ZN(W23534));
  NANDX1 G31952 (.A1(W5974), .A2(I1793), .ZN(W9897));
  NANDX1 G31953 (.A1(W2047), .A2(W15736), .ZN(W23536));
  NANDX1 G31954 (.A1(W989), .A2(I459), .ZN(W1235));
  NANDX1 G31955 (.A1(W3742), .A2(W9695), .ZN(W24347));
  NANDX1 G31956 (.A1(W6019), .A2(W7504), .ZN(O334));
  NANDX1 G31957 (.A1(W3602), .A2(W6156), .ZN(W9683));
  NANDX1 G31958 (.A1(W17240), .A2(I1792), .ZN(O2810));
  NANDX1 G31959 (.A1(W8794), .A2(W19953), .ZN(W23539));
  NANDX1 G31960 (.A1(W2374), .A2(W6984), .ZN(W9684));
  NANDX1 G31961 (.A1(W2257), .A2(W462), .ZN(W23542));
  NANDX1 G31962 (.A1(W3738), .A2(W8134), .ZN(W10998));
  NANDX1 G31963 (.A1(W1460), .A2(W19010), .ZN(W23543));
  NANDX1 G31964 (.A1(W3867), .A2(W4894), .ZN(W9686));
  NANDX1 G31965 (.A1(I608), .A2(W458), .ZN(W1231));
  NANDX1 G31966 (.A1(W5513), .A2(W20671), .ZN(W23546));
  NANDX1 G31967 (.A1(W7981), .A2(W16377), .ZN(W23512));
  NANDX1 G31968 (.A1(W611), .A2(I75), .ZN(W1265));
  NANDX1 G31969 (.A1(W868), .A2(I1444), .ZN(W1263));
  NANDX1 G31970 (.A1(W5533), .A2(W4931), .ZN(W23504));
  NANDX1 G31971 (.A1(W1004), .A2(I1067), .ZN(W1262));
  NANDX1 G31972 (.A1(I1495), .A2(W1088), .ZN(W1261));
  NANDX1 G31973 (.A1(W989), .A2(W4608), .ZN(O463));
  NANDX1 G31974 (.A1(I1859), .A2(W10622), .ZN(W24358));
  NANDX1 G31975 (.A1(W10654), .A2(W2084), .ZN(W11009));
  NANDX1 G31976 (.A1(W16423), .A2(W20410), .ZN(W23507));
  NANDX1 G31977 (.A1(W5812), .A2(W20460), .ZN(W23508));
  NANDX1 G31978 (.A1(I756), .A2(W1187), .ZN(W1256));
  NANDX1 G31979 (.A1(W4573), .A2(I1522), .ZN(W24357));
  NANDX1 G31980 (.A1(W9761), .A2(W10648), .ZN(W23509));
  NANDX1 G31981 (.A1(W6725), .A2(W13016), .ZN(W23510));
  NANDX1 G31982 (.A1(W6396), .A2(W5092), .ZN(W8782));
  NANDX1 G31983 (.A1(I400), .A2(W2), .ZN(W1254));
  NANDX1 G31984 (.A1(W20654), .A2(I934), .ZN(W24356));
  NANDX1 G31985 (.A1(I360), .A2(W32), .ZN(W1252));
  NANDX1 G31986 (.A1(W19704), .A2(W4156), .ZN(O2802));
  NANDX1 G31987 (.A1(I879), .A2(W20256), .ZN(W24355));
  NANDX1 G31988 (.A1(W17207), .A2(W19032), .ZN(W24354));
  NANDX1 G31989 (.A1(W22223), .A2(W22100), .ZN(W23517));
  NANDX1 G31990 (.A1(W15929), .A2(W17866), .ZN(W24353));
  NANDX1 G31991 (.A1(W17079), .A2(W21995), .ZN(W23518));
  NANDX1 G31992 (.A1(W13186), .A2(W13758), .ZN(W23520));
  NANDX1 G31993 (.A1(W5494), .A2(W18562), .ZN(O2803));
  NANDX1 G31994 (.A1(W5216), .A2(W9648), .ZN(O2804));
  NANDX1 G31995 (.A1(W3381), .A2(W538), .ZN(W10648));
  NANDX1 G31996 (.A1(W6270), .A2(I1264), .ZN(W10650));
  NANDX1 G31997 (.A1(W14495), .A2(W18663), .ZN(O3302));
  NANDX1 G31998 (.A1(W8037), .A2(W8447), .ZN(W21340));
  NANDX1 G31999 (.A1(W3272), .A2(I1402), .ZN(W8965));
  NANDX1 G32000 (.A1(W301), .A2(W1836), .ZN(W2737));
  NANDX1 G32001 (.A1(W1078), .A2(W7157), .ZN(W8967));
  NANDX1 G32002 (.A1(W2481), .A2(I74), .ZN(W2736));
  NANDX1 G32003 (.A1(I284), .A2(I285), .ZN(W142));
  NANDX1 G32004 (.A1(W713), .A2(W157), .ZN(W2734));
  NANDX1 G32005 (.A1(W1273), .A2(W7557), .ZN(W12032));
  NANDX1 G32006 (.A1(I1112), .A2(W851), .ZN(W10298));
  NANDX1 G32007 (.A1(W20962), .A2(W4461), .ZN(W21351));
  NANDX1 G32008 (.A1(W8915), .A2(W13959), .ZN(W21352));
  NANDX1 G32009 (.A1(I539), .A2(W4330), .ZN(W25105));
  NANDX1 G32010 (.A1(W949), .A2(W2557), .ZN(W2731));
  NANDX1 G32011 (.A1(W15927), .A2(W9566), .ZN(W21356));
  NANDX1 G32012 (.A1(I1738), .A2(W524), .ZN(O2224));
  NANDX1 G32013 (.A1(W7827), .A2(W16555), .ZN(W21339));
  NANDX1 G32014 (.A1(W3690), .A2(W5418), .ZN(W8971));
  NANDX1 G32015 (.A1(W4380), .A2(W1179), .ZN(O3300));
  NANDX1 G32016 (.A1(W8842), .A2(W11416), .ZN(W21364));
  NANDX1 G32017 (.A1(I543), .A2(I1352), .ZN(W8973));
  NANDX1 G32018 (.A1(W7215), .A2(W1185), .ZN(W12030));
  NANDX1 G32019 (.A1(W7073), .A2(W3891), .ZN(W12029));
  NANDX1 G32020 (.A1(W8127), .A2(W2842), .ZN(W12028));
  NANDX1 G32021 (.A1(I288), .A2(I289), .ZN(W144));
  NANDX1 G32022 (.A1(I290), .A2(I291), .ZN(W145));
  NANDX1 G32023 (.A1(W699), .A2(I1593), .ZN(W2727));
  NANDX1 G32024 (.A1(W5134), .A2(W3067), .ZN(O560));
  NANDX1 G32025 (.A1(W18557), .A2(W17693), .ZN(W25099));
  NANDX1 G32026 (.A1(W5670), .A2(W12529), .ZN(O2227));
  NANDX1 G32027 (.A1(W6012), .A2(W9414), .ZN(W12024));
  NANDX1 G32028 (.A1(W9765), .A2(W1918), .ZN(W12037));
  NANDX1 G32029 (.A1(W24420), .A2(W1051), .ZN(O3307));
  NANDX1 G32030 (.A1(W11426), .A2(W7944), .ZN(W12042));
  NANDX1 G32031 (.A1(I753), .A2(W6815), .ZN(W10295));
  NANDX1 G32032 (.A1(W1424), .A2(I1883), .ZN(W25118));
  NANDX1 G32033 (.A1(I1437), .A2(W2657), .ZN(W2756));
  NANDX1 G32034 (.A1(W11932), .A2(W6270), .ZN(W21313));
  NANDX1 G32035 (.A1(W3462), .A2(W19608), .ZN(W21315));
  NANDX1 G32036 (.A1(W2490), .A2(W681), .ZN(W2753));
  NANDX1 G32037 (.A1(I276), .A2(I277), .ZN(W138));
  NANDX1 G32038 (.A1(W1347), .A2(W2166), .ZN(W2747));
  NANDX1 G32039 (.A1(I1619), .A2(I471), .ZN(W2746));
  NANDX1 G32040 (.A1(W1227), .A2(W10884), .ZN(W25115));
  NANDX1 G32041 (.A1(W6031), .A2(W6611), .ZN(W12038));
  NANDX1 G32042 (.A1(W20076), .A2(I1739), .ZN(W21321));
  NANDX1 G32043 (.A1(W7533), .A2(W20057), .ZN(W21372));
  NANDX1 G32044 (.A1(W1432), .A2(I1196), .ZN(W2743));
  NANDX1 G32045 (.A1(W4433), .A2(W2602), .ZN(W8960));
  NANDX1 G32046 (.A1(W16376), .A2(W622), .ZN(W25113));
  NANDX1 G32047 (.A1(W1153), .A2(W1496), .ZN(W2742));
  NANDX1 G32048 (.A1(W19415), .A2(W19574), .ZN(O2216));
  NANDX1 G32049 (.A1(W2727), .A2(W2005), .ZN(W25112));
  NANDX1 G32050 (.A1(W165), .A2(W780), .ZN(W2740));
  NANDX1 G32051 (.A1(W631), .A2(W1167), .ZN(W2739));
  NANDX1 G32052 (.A1(W9236), .A2(W942), .ZN(W10124));
  NANDX1 G32053 (.A1(W11517), .A2(W20611), .ZN(W21332));
  NANDX1 G32054 (.A1(W2835), .A2(W21564), .ZN(O3305));
  NANDX1 G32055 (.A1(W2218), .A2(W11481), .ZN(W21333));
  NANDX1 G32056 (.A1(W315), .A2(W1591), .ZN(W2738));
  NANDX1 G32057 (.A1(W20891), .A2(W613), .ZN(W21336));
  NANDX1 G32058 (.A1(I476), .A2(W1189), .ZN(W2689));
  NANDX1 G32059 (.A1(W14583), .A2(W5906), .ZN(W21404));
  NANDX1 G32060 (.A1(I300), .A2(I301), .ZN(W150));
  NANDX1 G32061 (.A1(I302), .A2(I303), .ZN(W151));
  NANDX1 G32062 (.A1(I304), .A2(I305), .ZN(W152));
  NANDX1 G32063 (.A1(W8706), .A2(W7547), .ZN(W8987));
  NANDX1 G32064 (.A1(W2700), .A2(W4134), .ZN(W10114));
  NANDX1 G32065 (.A1(W1745), .A2(I1773), .ZN(W8989));
  NANDX1 G32066 (.A1(W1647), .A2(I468), .ZN(O380));
  NANDX1 G32067 (.A1(W3922), .A2(W11998), .ZN(W12001));
  NANDX1 G32068 (.A1(I308), .A2(I309), .ZN(W154));
  NANDX1 G32069 (.A1(W185), .A2(W12965), .ZN(O2237));
  NANDX1 G32070 (.A1(W2193), .A2(I246), .ZN(W2695));
  NANDX1 G32071 (.A1(I128), .A2(W15839), .ZN(O2239));
  NANDX1 G32072 (.A1(W4782), .A2(W6907), .ZN(W8992));
  NANDX1 G32073 (.A1(W884), .A2(I1569), .ZN(W2692));
  NANDX1 G32074 (.A1(I298), .A2(I299), .ZN(W149));
  NANDX1 G32075 (.A1(I312), .A2(I313), .ZN(W156));
  NANDX1 G32076 (.A1(W2698), .A2(W6278), .ZN(O2240));
  NANDX1 G32077 (.A1(I679), .A2(W1310), .ZN(W11997));
  NANDX1 G32078 (.A1(W10632), .A2(W4555), .ZN(W11995));
  NANDX1 G32079 (.A1(W15604), .A2(W1565), .ZN(O3290));
  NANDX1 G32080 (.A1(W21093), .A2(W5711), .ZN(W25082));
  NANDX1 G32081 (.A1(W6552), .A2(W9988), .ZN(W11994));
  NANDX1 G32082 (.A1(W2628), .A2(W15055), .ZN(O2242));
  NANDX1 G32083 (.A1(W742), .A2(I1571), .ZN(W8993));
  NANDX1 G32084 (.A1(I314), .A2(I315), .ZN(W157));
  NANDX1 G32085 (.A1(I435), .A2(W1405), .ZN(W2684));
  NANDX1 G32086 (.A1(I318), .A2(I319), .ZN(W159));
  NANDX1 G32087 (.A1(W2569), .A2(I943), .ZN(W2683));
  NANDX1 G32088 (.A1(I1762), .A2(W20947), .ZN(W21429));
  NANDX1 G32089 (.A1(W8945), .A2(W621), .ZN(W10116));
  NANDX1 G32090 (.A1(W10191), .A2(W1302), .ZN(W12023));
  NANDX1 G32091 (.A1(W8477), .A2(W2257), .ZN(O2228));
  NANDX1 G32092 (.A1(W15440), .A2(W8677), .ZN(W21376));
  NANDX1 G32093 (.A1(W11194), .A2(W4946), .ZN(O3297));
  NANDX1 G32094 (.A1(W18644), .A2(W2524), .ZN(W25096));
  NANDX1 G32095 (.A1(I1702), .A2(W2897), .ZN(O558));
  NANDX1 G32096 (.A1(W4046), .A2(W534), .ZN(W21378));
  NANDX1 G32097 (.A1(W6979), .A2(I70), .ZN(O379));
  NANDX1 G32098 (.A1(I17), .A2(W15605), .ZN(W21380));
  NANDX1 G32099 (.A1(W622), .A2(W989), .ZN(W8981));
  NANDX1 G32100 (.A1(W2282), .A2(W1111), .ZN(W2719));
  NANDX1 G32101 (.A1(W2986), .A2(W300), .ZN(W12015));
  NANDX1 G32102 (.A1(W7748), .A2(W5091), .ZN(W8983));
  NANDX1 G32103 (.A1(I1281), .A2(W898), .ZN(W2709));
  NANDX1 G32104 (.A1(W3103), .A2(W9), .ZN(W10292));
  NANDX1 G32105 (.A1(W2799), .A2(W11175), .ZN(W12012));
  NANDX1 G32106 (.A1(W2589), .A2(W128), .ZN(W2707));
  NANDX1 G32107 (.A1(W18197), .A2(W12504), .ZN(O2233));
  NANDX1 G32108 (.A1(W8621), .A2(W11952), .ZN(W12011));
  NANDX1 G32109 (.A1(W5511), .A2(W16646), .ZN(W25094));
  NANDX1 G32110 (.A1(W20469), .A2(W17406), .ZN(O2236));
  NANDX1 G32111 (.A1(I296), .A2(I297), .ZN(W148));
  NANDX1 G32112 (.A1(W219), .A2(W4620), .ZN(W8985));
  NANDX1 G32113 (.A1(W3392), .A2(W210), .ZN(W12006));
  NANDX1 G32114 (.A1(W16885), .A2(W15221), .ZN(W21400));
  NANDX1 G32115 (.A1(W2190), .A2(W5245), .ZN(W25093));
  NANDX1 G32116 (.A1(I1975), .A2(W608), .ZN(W2704));
  NANDX1 G32117 (.A1(W5190), .A2(W19335), .ZN(W21402));
  NANDX1 G32118 (.A1(W14784), .A2(W13749), .ZN(W21403));
  NANDX1 G32119 (.A1(W6649), .A2(W5849), .ZN(O3315));
  NANDX1 G32120 (.A1(W19149), .A2(W7142), .ZN(W21221));
  NANDX1 G32121 (.A1(I455), .A2(W453), .ZN(W2809));
  NANDX1 G32122 (.A1(W821), .A2(W847), .ZN(W2808));
  NANDX1 G32123 (.A1(W21638), .A2(W15943), .ZN(O3316));
  NANDX1 G32124 (.A1(W868), .A2(W16115), .ZN(O2186));
  NANDX1 G32125 (.A1(W18384), .A2(W1150), .ZN(W21225));
  NANDX1 G32126 (.A1(W2059), .A2(W6251), .ZN(W8924));
  NANDX1 G32127 (.A1(W7204), .A2(I1648), .ZN(W12072));
  NANDX1 G32128 (.A1(W13130), .A2(W18049), .ZN(W21231));
  NANDX1 G32129 (.A1(W2401), .A2(I652), .ZN(W2805));
  NANDX1 G32130 (.A1(W1623), .A2(W2648), .ZN(W2802));
  NANDX1 G32131 (.A1(W11112), .A2(I564), .ZN(W12071));
  NANDX1 G32132 (.A1(I658), .A2(W82), .ZN(W2799));
  NANDX1 G32133 (.A1(I1830), .A2(W2750), .ZN(W8925));
  NANDX1 G32134 (.A1(W4528), .A2(W20856), .ZN(W21235));
  NANDX1 G32135 (.A1(W18494), .A2(W14036), .ZN(O2185));
  NANDX1 G32136 (.A1(W5861), .A2(W3412), .ZN(W8926));
  NANDX1 G32137 (.A1(I1002), .A2(I1087), .ZN(W2796));
  NANDX1 G32138 (.A1(W4047), .A2(W11314), .ZN(W21239));
  NANDX1 G32139 (.A1(I917), .A2(I1711), .ZN(W2795));
  NANDX1 G32140 (.A1(W2536), .A2(W1512), .ZN(W2793));
  NANDX1 G32141 (.A1(I220), .A2(I221), .ZN(W110));
  NANDX1 G32142 (.A1(W16539), .A2(W2742), .ZN(W25149));
  NANDX1 G32143 (.A1(W17991), .A2(W2359), .ZN(O2191));
  NANDX1 G32144 (.A1(I222), .A2(I223), .ZN(W111));
  NANDX1 G32145 (.A1(I226), .A2(I227), .ZN(W113));
  NANDX1 G32146 (.A1(I1156), .A2(I700), .ZN(W2790));
  NANDX1 G32147 (.A1(W2267), .A2(W2372), .ZN(W2789));
  NANDX1 G32148 (.A1(I679), .A2(I474), .ZN(W2788));
  NANDX1 G32149 (.A1(W2468), .A2(I1589), .ZN(W2787));
  NANDX1 G32150 (.A1(W2500), .A2(W1351), .ZN(W2819));
  NANDX1 G32151 (.A1(W4054), .A2(W6946), .ZN(W8908));
  NANDX1 G32152 (.A1(W4053), .A2(W10217), .ZN(W21193));
  NANDX1 G32153 (.A1(W18231), .A2(W8764), .ZN(O2179));
  NANDX1 G32154 (.A1(I1981), .A2(W221), .ZN(W2827));
  NANDX1 G32155 (.A1(I128), .A2(W292), .ZN(W2826));
  NANDX1 G32156 (.A1(I206), .A2(I207), .ZN(W103));
  NANDX1 G32157 (.A1(W9352), .A2(W3159), .ZN(W21198));
  NANDX1 G32158 (.A1(W2107), .A2(I1317), .ZN(W2824));
  NANDX1 G32159 (.A1(I208), .A2(I209), .ZN(W104));
  NANDX1 G32160 (.A1(W5524), .A2(W19028), .ZN(W21200));
  NANDX1 G32161 (.A1(W13740), .A2(W12885), .ZN(W25164));
  NANDX1 G32162 (.A1(I791), .A2(W13277), .ZN(W21201));
  NANDX1 G32163 (.A1(W9401), .A2(W6624), .ZN(W25163));
  NANDX1 G32164 (.A1(W2645), .A2(W7871), .ZN(W10132));
  NANDX1 G32165 (.A1(W7428), .A2(W17308), .ZN(O2193));
  NANDX1 G32166 (.A1(W10637), .A2(W16775), .ZN(O2182));
  NANDX1 G32167 (.A1(W13609), .A2(W12047), .ZN(O2183));
  NANDX1 G32168 (.A1(W10195), .A2(W1417), .ZN(W12082));
  NANDX1 G32169 (.A1(W11514), .A2(W13622), .ZN(W21208));
  NANDX1 G32170 (.A1(W10695), .A2(W11268), .ZN(W12077));
  NANDX1 G32171 (.A1(I212), .A2(I213), .ZN(W106));
  NANDX1 G32172 (.A1(I214), .A2(I215), .ZN(W107));
  NANDX1 G32173 (.A1(W1702), .A2(I1500), .ZN(W2814));
  NANDX1 G32174 (.A1(W2540), .A2(W1511), .ZN(W2812));
  NANDX1 G32175 (.A1(W5482), .A2(I1743), .ZN(W8916));
  NANDX1 G32176 (.A1(I1073), .A2(I748), .ZN(W8919));
  NANDX1 G32177 (.A1(W4746), .A2(W619), .ZN(W8921));
  NANDX1 G32178 (.A1(I1323), .A2(W74), .ZN(W2811));
  NANDX1 G32179 (.A1(I826), .A2(W24089), .ZN(W25157));
  NANDX1 G32180 (.A1(W8624), .A2(W6778), .ZN(W21292));
  NANDX1 G32181 (.A1(W7580), .A2(W19350), .ZN(W21275));
  NANDX1 G32182 (.A1(I254), .A2(I255), .ZN(W127));
  NANDX1 G32183 (.A1(W21955), .A2(W18502), .ZN(O3311));
  NANDX1 G32184 (.A1(I258), .A2(I259), .ZN(W129));
  NANDX1 G32185 (.A1(W2004), .A2(W1672), .ZN(W2770));
  NANDX1 G32186 (.A1(W1744), .A2(I588), .ZN(W21281));
  NANDX1 G32187 (.A1(W271), .A2(I1704), .ZN(W8943));
  NANDX1 G32188 (.A1(W907), .A2(I474), .ZN(W8944));
  NANDX1 G32189 (.A1(W13318), .A2(W8059), .ZN(W21287));
  NANDX1 G32190 (.A1(W5364), .A2(W6454), .ZN(O378));
  NANDX1 G32191 (.A1(W7121), .A2(W11757), .ZN(W21289));
  NANDX1 G32192 (.A1(W1844), .A2(W9295), .ZN(W12048));
  NANDX1 G32193 (.A1(W7670), .A2(W9359), .ZN(W10128));
  NANDX1 G32194 (.A1(W8901), .A2(W3926), .ZN(W8946));
  NANDX1 G32195 (.A1(W10103), .A2(W1169), .ZN(W10284));
  NANDX1 G32196 (.A1(W14128), .A2(W9273), .ZN(W21293));
  NANDX1 G32197 (.A1(W5922), .A2(I1318), .ZN(W21294));
  NANDX1 G32198 (.A1(W23184), .A2(W638), .ZN(O3310));
  NANDX1 G32199 (.A1(I268), .A2(I269), .ZN(W134));
  NANDX1 G32200 (.A1(W2753), .A2(W2852), .ZN(W8947));
  NANDX1 G32201 (.A1(W10227), .A2(W4103), .ZN(W12045));
  NANDX1 G32202 (.A1(W14095), .A2(W20830), .ZN(W21296));
  NANDX1 G32203 (.A1(W4886), .A2(W1768), .ZN(W12044));
  NANDX1 G32204 (.A1(W1616), .A2(I1236), .ZN(W2766));
  NANDX1 G32205 (.A1(I468), .A2(W9161), .ZN(W21300));
  NANDX1 G32206 (.A1(W10881), .A2(W13691), .ZN(W21301));
  NANDX1 G32207 (.A1(W20967), .A2(W11711), .ZN(O2206));
  NANDX1 G32208 (.A1(W1334), .A2(W1875), .ZN(W25124));
  NANDX1 G32209 (.A1(W5552), .A2(W3585), .ZN(W12043));
  NANDX1 G32210 (.A1(W2643), .A2(I1762), .ZN(W2779));
  NANDX1 G32211 (.A1(I22), .A2(I670), .ZN(W12066));
  NANDX1 G32212 (.A1(I228), .A2(I229), .ZN(W114));
  NANDX1 G32213 (.A1(I499), .A2(W7378), .ZN(W8930));
  NANDX1 G32214 (.A1(I232), .A2(I233), .ZN(W116));
  NANDX1 G32215 (.A1(W4562), .A2(W13556), .ZN(W21254));
  NANDX1 G32216 (.A1(I1293), .A2(I526), .ZN(W8931));
  NANDX1 G32217 (.A1(W8254), .A2(W5475), .ZN(W10281));
  NANDX1 G32218 (.A1(W14365), .A2(W11855), .ZN(W25145));
  NANDX1 G32219 (.A1(W2021), .A2(W4732), .ZN(W21255));
  NANDX1 G32220 (.A1(I643), .A2(W1897), .ZN(W2782));
  NANDX1 G32221 (.A1(W10477), .A2(I948), .ZN(W12062));
  NANDX1 G32222 (.A1(W20712), .A2(W1088), .ZN(W25144));
  NANDX1 G32223 (.A1(W2750), .A2(W2636), .ZN(W2780));
  NANDX1 G32224 (.A1(W15019), .A2(W20668), .ZN(W21257));
  NANDX1 G32225 (.A1(W11165), .A2(I555), .ZN(W11991));
  NANDX1 G32226 (.A1(I236), .A2(I237), .ZN(W118));
  NANDX1 G32227 (.A1(I238), .A2(I239), .ZN(W119));
  NANDX1 G32228 (.A1(W1295), .A2(W9765), .ZN(O2194));
  NANDX1 G32229 (.A1(W960), .A2(W8395), .ZN(W21259));
  NANDX1 G32230 (.A1(I463), .A2(W5372), .ZN(W8934));
  NANDX1 G32231 (.A1(W10268), .A2(W6988), .ZN(W12059));
  NANDX1 G32232 (.A1(W2957), .A2(W7978), .ZN(W21268));
  NANDX1 G32233 (.A1(W953), .A2(W18693), .ZN(W21270));
  NANDX1 G32234 (.A1(W24927), .A2(W10807), .ZN(W25138));
  NANDX1 G32235 (.A1(I702), .A2(W2116), .ZN(W2776));
  NANDX1 G32236 (.A1(W9541), .A2(W5350), .ZN(O2197));
  NANDX1 G32237 (.A1(W3537), .A2(W8050), .ZN(W8937));
  NANDX1 G32238 (.A1(W7772), .A2(W5370), .ZN(W10282));
  NANDX1 G32239 (.A1(I242), .A2(I243), .ZN(W121));
  NANDX1 G32240 (.A1(W12150), .A2(W4486), .ZN(W21589));
  NANDX1 G32241 (.A1(I1324), .A2(W1324), .ZN(W2562));
  NANDX1 G32242 (.A1(W2362), .A2(W6398), .ZN(W21575));
  NANDX1 G32243 (.A1(I390), .A2(I391), .ZN(W195));
  NANDX1 G32244 (.A1(I725), .A2(W925), .ZN(W2561));
  NANDX1 G32245 (.A1(W103), .A2(W6600), .ZN(W21579));
  NANDX1 G32246 (.A1(W20086), .A2(W3820), .ZN(W21580));
  NANDX1 G32247 (.A1(I191), .A2(W5799), .ZN(W10340));
  NANDX1 G32248 (.A1(W5079), .A2(W6683), .ZN(W25025));
  NANDX1 G32249 (.A1(W6123), .A2(I1244), .ZN(W10086));
  NANDX1 G32250 (.A1(I858), .A2(I1719), .ZN(W11933));
  NANDX1 G32251 (.A1(W6837), .A2(W2429), .ZN(W25024));
  NANDX1 G32252 (.A1(W393), .A2(W2788), .ZN(W9046));
  NANDX1 G32253 (.A1(I392), .A2(I393), .ZN(W196));
  NANDX1 G32254 (.A1(W4379), .A2(W7251), .ZN(W11932));
  NANDX1 G32255 (.A1(W3114), .A2(W2811), .ZN(W21587));
  NANDX1 G32256 (.A1(I1652), .A2(W9742), .ZN(O2283));
  NANDX1 G32257 (.A1(W19391), .A2(W11737), .ZN(W21590));
  NANDX1 G32258 (.A1(W13753), .A2(W12960), .ZN(O3270));
  NANDX1 G32259 (.A1(I176), .A2(W2127), .ZN(W2554));
  NANDX1 G32260 (.A1(W195), .A2(W385), .ZN(W2552));
  NANDX1 G32261 (.A1(I32), .A2(W1495), .ZN(W2549));
  NANDX1 G32262 (.A1(W13747), .A2(W10405), .ZN(O3268));
  NANDX1 G32263 (.A1(W4494), .A2(W7040), .ZN(W9054));
  NANDX1 G32264 (.A1(W3554), .A2(W2005), .ZN(W10347));
  NANDX1 G32265 (.A1(W19526), .A2(W3030), .ZN(W21600));
  NANDX1 G32266 (.A1(W5053), .A2(W4842), .ZN(W9055));
  NANDX1 G32267 (.A1(W3790), .A2(W20275), .ZN(W21601));
  NANDX1 G32268 (.A1(I313), .A2(W1769), .ZN(W2547));
  NANDX1 G32269 (.A1(W8158), .A2(W15616), .ZN(W21605));
  NANDX1 G32270 (.A1(W8290), .A2(W2431), .ZN(W10082));
  NANDX1 G32271 (.A1(I296), .A2(I85), .ZN(W2574));
  NANDX1 G32272 (.A1(W15179), .A2(W4604), .ZN(W21544));
  NANDX1 G32273 (.A1(W3888), .A2(W10594), .ZN(W21545));
  NANDX1 G32274 (.A1(W100), .A2(W6277), .ZN(W10090));
  NANDX1 G32275 (.A1(W9592), .A2(I1894), .ZN(W10332));
  NANDX1 G32276 (.A1(W4067), .A2(W8323), .ZN(W10087));
  NANDX1 G32277 (.A1(W11249), .A2(W2673), .ZN(O551));
  NANDX1 G32278 (.A1(W258), .A2(W16554), .ZN(O3273));
  NANDX1 G32279 (.A1(W2528), .A2(W6654), .ZN(W11942));
  NANDX1 G32280 (.A1(W9102), .A2(W7578), .ZN(W11941));
  NANDX1 G32281 (.A1(W24931), .A2(W19102), .ZN(W25034));
  NANDX1 G32282 (.A1(I1394), .A2(W16988), .ZN(W25033));
  NANDX1 G32283 (.A1(W1832), .A2(I1148), .ZN(W2576));
  NANDX1 G32284 (.A1(I109), .A2(W545), .ZN(W2575));
  NANDX1 G32285 (.A1(W12384), .A2(W16875), .ZN(W21551));
  NANDX1 G32286 (.A1(W6710), .A2(W6172), .ZN(W11923));
  NANDX1 G32287 (.A1(W1717), .A2(W397), .ZN(W2573));
  NANDX1 G32288 (.A1(W534), .A2(W863), .ZN(W2572));
  NANDX1 G32289 (.A1(W1299), .A2(W1824), .ZN(W2571));
  NANDX1 G32290 (.A1(I386), .A2(I387), .ZN(W193));
  NANDX1 G32291 (.A1(W2937), .A2(W2765), .ZN(W9040));
  NANDX1 G32292 (.A1(W1612), .A2(W867), .ZN(W2569));
  NANDX1 G32293 (.A1(I388), .A2(I389), .ZN(W194));
  NANDX1 G32294 (.A1(W2653), .A2(W5874), .ZN(W9042));
  NANDX1 G32295 (.A1(W2291), .A2(W3248), .ZN(W11936));
  NANDX1 G32296 (.A1(W21301), .A2(W6857), .ZN(W25029));
  NANDX1 G32297 (.A1(W5868), .A2(W4525), .ZN(W9044));
  NANDX1 G32298 (.A1(W11122), .A2(W18654), .ZN(O2281));
  NANDX1 G32299 (.A1(W3808), .A2(W300), .ZN(W25027));
  NANDX1 G32300 (.A1(I521), .A2(W6636), .ZN(O2282));
  NANDX1 G32301 (.A1(W2128), .A2(W21143), .ZN(W21654));
  NANDX1 G32302 (.A1(W10014), .A2(I0), .ZN(W11915));
  NANDX1 G32303 (.A1(I392), .A2(W620), .ZN(W2532));
  NANDX1 G32304 (.A1(W2403), .A2(W2347), .ZN(W2531));
  NANDX1 G32305 (.A1(I432), .A2(I433), .ZN(W216));
  NANDX1 G32306 (.A1(W19133), .A2(W7955), .ZN(W25007));
  NANDX1 G32307 (.A1(I436), .A2(I437), .ZN(W218));
  NANDX1 G32308 (.A1(W5688), .A2(W5685), .ZN(W11914));
  NANDX1 G32309 (.A1(I1148), .A2(I1516), .ZN(W2526));
  NANDX1 G32310 (.A1(W410), .A2(W6869), .ZN(W10359));
  NANDX1 G32311 (.A1(W14109), .A2(W8129), .ZN(W25006));
  NANDX1 G32312 (.A1(W110), .A2(W2295), .ZN(W9067));
  NANDX1 G32313 (.A1(W1686), .A2(I450), .ZN(W2524));
  NANDX1 G32314 (.A1(I309), .A2(W3259), .ZN(W21651));
  NANDX1 G32315 (.A1(W1017), .A2(W2366), .ZN(W2523));
  NANDX1 G32316 (.A1(W3223), .A2(W4678), .ZN(W11911));
  NANDX1 G32317 (.A1(W11171), .A2(W10151), .ZN(W21644));
  NANDX1 G32318 (.A1(W2413), .A2(W2531), .ZN(W9068));
  NANDX1 G32319 (.A1(I438), .A2(I439), .ZN(W219));
  NANDX1 G32320 (.A1(W4430), .A2(W8682), .ZN(W10361));
  NANDX1 G32321 (.A1(W2210), .A2(W11039), .ZN(W11909));
  NANDX1 G32322 (.A1(W1929), .A2(W6493), .ZN(W11907));
  NANDX1 G32323 (.A1(W8222), .A2(W4587), .ZN(W21660));
  NANDX1 G32324 (.A1(W16477), .A2(W7194), .ZN(W25003));
  NANDX1 G32325 (.A1(W14726), .A2(W2121), .ZN(W21662));
  NANDX1 G32326 (.A1(I1392), .A2(I682), .ZN(W2516));
  NANDX1 G32327 (.A1(W341), .A2(W1152), .ZN(W2515));
  NANDX1 G32328 (.A1(W6981), .A2(W10499), .ZN(O546));
  NANDX1 G32329 (.A1(W17746), .A2(W7731), .ZN(W21667));
  NANDX1 G32330 (.A1(W13135), .A2(W15272), .ZN(O3266));
  NANDX1 G32331 (.A1(W11027), .A2(W10950), .ZN(O2305));
  NANDX1 G32332 (.A1(I422), .A2(I423), .ZN(W211));
  NANDX1 G32333 (.A1(W1236), .A2(W2064), .ZN(W2542));
  NANDX1 G32334 (.A1(W8600), .A2(W14335), .ZN(W21610));
  NANDX1 G32335 (.A1(W5676), .A2(W1034), .ZN(W11922));
  NANDX1 G32336 (.A1(W15465), .A2(W16215), .ZN(W21612));
  NANDX1 G32337 (.A1(I1055), .A2(W1151), .ZN(W2541));
  NANDX1 G32338 (.A1(W8601), .A2(W4097), .ZN(W10348));
  NANDX1 G32339 (.A1(W5785), .A2(I1799), .ZN(W11920));
  NANDX1 G32340 (.A1(W15632), .A2(W20584), .ZN(W21615));
  NANDX1 G32341 (.A1(W5456), .A2(W19447), .ZN(W21617));
  NANDX1 G32342 (.A1(I404), .A2(I405), .ZN(W202));
  NANDX1 G32343 (.A1(W1662), .A2(W17992), .ZN(W21624));
  NANDX1 G32344 (.A1(I408), .A2(I409), .ZN(W204));
  NANDX1 G32345 (.A1(W8770), .A2(W942), .ZN(W10349));
  NANDX1 G32346 (.A1(I1053), .A2(I272), .ZN(W2538));
  NANDX1 G32347 (.A1(I1546), .A2(W7169), .ZN(W10091));
  NANDX1 G32348 (.A1(I1158), .A2(W9469), .ZN(W10352));
  NANDX1 G32349 (.A1(I1976), .A2(W6974), .ZN(W11918));
  NANDX1 G32350 (.A1(W3836), .A2(W12387), .ZN(W21632));
  NANDX1 G32351 (.A1(I1994), .A2(W5283), .ZN(O2299));
  NANDX1 G32352 (.A1(W15191), .A2(W1346), .ZN(W25010));
  NANDX1 G32353 (.A1(I983), .A2(I582), .ZN(W2536));
  NANDX1 G32354 (.A1(I832), .A2(I1919), .ZN(W2535));
  NANDX1 G32355 (.A1(I428), .A2(I429), .ZN(W214));
  NANDX1 G32356 (.A1(W13370), .A2(W423), .ZN(W21637));
  NANDX1 G32357 (.A1(W6200), .A2(W14418), .ZN(W21638));
  NANDX1 G32358 (.A1(W5013), .A2(W874), .ZN(W9064));
  NANDX1 G32359 (.A1(I1367), .A2(W2960), .ZN(W11916));
  NANDX1 G32360 (.A1(W3980), .A2(W3563), .ZN(W10357));
  NANDX1 G32361 (.A1(W1602), .A2(I1392), .ZN(W2533));
  NANDX1 G32362 (.A1(W20232), .A2(W6671), .ZN(W25063));
  NANDX1 G32363 (.A1(I350), .A2(I351), .ZN(W175));
  NANDX1 G32364 (.A1(W2795), .A2(W8124), .ZN(W11977));
  NANDX1 G32365 (.A1(W6705), .A2(W45), .ZN(W25064));
  NANDX1 G32366 (.A1(W475), .A2(I960), .ZN(W2658));
  NANDX1 G32367 (.A1(W476), .A2(W1942), .ZN(W2656));
  NANDX1 G32368 (.A1(W9065), .A2(W33), .ZN(O2250));
  NANDX1 G32369 (.A1(W14976), .A2(W7987), .ZN(W21466));
  NANDX1 G32370 (.A1(W16053), .A2(W19916), .ZN(W21467));
  NANDX1 G32371 (.A1(W3463), .A2(W6730), .ZN(W21468));
  NANDX1 G32372 (.A1(W8993), .A2(W9359), .ZN(W21469));
  NANDX1 G32373 (.A1(I1111), .A2(W1687), .ZN(W9007));
  NANDX1 G32374 (.A1(W10537), .A2(W2746), .ZN(W11974));
  NANDX1 G32375 (.A1(I564), .A2(I1976), .ZN(W2650));
  NANDX1 G32376 (.A1(I352), .A2(I353), .ZN(W176));
  NANDX1 G32377 (.A1(I1322), .A2(I194), .ZN(W2649));
  NANDX1 G32378 (.A1(W1774), .A2(W2237), .ZN(W2660));
  NANDX1 G32379 (.A1(W2800), .A2(W23490), .ZN(O3284));
  NANDX1 G32380 (.A1(W141), .A2(W1561), .ZN(W2643));
  NANDX1 G32381 (.A1(I354), .A2(I355), .ZN(W177));
  NANDX1 G32382 (.A1(I974), .A2(I1864), .ZN(W2640));
  NANDX1 G32383 (.A1(W6920), .A2(W8556), .ZN(W10098));
  NANDX1 G32384 (.A1(W1519), .A2(I1465), .ZN(W2639));
  NANDX1 G32385 (.A1(W6944), .A2(W3879), .ZN(W9011));
  NANDX1 G32386 (.A1(I356), .A2(I357), .ZN(W178));
  NANDX1 G32387 (.A1(W1475), .A2(W458), .ZN(W2637));
  NANDX1 G32388 (.A1(W6085), .A2(W9566), .ZN(O554));
  NANDX1 G32389 (.A1(W16622), .A2(W9435), .ZN(W25056));
  NANDX1 G32390 (.A1(W6131), .A2(W4905), .ZN(W10097));
  NANDX1 G32391 (.A1(I360), .A2(I361), .ZN(W180));
  NANDX1 G32392 (.A1(W23848), .A2(W17059), .ZN(W25053));
  NANDX1 G32393 (.A1(I1602), .A2(W2405), .ZN(W2668));
  NANDX1 G32394 (.A1(I322), .A2(I323), .ZN(W161));
  NANDX1 G32395 (.A1(I1594), .A2(W2175), .ZN(W2676));
  NANDX1 G32396 (.A1(W828), .A2(W7343), .ZN(W8996));
  NANDX1 G32397 (.A1(W17021), .A2(W20908), .ZN(W21436));
  NANDX1 G32398 (.A1(W23399), .A2(W17574), .ZN(W25076));
  NANDX1 G32399 (.A1(I328), .A2(I329), .ZN(W164));
  NANDX1 G32400 (.A1(I1962), .A2(W5277), .ZN(W11988));
  NANDX1 G32401 (.A1(W4579), .A2(I306), .ZN(W11986));
  NANDX1 G32402 (.A1(W1458), .A2(W5340), .ZN(W10105));
  NANDX1 G32403 (.A1(I447), .A2(W2085), .ZN(W2670));
  NANDX1 G32404 (.A1(W8334), .A2(W5978), .ZN(W11985));
  NANDX1 G32405 (.A1(W17819), .A2(W7116), .ZN(O2246));
  NANDX1 G32406 (.A1(W10030), .A2(W3164), .ZN(W10101));
  NANDX1 G32407 (.A1(I382), .A2(W1605), .ZN(W8999));
  NANDX1 G32408 (.A1(W1802), .A2(W3503), .ZN(W11964));
  NANDX1 G32409 (.A1(W143), .A2(W3491), .ZN(W9002));
  NANDX1 G32410 (.A1(W539), .A2(W1661), .ZN(W2666));
  NANDX1 G32411 (.A1(I348), .A2(I349), .ZN(W174));
  NANDX1 G32412 (.A1(W612), .A2(W1205), .ZN(W2663));
  NANDX1 G32413 (.A1(W16853), .A2(W22956), .ZN(O3285));
  NANDX1 G32414 (.A1(W6630), .A2(W10176), .ZN(W10318));
  NANDX1 G32415 (.A1(I1439), .A2(I1128), .ZN(W21454));
  NANDX1 G32416 (.A1(W9832), .A2(W4531), .ZN(W21455));
  NANDX1 G32417 (.A1(W530), .A2(I1208), .ZN(W2662));
  NANDX1 G32418 (.A1(W21414), .A2(W7431), .ZN(W25065));
  NANDX1 G32419 (.A1(I838), .A2(I1547), .ZN(W9004));
  NANDX1 G32420 (.A1(W6518), .A2(W2957), .ZN(W10099));
  NANDX1 G32421 (.A1(W9028), .A2(W19301), .ZN(W21459));
  NANDX1 G32422 (.A1(W1772), .A2(W5170), .ZN(W9005));
  NANDX1 G32423 (.A1(W11230), .A2(W6598), .ZN(W21524));
  NANDX1 G32424 (.A1(W8105), .A2(W5339), .ZN(W9025));
  NANDX1 G32425 (.A1(W6238), .A2(W8494), .ZN(W9026));
  NANDX1 G32426 (.A1(W565), .A2(W8174), .ZN(W11953));
  NANDX1 G32427 (.A1(I370), .A2(I371), .ZN(W185));
  NANDX1 G32428 (.A1(I918), .A2(I1214), .ZN(W2602));
  NANDX1 G32429 (.A1(W96), .A2(W20060), .ZN(W21519));
  NANDX1 G32430 (.A1(W9178), .A2(W9679), .ZN(W11952));
  NANDX1 G32431 (.A1(W173), .A2(I884), .ZN(W2599));
  NANDX1 G32432 (.A1(W442), .A2(W1838), .ZN(W2598));
  NANDX1 G32433 (.A1(W4735), .A2(W13524), .ZN(O3275));
  NANDX1 G32434 (.A1(W17198), .A2(I905), .ZN(W25038));
  NANDX1 G32435 (.A1(I104), .A2(W1196), .ZN(W2597));
  NANDX1 G32436 (.A1(W20722), .A2(W11986), .ZN(W21521));
  NANDX1 G32437 (.A1(W2936), .A2(W6262), .ZN(W11951));
  NANDX1 G32438 (.A1(W1488), .A2(W1284), .ZN(W2613));
  NANDX1 G32439 (.A1(W5333), .A2(W9782), .ZN(W11950));
  NANDX1 G32440 (.A1(W957), .A2(I1314), .ZN(W2591));
  NANDX1 G32441 (.A1(W3548), .A2(W2601), .ZN(W9027));
  NANDX1 G32442 (.A1(W5864), .A2(W380), .ZN(W9028));
  NANDX1 G32443 (.A1(W19064), .A2(W21037), .ZN(W21534));
  NANDX1 G32444 (.A1(W6909), .A2(W8462), .ZN(W9029));
  NANDX1 G32445 (.A1(W17996), .A2(W17621), .ZN(O2273));
  NANDX1 G32446 (.A1(W1417), .A2(I1862), .ZN(W11945));
  NANDX1 G32447 (.A1(W246), .A2(W634), .ZN(W2586));
  NANDX1 G32448 (.A1(W2435), .A2(W8562), .ZN(W11944));
  NANDX1 G32449 (.A1(W16141), .A2(W3602), .ZN(W21541));
  NANDX1 G32450 (.A1(W21442), .A2(W1278), .ZN(W21542));
  NANDX1 G32451 (.A1(W10426), .A2(W7120), .ZN(W21543));
  NANDX1 G32452 (.A1(W2283), .A2(W840), .ZN(W2584));
  NANDX1 G32453 (.A1(W3183), .A2(W5731), .ZN(W11957));
  NANDX1 G32454 (.A1(W8177), .A2(W5205), .ZN(W21487));
  NANDX1 G32455 (.A1(W2307), .A2(W1400), .ZN(W2631));
  NANDX1 G32456 (.A1(W7404), .A2(I530), .ZN(O3279));
  NANDX1 G32457 (.A1(I1950), .A2(I1554), .ZN(W2630));
  NANDX1 G32458 (.A1(W835), .A2(W1359), .ZN(O362));
  NANDX1 G32459 (.A1(I498), .A2(W884), .ZN(W2629));
  NANDX1 G32460 (.A1(W674), .A2(W1621), .ZN(W2628));
  NANDX1 G32461 (.A1(W2274), .A2(W2173), .ZN(W2625));
  NANDX1 G32462 (.A1(W1970), .A2(W1862), .ZN(W2623));
  NANDX1 G32463 (.A1(W1744), .A2(W377), .ZN(W2622));
  NANDX1 G32464 (.A1(W11071), .A2(W13365), .ZN(W21494));
  NANDX1 G32465 (.A1(W2340), .A2(W258), .ZN(W11958));
  NANDX1 G32466 (.A1(W351), .A2(W206), .ZN(W2619));
  NANDX1 G32467 (.A1(W6633), .A2(W10522), .ZN(O2260));
  NANDX1 G32468 (.A1(W8535), .A2(W2249), .ZN(W12088));
  NANDX1 G32469 (.A1(W230), .A2(W2560), .ZN(W2618));
  NANDX1 G32470 (.A1(W19461), .A2(W557), .ZN(O2263));
  NANDX1 G32471 (.A1(W17947), .A2(W18000), .ZN(W25044));
  NANDX1 G32472 (.A1(W14125), .A2(W16846), .ZN(W21504));
  NANDX1 G32473 (.A1(I584), .A2(W609), .ZN(W2616));
  NANDX1 G32474 (.A1(W6443), .A2(W20643), .ZN(O2264));
  NANDX1 G32475 (.A1(W5321), .A2(W3504), .ZN(W11956));
  NANDX1 G32476 (.A1(W18586), .A2(W16141), .ZN(W21509));
  NANDX1 G32477 (.A1(W17074), .A2(W1508), .ZN(W25041));
  NANDX1 G32478 (.A1(W8213), .A2(W1197), .ZN(W9024));
  NANDX1 G32479 (.A1(W14874), .A2(W13345), .ZN(W21511));
  NANDX1 G32480 (.A1(I1814), .A2(I1346), .ZN(W2614));
  NANDX1 G32481 (.A1(W19520), .A2(W18801), .ZN(W25040));
  NANDX1 G32482 (.A1(W3509), .A2(I770), .ZN(O2266));
  NANDX1 G32483 (.A1(W3197), .A2(W18933), .ZN(W20885));
  NANDX1 G32484 (.A1(W18589), .A2(W17810), .ZN(W25272));
  NANDX1 G32485 (.A1(W5586), .A2(W9215), .ZN(W20874));
  NANDX1 G32486 (.A1(W2972), .A2(W14546), .ZN(W20876));
  NANDX1 G32487 (.A1(W3013), .A2(I595), .ZN(W3034));
  NANDX1 G32488 (.A1(W15688), .A2(W7473), .ZN(W20878));
  NANDX1 G32489 (.A1(W3153), .A2(W1858), .ZN(W8823));
  NANDX1 G32490 (.A1(W9705), .A2(W12236), .ZN(W20881));
  NANDX1 G32491 (.A1(W22977), .A2(W1655), .ZN(W25270));
  NANDX1 G32492 (.A1(W479), .A2(W2612), .ZN(W10170));
  NANDX1 G32493 (.A1(W1037), .A2(W10565), .ZN(W12239));
  NANDX1 G32494 (.A1(W2273), .A2(W5264), .ZN(W10169));
  NANDX1 G32495 (.A1(W3575), .A2(W10800), .ZN(W20883));
  NANDX1 G32496 (.A1(W1296), .A2(W2093), .ZN(O3350));
  NANDX1 G32497 (.A1(W2730), .A2(W15372), .ZN(W20884));
  NANDX1 G32498 (.A1(W1137), .A2(W9199), .ZN(W25266));
  NANDX1 G32499 (.A1(W176), .A2(W2421), .ZN(W8818));
  NANDX1 G32500 (.A1(W1190), .A2(W2928), .ZN(W3032));
  NANDX1 G32501 (.A1(W15722), .A2(W18435), .ZN(W20887));
  NANDX1 G32502 (.A1(W3391), .A2(W8079), .ZN(W20888));
  NANDX1 G32503 (.A1(W3250), .A2(W2489), .ZN(O369));
  NANDX1 G32504 (.A1(W17165), .A2(W10952), .ZN(W20889));
  NANDX1 G32505 (.A1(W11981), .A2(W10520), .ZN(W20892));
  NANDX1 G32506 (.A1(I1050), .A2(I1193), .ZN(W8825));
  NANDX1 G32507 (.A1(I84), .A2(I85), .ZN(W42));
  NANDX1 G32508 (.A1(I352), .A2(W10190), .ZN(O2106));
  NANDX1 G32509 (.A1(W184), .A2(W1375), .ZN(W3024));
  NANDX1 G32510 (.A1(W19969), .A2(W822), .ZN(W20895));
  NANDX1 G32511 (.A1(W6123), .A2(W2655), .ZN(W20896));
  NANDX1 G32512 (.A1(W3156), .A2(W1612), .ZN(W8828));
  NANDX1 G32513 (.A1(I380), .A2(W437), .ZN(W3023));
  NANDX1 G32514 (.A1(W1179), .A2(I798), .ZN(W3055));
  NANDX1 G32515 (.A1(W3189), .A2(W6631), .ZN(W8812));
  NANDX1 G32516 (.A1(I875), .A2(W16337), .ZN(W25290));
  NANDX1 G32517 (.A1(W1341), .A2(I421), .ZN(W3062));
  NANDX1 G32518 (.A1(W12872), .A2(W3641), .ZN(O3360));
  NANDX1 G32519 (.A1(W14579), .A2(W7625), .ZN(W20854));
  NANDX1 G32520 (.A1(W8013), .A2(I1091), .ZN(W10209));
  NANDX1 G32521 (.A1(I54), .A2(I55), .ZN(W27));
  NANDX1 G32522 (.A1(I60), .A2(I61), .ZN(W30));
  NANDX1 G32523 (.A1(W5903), .A2(W6231), .ZN(W10177));
  NANDX1 G32524 (.A1(W18352), .A2(W22729), .ZN(W25283));
  NANDX1 G32525 (.A1(W2209), .A2(I1894), .ZN(W3058));
  NANDX1 G32526 (.A1(W18022), .A2(W13345), .ZN(W20859));
  NANDX1 G32527 (.A1(W2808), .A2(W2635), .ZN(W12248));
  NANDX1 G32528 (.A1(I576), .A2(W8067), .ZN(W12247));
  NANDX1 G32529 (.A1(W3645), .A2(W4787), .ZN(W12235));
  NANDX1 G32530 (.A1(W2508), .A2(W2164), .ZN(O28));
  NANDX1 G32531 (.A1(W9660), .A2(W12135), .ZN(W12246));
  NANDX1 G32532 (.A1(W11131), .A2(W11617), .ZN(W12244));
  NANDX1 G32533 (.A1(W2518), .A2(W2024), .ZN(W3050));
  NANDX1 G32534 (.A1(I1486), .A2(W2834), .ZN(W3049));
  NANDX1 G32535 (.A1(I246), .A2(I123), .ZN(W3048));
  NANDX1 G32536 (.A1(W8417), .A2(W7491), .ZN(W10175));
  NANDX1 G32537 (.A1(I1467), .A2(W6516), .ZN(W10173));
  NANDX1 G32538 (.A1(W5709), .A2(W10425), .ZN(W12242));
  NANDX1 G32539 (.A1(W6665), .A2(W18226), .ZN(W20869));
  NANDX1 G32540 (.A1(W1537), .A2(W1806), .ZN(W3044));
  NANDX1 G32541 (.A1(W8041), .A2(W6125), .ZN(W10212));
  NANDX1 G32542 (.A1(W6985), .A2(W3875), .ZN(W20870));
  NANDX1 G32543 (.A1(W2240), .A2(I1321), .ZN(W3042));
  NANDX1 G32544 (.A1(I102), .A2(I103), .ZN(W51));
  NANDX1 G32545 (.A1(W4188), .A2(W17897), .ZN(O2110));
  NANDX1 G32546 (.A1(W12824), .A2(W2980), .ZN(W20928));
  NANDX1 G32547 (.A1(W8693), .A2(W19301), .ZN(O2111));
  NANDX1 G32548 (.A1(I1651), .A2(W902), .ZN(W2994));
  NANDX1 G32549 (.A1(W1744), .A2(I1108), .ZN(W2993));
  NANDX1 G32550 (.A1(I737), .A2(W470), .ZN(W2992));
  NANDX1 G32551 (.A1(W4275), .A2(W15746), .ZN(W20931));
  NANDX1 G32552 (.A1(W2320), .A2(W15644), .ZN(W25255));
  NANDX1 G32553 (.A1(W5657), .A2(W8100), .ZN(W12222));
  NANDX1 G32554 (.A1(W2548), .A2(W2795), .ZN(W10230));
  NANDX1 G32555 (.A1(W13872), .A2(W10198), .ZN(W20936));
  NANDX1 G32556 (.A1(W793), .A2(W14826), .ZN(O2115));
  NANDX1 G32557 (.A1(W803), .A2(W6194), .ZN(W20938));
  NANDX1 G32558 (.A1(W20312), .A2(W7084), .ZN(W20939));
  NANDX1 G32559 (.A1(I872), .A2(W2129), .ZN(W2988));
  NANDX1 G32560 (.A1(W7377), .A2(W288), .ZN(W8836));
  NANDX1 G32561 (.A1(W8471), .A2(W5469), .ZN(W8844));
  NANDX1 G32562 (.A1(I1794), .A2(W944), .ZN(W2987));
  NANDX1 G32563 (.A1(W854), .A2(I1210), .ZN(W2982));
  NANDX1 G32564 (.A1(W10942), .A2(W15439), .ZN(W20940));
  NANDX1 G32565 (.A1(W5907), .A2(W5225), .ZN(O2116));
  NANDX1 G32566 (.A1(W1374), .A2(W8016), .ZN(W12221));
  NANDX1 G32567 (.A1(W14954), .A2(W18845), .ZN(O2117));
  NANDX1 G32568 (.A1(W1409), .A2(I958), .ZN(W2978));
  NANDX1 G32569 (.A1(W6038), .A2(W155), .ZN(W12219));
  NANDX1 G32570 (.A1(W593), .A2(W11242), .ZN(W12216));
  NANDX1 G32571 (.A1(W1170), .A2(I1447), .ZN(W2973));
  NANDX1 G32572 (.A1(W10533), .A2(W10254), .ZN(O2119));
  NANDX1 G32573 (.A1(W18000), .A2(W1234), .ZN(W20951));
  NANDX1 G32574 (.A1(W7610), .A2(W5), .ZN(W12212));
  NANDX1 G32575 (.A1(I94), .A2(I95), .ZN(W47));
  NANDX1 G32576 (.A1(W11083), .A2(W105), .ZN(W20900));
  NANDX1 G32577 (.A1(W8316), .A2(W869), .ZN(W10221));
  NANDX1 G32578 (.A1(W8820), .A2(W7231), .ZN(W8831));
  NANDX1 G32579 (.A1(W5983), .A2(W7235), .ZN(W12230));
  NANDX1 G32580 (.A1(W220), .A2(W751), .ZN(W3018));
  NANDX1 G32581 (.A1(W2433), .A2(W992), .ZN(W3017));
  NANDX1 G32582 (.A1(W3844), .A2(W9354), .ZN(W20905));
  NANDX1 G32583 (.A1(W923), .A2(W739), .ZN(W3016));
  NANDX1 G32584 (.A1(W9503), .A2(W9753), .ZN(W10226));
  NANDX1 G32585 (.A1(W5307), .A2(W5116), .ZN(W20910));
  NANDX1 G32586 (.A1(W13477), .A2(W7283), .ZN(W20911));
  NANDX1 G32587 (.A1(W2271), .A2(W2313), .ZN(W3015));
  NANDX1 G32588 (.A1(W1252), .A2(W1534), .ZN(W3012));
  NANDX1 G32589 (.A1(I1163), .A2(W1600), .ZN(W3010));
  NANDX1 G32590 (.A1(W7179), .A2(W2450), .ZN(W8810));
  NANDX1 G32591 (.A1(W2522), .A2(W1388), .ZN(W3008));
  NANDX1 G32592 (.A1(I1236), .A2(W888), .ZN(W3006));
  NANDX1 G32593 (.A1(W1146), .A2(W1379), .ZN(W10167));
  NANDX1 G32594 (.A1(W5592), .A2(W1361), .ZN(O581));
  NANDX1 G32595 (.A1(W369), .A2(W8196), .ZN(W20916));
  NANDX1 G32596 (.A1(W8231), .A2(W11060), .ZN(W12226));
  NANDX1 G32597 (.A1(W10273), .A2(W19324), .ZN(O2109));
  NANDX1 G32598 (.A1(W20269), .A2(W8181), .ZN(W20923));
  NANDX1 G32599 (.A1(W9787), .A2(W2575), .ZN(W12225));
  NANDX1 G32600 (.A1(I422), .A2(W18731), .ZN(O3346));
  NANDX1 G32601 (.A1(W10087), .A2(W14817), .ZN(W25256));
  NANDX1 G32602 (.A1(W1588), .A2(W6832), .ZN(W8834));
  NANDX1 G32603 (.A1(W7299), .A2(W8672), .ZN(W10166));
  NANDX1 G32604 (.A1(I1044), .A2(W9841), .ZN(O580));
  NANDX1 G32605 (.A1(W1029), .A2(I1042), .ZN(W3103));
  NANDX1 G32606 (.A1(W20287), .A2(I444), .ZN(W20777));
  NANDX1 G32607 (.A1(W906), .A2(W767), .ZN(W3113));
  NANDX1 G32608 (.A1(I16), .A2(I17), .ZN(W8));
  NANDX1 G32609 (.A1(W12865), .A2(W5477), .ZN(O3378));
  NANDX1 G32610 (.A1(W8440), .A2(W1280), .ZN(W12282));
  NANDX1 G32611 (.A1(W55), .A2(I1466), .ZN(W3111));
  NANDX1 G32612 (.A1(W12751), .A2(W10107), .ZN(W20779));
  NANDX1 G32613 (.A1(W7391), .A2(W7052), .ZN(W12281));
  NANDX1 G32614 (.A1(I18), .A2(I19), .ZN(W9));
  NANDX1 G32615 (.A1(I22), .A2(I23), .ZN(W11));
  NANDX1 G32616 (.A1(W7133), .A2(W2557), .ZN(O2081));
  NANDX1 G32617 (.A1(W9251), .A2(W8165), .ZN(W12280));
  NANDX1 G32618 (.A1(W5949), .A2(W3181), .ZN(W8795));
  NANDX1 G32619 (.A1(W2449), .A2(W2479), .ZN(W3105));
  NANDX1 G32620 (.A1(W2462), .A2(W6362), .ZN(W8796));
  NANDX1 G32621 (.A1(W8557), .A2(W1568), .ZN(W8790));
  NANDX1 G32622 (.A1(W6834), .A2(W9725), .ZN(O589));
  NANDX1 G32623 (.A1(W3157), .A2(W4339), .ZN(O247));
  NANDX1 G32624 (.A1(W2407), .A2(W8983), .ZN(W12278));
  NANDX1 G32625 (.A1(W4478), .A2(W1365), .ZN(W10183));
  NANDX1 G32626 (.A1(W1754), .A2(W171), .ZN(W3100));
  NANDX1 G32627 (.A1(W1019), .A2(W125), .ZN(W3099));
  NANDX1 G32628 (.A1(W1875), .A2(I681), .ZN(W12275));
  NANDX1 G32629 (.A1(W17993), .A2(W12207), .ZN(W25328));
  NANDX1 G32630 (.A1(I28), .A2(I29), .ZN(W14));
  NANDX1 G32631 (.A1(I748), .A2(W8289), .ZN(W10197));
  NANDX1 G32632 (.A1(W18572), .A2(W13698), .ZN(W25327));
  NANDX1 G32633 (.A1(W2216), .A2(W445), .ZN(W3095));
  NANDX1 G32634 (.A1(I980), .A2(I756), .ZN(O29));
  NANDX1 G32635 (.A1(W10098), .A2(W1347), .ZN(W10182));
  NANDX1 G32636 (.A1(I601), .A2(W20060), .ZN(W25337));
  NANDX1 G32637 (.A1(W16346), .A2(W14261), .ZN(O2073));
  NANDX1 G32638 (.A1(W1614), .A2(W7724), .ZN(W20755));
  NANDX1 G32639 (.A1(W11580), .A2(W11698), .ZN(W12293));
  NANDX1 G32640 (.A1(W2603), .A2(W15531), .ZN(W20757));
  NANDX1 G32641 (.A1(W752), .A2(W1753), .ZN(W3128));
  NANDX1 G32642 (.A1(W13475), .A2(W3285), .ZN(W20758));
  NANDX1 G32643 (.A1(W11812), .A2(I271), .ZN(W12291));
  NANDX1 G32644 (.A1(I1357), .A2(W15394), .ZN(W20760));
  NANDX1 G32645 (.A1(I4), .A2(I5), .ZN(W2));
  NANDX1 G32646 (.A1(W11313), .A2(W13646), .ZN(O2074));
  NANDX1 G32647 (.A1(W25240), .A2(W10813), .ZN(O3381));
  NANDX1 G32648 (.A1(I12), .A2(I13), .ZN(W6));
  NANDX1 G32649 (.A1(W705), .A2(W388), .ZN(W3127));
  NANDX1 G32650 (.A1(W4975), .A2(W3464), .ZN(W8788));
  NANDX1 G32651 (.A1(I514), .A2(I1577), .ZN(W3093));
  NANDX1 G32652 (.A1(W7440), .A2(W10702), .ZN(W20764));
  NANDX1 G32653 (.A1(W7083), .A2(W11951), .ZN(O590));
  NANDX1 G32654 (.A1(W3076), .A2(W15692), .ZN(W20767));
  NANDX1 G32655 (.A1(W22276), .A2(W18888), .ZN(O3380));
  NANDX1 G32656 (.A1(W5872), .A2(W10612), .ZN(W12286));
  NANDX1 G32657 (.A1(W12064), .A2(W3607), .ZN(W12285));
  NANDX1 G32658 (.A1(W2781), .A2(W10736), .ZN(W20771));
  NANDX1 G32659 (.A1(W8018), .A2(I1333), .ZN(W10191));
  NANDX1 G32660 (.A1(W2297), .A2(W846), .ZN(W3117));
  NANDX1 G32661 (.A1(W9311), .A2(W7115), .ZN(W12284));
  NANDX1 G32662 (.A1(W20531), .A2(W16310), .ZN(W20772));
  NANDX1 G32663 (.A1(W14528), .A2(W14425), .ZN(O2077));
  NANDX1 G32664 (.A1(W677), .A2(W7955), .ZN(W20775));
  NANDX1 G32665 (.A1(W7163), .A2(W469), .ZN(W10184));
  NANDX1 G32666 (.A1(W9860), .A2(W2219), .ZN(W20843));
  NANDX1 G32667 (.A1(W1887), .A2(W2236), .ZN(W3078));
  NANDX1 G32668 (.A1(I483), .A2(W1620), .ZN(W3077));
  NANDX1 G32669 (.A1(W7695), .A2(I1051), .ZN(W10204));
  NANDX1 G32670 (.A1(W181), .A2(I1953), .ZN(W3074));
  NANDX1 G32671 (.A1(W6919), .A2(W6982), .ZN(W12259));
  NANDX1 G32672 (.A1(W12057), .A2(W13728), .ZN(W20832));
  NANDX1 G32673 (.A1(W6716), .A2(W12387), .ZN(W20833));
  NANDX1 G32674 (.A1(I44), .A2(I45), .ZN(W22));
  NANDX1 G32675 (.A1(I80), .A2(W2920), .ZN(W3073));
  NANDX1 G32676 (.A1(W20260), .A2(W14010), .ZN(O2096));
  NANDX1 G32677 (.A1(W5183), .A2(W7727), .ZN(W8805));
  NANDX1 G32678 (.A1(W88), .A2(W1643), .ZN(W3071));
  NANDX1 G32679 (.A1(W3183), .A2(W7811), .ZN(W20838));
  NANDX1 G32680 (.A1(W11870), .A2(W3226), .ZN(O3364));
  NANDX1 G32681 (.A1(W10895), .A2(W10588), .ZN(W20827));
  NANDX1 G32682 (.A1(W14666), .A2(W18189), .ZN(O2098));
  NANDX1 G32683 (.A1(W4205), .A2(W1485), .ZN(O3363));
  NANDX1 G32684 (.A1(W24502), .A2(W124), .ZN(W25297));
  NANDX1 G32685 (.A1(W13427), .A2(W12854), .ZN(W20845));
  NANDX1 G32686 (.A1(W6120), .A2(W6417), .ZN(W12255));
  NANDX1 G32687 (.A1(W9862), .A2(W6609), .ZN(W12254));
  NANDX1 G32688 (.A1(W1607), .A2(W18111), .ZN(O3361));
  NANDX1 G32689 (.A1(W2957), .A2(I104), .ZN(W3068));
  NANDX1 G32690 (.A1(W1611), .A2(W7822), .ZN(W10207));
  NANDX1 G32691 (.A1(W9353), .A2(W4846), .ZN(W12252));
  NANDX1 G32692 (.A1(W15548), .A2(W22615), .ZN(W25293));
  NANDX1 G32693 (.A1(W1612), .A2(I1230), .ZN(W3065));
  NANDX1 G32694 (.A1(W7868), .A2(W17521), .ZN(W20847));
  NANDX1 G32695 (.A1(W14545), .A2(W18630), .ZN(W20850));
  NANDX1 G32696 (.A1(W6118), .A2(W2010), .ZN(W10203));
  NANDX1 G32697 (.A1(W17072), .A2(W8332), .ZN(W25323));
  NANDX1 G32698 (.A1(W19080), .A2(W23184), .ZN(O3373));
  NANDX1 G32699 (.A1(W480), .A2(W2286), .ZN(W12273));
  NANDX1 G32700 (.A1(W5134), .A2(W7126), .ZN(W10199));
  NANDX1 G32701 (.A1(W9035), .A2(W19623), .ZN(O3371));
  NANDX1 G32702 (.A1(I1636), .A2(W593), .ZN(W3090));
  NANDX1 G32703 (.A1(W4429), .A2(W9042), .ZN(W20800));
  NANDX1 G32704 (.A1(I1342), .A2(W3271), .ZN(O587));
  NANDX1 G32705 (.A1(W32), .A2(W6518), .ZN(W8801));
  NANDX1 G32706 (.A1(W17359), .A2(W14310), .ZN(O3370));
  NANDX1 G32707 (.A1(W10456), .A2(W1145), .ZN(O586));
  NANDX1 G32708 (.A1(W13307), .A2(W1686), .ZN(W25314));
  NANDX1 G32709 (.A1(W5443), .A2(W4824), .ZN(W8802));
  NANDX1 G32710 (.A1(W2084), .A2(W2093), .ZN(W8804));
  NANDX1 G32711 (.A1(W7336), .A2(W7572), .ZN(W12211));
  NANDX1 G32712 (.A1(W340), .A2(W15919), .ZN(W25311));
  NANDX1 G32713 (.A1(W16269), .A2(W5775), .ZN(O2088));
  NANDX1 G32714 (.A1(W8489), .A2(W6357), .ZN(W12267));
  NANDX1 G32715 (.A1(W9727), .A2(I676), .ZN(W25308));
  NANDX1 G32716 (.A1(W18539), .A2(W18660), .ZN(W20815));
  NANDX1 G32717 (.A1(W2878), .A2(W2355), .ZN(W12265));
  NANDX1 G32718 (.A1(W18602), .A2(W3780), .ZN(O2090));
  NANDX1 G32719 (.A1(W774), .A2(W1539), .ZN(W3083));
  NANDX1 G32720 (.A1(W6133), .A2(W5587), .ZN(W12264));
  NANDX1 G32721 (.A1(I38), .A2(I39), .ZN(W19));
  NANDX1 G32722 (.A1(W9760), .A2(W1347), .ZN(W20819));
  NANDX1 G32723 (.A1(W14277), .A2(W5019), .ZN(O3367));
  NANDX1 G32724 (.A1(W295), .A2(W1679), .ZN(O3365));
  NANDX1 G32725 (.A1(W8348), .A2(W2920), .ZN(W20824));
  NANDX1 G32726 (.A1(W398), .A2(W2492), .ZN(O25));
  NANDX1 G32727 (.A1(W1302), .A2(I575), .ZN(W2882));
  NANDX1 G32728 (.A1(W20254), .A2(W7594), .ZN(W21102));
  NANDX1 G32729 (.A1(W16287), .A2(W6842), .ZN(O2151));
  NANDX1 G32730 (.A1(W850), .A2(I832), .ZN(W2881));
  NANDX1 G32731 (.A1(I1962), .A2(W15027), .ZN(O2152));
  NANDX1 G32732 (.A1(I164), .A2(I165), .ZN(W82));
  NANDX1 G32733 (.A1(W24693), .A2(W2524), .ZN(O3328));
  NANDX1 G32734 (.A1(W16654), .A2(W9219), .ZN(W21115));
  NANDX1 G32735 (.A1(W1640), .A2(I398), .ZN(W10141));
  NANDX1 G32736 (.A1(I102), .A2(W10799), .ZN(W21120));
  NANDX1 G32737 (.A1(W2946), .A2(W7647), .ZN(W8891));
  NANDX1 G32738 (.A1(W18133), .A2(W2480), .ZN(W21121));
  NANDX1 G32739 (.A1(W13321), .A2(W8710), .ZN(W21122));
  NANDX1 G32740 (.A1(W770), .A2(W19926), .ZN(W21123));
  NANDX1 G32741 (.A1(W4877), .A2(W10018), .ZN(W12127));
  NANDX1 G32742 (.A1(W1876), .A2(W9022), .ZN(W25201));
  NANDX1 G32743 (.A1(W8102), .A2(W10285), .ZN(W12122));
  NANDX1 G32744 (.A1(W13483), .A2(W24869), .ZN(W25198));
  NANDX1 G32745 (.A1(I564), .A2(W10468), .ZN(W25197));
  NANDX1 G32746 (.A1(W166), .A2(I1121), .ZN(W2872));
  NANDX1 G32747 (.A1(W16911), .A2(W16210), .ZN(W25193));
  NANDX1 G32748 (.A1(W16399), .A2(I1633), .ZN(W25192));
  NANDX1 G32749 (.A1(W1914), .A2(W3900), .ZN(W12118));
  NANDX1 G32750 (.A1(W23342), .A2(W4663), .ZN(O3326));
  NANDX1 G32751 (.A1(W9485), .A2(W644), .ZN(W21131));
  NANDX1 G32752 (.A1(W16980), .A2(W9268), .ZN(W21132));
  NANDX1 G32753 (.A1(W9704), .A2(W9288), .ZN(O567));
  NANDX1 G32754 (.A1(W3742), .A2(W8055), .ZN(W21134));
  NANDX1 G32755 (.A1(I603), .A2(I1940), .ZN(W2867));
  NANDX1 G32756 (.A1(I681), .A2(W1828), .ZN(W25189));
  NANDX1 G32757 (.A1(W10184), .A2(W19199), .ZN(O2145));
  NANDX1 G32758 (.A1(W9685), .A2(W2866), .ZN(W10250));
  NANDX1 G32759 (.A1(I1022), .A2(I391), .ZN(W2900));
  NANDX1 G32760 (.A1(W9174), .A2(W14593), .ZN(W21073));
  NANDX1 G32761 (.A1(I1123), .A2(W959), .ZN(W12154));
  NANDX1 G32762 (.A1(W8296), .A2(W14637), .ZN(W21077));
  NANDX1 G32763 (.A1(W4247), .A2(W11922), .ZN(W12153));
  NANDX1 G32764 (.A1(W14981), .A2(W7442), .ZN(O3330));
  NANDX1 G32765 (.A1(W12562), .A2(W12556), .ZN(W21078));
  NANDX1 G32766 (.A1(W8467), .A2(W3314), .ZN(W10252));
  NANDX1 G32767 (.A1(W2214), .A2(W4164), .ZN(W8874));
  NANDX1 G32768 (.A1(W9420), .A2(W4021), .ZN(W10260));
  NANDX1 G32769 (.A1(W12996), .A2(W7636), .ZN(W21087));
  NANDX1 G32770 (.A1(W5981), .A2(W3746), .ZN(O571));
  NANDX1 G32771 (.A1(W13625), .A2(W22826), .ZN(W25211));
  NANDX1 G32772 (.A1(W3789), .A2(W5251), .ZN(W21136));
  NANDX1 G32773 (.A1(W3281), .A2(W5559), .ZN(W12139));
  NANDX1 G32774 (.A1(I144), .A2(I145), .ZN(W72));
  NANDX1 G32775 (.A1(W934), .A2(W1589), .ZN(W2889));
  NANDX1 G32776 (.A1(W14747), .A2(I1706), .ZN(W25210));
  NANDX1 G32777 (.A1(W4031), .A2(W1932), .ZN(O367));
  NANDX1 G32778 (.A1(W6466), .A2(W4253), .ZN(W10146));
  NANDX1 G32779 (.A1(W1366), .A2(I910), .ZN(W2886));
  NANDX1 G32780 (.A1(W9125), .A2(W4800), .ZN(O2146));
  NANDX1 G32781 (.A1(W24311), .A2(W5114), .ZN(W25207));
  NANDX1 G32782 (.A1(W2397), .A2(W6843), .ZN(W25206));
  NANDX1 G32783 (.A1(I156), .A2(I157), .ZN(W78));
  NANDX1 G32784 (.A1(W12215), .A2(W13482), .ZN(O2147));
  NANDX1 G32785 (.A1(I1562), .A2(I919), .ZN(W10266));
  NANDX1 G32786 (.A1(W12311), .A2(W797), .ZN(O2149));
  NANDX1 G32787 (.A1(W20473), .A2(W9612), .ZN(W21179));
  NANDX1 G32788 (.A1(W6218), .A2(W9891), .ZN(W21168));
  NANDX1 G32789 (.A1(W11143), .A2(W9839), .ZN(W21169));
  NANDX1 G32790 (.A1(W18768), .A2(W9960), .ZN(W21170));
  NANDX1 G32791 (.A1(W1645), .A2(W1548), .ZN(W2838));
  NANDX1 G32792 (.A1(W22018), .A2(W10921), .ZN(W25178));
  NANDX1 G32793 (.A1(W19847), .A2(W9592), .ZN(W21171));
  NANDX1 G32794 (.A1(W1676), .A2(W23100), .ZN(W25177));
  NANDX1 G32795 (.A1(W18907), .A2(W13128), .ZN(W21173));
  NANDX1 G32796 (.A1(W7072), .A2(W13917), .ZN(W21176));
  NANDX1 G32797 (.A1(I1954), .A2(W1130), .ZN(W2837));
  NANDX1 G32798 (.A1(W8706), .A2(W3977), .ZN(W8904));
  NANDX1 G32799 (.A1(I176), .A2(W2629), .ZN(W8905));
  NANDX1 G32800 (.A1(W5782), .A2(I1419), .ZN(W10276));
  NANDX1 G32801 (.A1(W18312), .A2(W12104), .ZN(W25175));
  NANDX1 G32802 (.A1(W986), .A2(W8357), .ZN(W12093));
  NANDX1 G32803 (.A1(I682), .A2(I1786), .ZN(W2840));
  NANDX1 G32804 (.A1(W18819), .A2(W19264), .ZN(W21180));
  NANDX1 G32805 (.A1(W6195), .A2(W9995), .ZN(W10277));
  NANDX1 G32806 (.A1(W8139), .A2(W16101), .ZN(O2172));
  NANDX1 G32807 (.A1(W13712), .A2(W13281), .ZN(O3321));
  NANDX1 G32808 (.A1(W10626), .A2(W5539), .ZN(W25172));
  NANDX1 G32809 (.A1(W4080), .A2(W2574), .ZN(W12091));
  NANDX1 G32810 (.A1(W16303), .A2(W11478), .ZN(W21183));
  NANDX1 G32811 (.A1(W8189), .A2(W4159), .ZN(W8906));
  NANDX1 G32812 (.A1(I194), .A2(I195), .ZN(W97));
  NANDX1 G32813 (.A1(I196), .A2(I197), .ZN(W98));
  NANDX1 G32814 (.A1(W7040), .A2(W6414), .ZN(O376));
  NANDX1 G32815 (.A1(W1513), .A2(W223), .ZN(W2830));
  NANDX1 G32816 (.A1(W774), .A2(I1459), .ZN(W2828));
  NANDX1 G32817 (.A1(I202), .A2(I203), .ZN(W101));
  NANDX1 G32818 (.A1(W17376), .A2(I612), .ZN(W25187));
  NANDX1 G32819 (.A1(I489), .A2(W5158), .ZN(W8896));
  NANDX1 G32820 (.A1(W4517), .A2(W6729), .ZN(W12110));
  NANDX1 G32821 (.A1(W4621), .A2(W7522), .ZN(W12107));
  NANDX1 G32822 (.A1(W13345), .A2(W13291), .ZN(O2160));
  NANDX1 G32823 (.A1(I1478), .A2(W1413), .ZN(W2862));
  NANDX1 G32824 (.A1(W16616), .A2(W7208), .ZN(W21143));
  NANDX1 G32825 (.A1(W4037), .A2(W1234), .ZN(W21144));
  NANDX1 G32826 (.A1(W2275), .A2(W2198), .ZN(W2861));
  NANDX1 G32827 (.A1(W2065), .A2(I785), .ZN(W2860));
  NANDX1 G32828 (.A1(W4964), .A2(W157), .ZN(O3324));
  NANDX1 G32829 (.A1(W21122), .A2(W2867), .ZN(O2161));
  NANDX1 G32830 (.A1(W5639), .A2(W687), .ZN(W12104));
  NANDX1 G32831 (.A1(W3140), .A2(W5408), .ZN(W21152));
  NANDX1 G32832 (.A1(W9319), .A2(W4348), .ZN(W12103));
  NANDX1 G32833 (.A1(I863), .A2(W8443), .ZN(W12158));
  NANDX1 G32834 (.A1(W23652), .A2(W15490), .ZN(W25186));
  NANDX1 G32835 (.A1(W9130), .A2(W5770), .ZN(O2163));
  NANDX1 G32836 (.A1(W25119), .A2(W16387), .ZN(W25185));
  NANDX1 G32837 (.A1(W4489), .A2(W9073), .ZN(W12100));
  NANDX1 G32838 (.A1(W10517), .A2(I332), .ZN(O2164));
  NANDX1 G32839 (.A1(W6124), .A2(W10091), .ZN(W10272));
  NANDX1 G32840 (.A1(W7919), .A2(W7266), .ZN(W8901));
  NANDX1 G32841 (.A1(W1230), .A2(W806), .ZN(W2856));
  NANDX1 G32842 (.A1(W16962), .A2(I525), .ZN(W21157));
  NANDX1 G32843 (.A1(W16498), .A2(W6126), .ZN(W21161));
  NANDX1 G32844 (.A1(I998), .A2(W209), .ZN(W2852));
  NANDX1 G32845 (.A1(W3134), .A2(I82), .ZN(W8902));
  NANDX1 G32846 (.A1(W1005), .A2(W793), .ZN(W12097));
  NANDX1 G32847 (.A1(I404), .A2(W535), .ZN(W2846));
  NANDX1 G32848 (.A1(W39), .A2(W787), .ZN(W21006));
  NANDX1 G32849 (.A1(I94), .A2(W1594), .ZN(W2956));
  NANDX1 G32850 (.A1(W5601), .A2(W2859), .ZN(O578));
  NANDX1 G32851 (.A1(W7077), .A2(I1566), .ZN(W20993));
  NANDX1 G32852 (.A1(W2922), .A2(W2323), .ZN(W8854));
  NANDX1 G32853 (.A1(W2745), .A2(W17273), .ZN(W25243));
  NANDX1 G32854 (.A1(W1654), .A2(W1053), .ZN(W2952));
  NANDX1 G32855 (.A1(W11618), .A2(W3611), .ZN(W20995));
  NANDX1 G32856 (.A1(W238), .A2(I858), .ZN(W2951));
  NANDX1 G32857 (.A1(W20170), .A2(I486), .ZN(O2132));
  NANDX1 G32858 (.A1(W5584), .A2(W15793), .ZN(W25242));
  NANDX1 G32859 (.A1(W8750), .A2(W2979), .ZN(W10235));
  NANDX1 G32860 (.A1(W10999), .A2(W4358), .ZN(W12198));
  NANDX1 G32861 (.A1(W8118), .A2(I1852), .ZN(W8856));
  NANDX1 G32862 (.A1(W19667), .A2(W6611), .ZN(W25241));
  NANDX1 G32863 (.A1(W218), .A2(W5118), .ZN(W10157));
  NANDX1 G32864 (.A1(W9654), .A2(W5875), .ZN(O3342));
  NANDX1 G32865 (.A1(I771), .A2(I874), .ZN(W2945));
  NANDX1 G32866 (.A1(W6417), .A2(W4320), .ZN(W21007));
  NANDX1 G32867 (.A1(I261), .A2(I1925), .ZN(W2944));
  NANDX1 G32868 (.A1(W4802), .A2(W2983), .ZN(W12193));
  NANDX1 G32869 (.A1(W3889), .A2(W4135), .ZN(O576));
  NANDX1 G32870 (.A1(W20156), .A2(W22179), .ZN(W25240));
  NANDX1 G32871 (.A1(W9914), .A2(W3183), .ZN(W10154));
  NANDX1 G32872 (.A1(W6827), .A2(I806), .ZN(O251));
  NANDX1 G32873 (.A1(W9722), .A2(I1665), .ZN(O2135));
  NANDX1 G32874 (.A1(W1410), .A2(I220), .ZN(W2933));
  NANDX1 G32875 (.A1(W16929), .A2(W8067), .ZN(W25239));
  NANDX1 G32876 (.A1(W17470), .A2(W4300), .ZN(W21013));
  NANDX1 G32877 (.A1(W5487), .A2(W9195), .ZN(W10153));
  NANDX1 G32878 (.A1(I771), .A2(W5761), .ZN(W12188));
  NANDX1 G32879 (.A1(W12149), .A2(W18988), .ZN(W20974));
  NANDX1 G32880 (.A1(W6029), .A2(W13623), .ZN(W20957));
  NANDX1 G32881 (.A1(W831), .A2(W2488), .ZN(W2971));
  NANDX1 G32882 (.A1(I1818), .A2(W1706), .ZN(W2970));
  NANDX1 G32883 (.A1(W2695), .A2(W9722), .ZN(W10164));
  NANDX1 G32884 (.A1(W6125), .A2(W3424), .ZN(W8846));
  NANDX1 G32885 (.A1(W2494), .A2(W14733), .ZN(W20961));
  NANDX1 G32886 (.A1(W2862), .A2(W887), .ZN(W2969));
  NANDX1 G32887 (.A1(W409), .A2(I1489), .ZN(W20962));
  NANDX1 G32888 (.A1(W2371), .A2(W3278), .ZN(W20966));
  NANDX1 G32889 (.A1(W1647), .A2(W3411), .ZN(W25251));
  NANDX1 G32890 (.A1(I244), .A2(W18022), .ZN(W20970));
  NANDX1 G32891 (.A1(W7190), .A2(I1662), .ZN(W8849));
  NANDX1 G32892 (.A1(W1358), .A2(W4190), .ZN(O2124));
  NANDX1 G32893 (.A1(W7414), .A2(W7138), .ZN(W8851));
  NANDX1 G32894 (.A1(W4012), .A2(W757), .ZN(W12185));
  NANDX1 G32895 (.A1(W774), .A2(W2910), .ZN(W2968));
  NANDX1 G32896 (.A1(W15066), .A2(W11637), .ZN(W20979));
  NANDX1 G32897 (.A1(W24710), .A2(W19129), .ZN(O3343));
  NANDX1 G32898 (.A1(W11750), .A2(W6353), .ZN(W20980));
  NANDX1 G32899 (.A1(W1623), .A2(W1787), .ZN(W2967));
  NANDX1 G32900 (.A1(I108), .A2(I109), .ZN(W54));
  NANDX1 G32901 (.A1(W1118), .A2(W6005), .ZN(O2129));
  NANDX1 G32902 (.A1(W935), .A2(I1828), .ZN(W2963));
  NANDX1 G32903 (.A1(W9666), .A2(W9262), .ZN(W20985));
  NANDX1 G32904 (.A1(W2720), .A2(W19405), .ZN(W25247));
  NANDX1 G32905 (.A1(I630), .A2(W278), .ZN(W2958));
  NANDX1 G32906 (.A1(I116), .A2(I117), .ZN(W58));
  NANDX1 G32907 (.A1(W3602), .A2(W5436), .ZN(W12204));
  NANDX1 G32908 (.A1(W8766), .A2(W595), .ZN(W10158));
  NANDX1 G32909 (.A1(W15964), .A2(W11529), .ZN(W21055));
  NANDX1 G32910 (.A1(W1518), .A2(W967), .ZN(W10247));
  NANDX1 G32911 (.A1(W13891), .A2(W15740), .ZN(W25231));
  NANDX1 G32912 (.A1(W7790), .A2(I257), .ZN(W25230));
  NANDX1 G32913 (.A1(W1836), .A2(I1345), .ZN(W10249));
  NANDX1 G32914 (.A1(W3888), .A2(I1008), .ZN(W12169));
  NANDX1 G32915 (.A1(W1358), .A2(W7943), .ZN(W21046));
  NANDX1 G32916 (.A1(I1419), .A2(W10472), .ZN(W12167));
  NANDX1 G32917 (.A1(W1992), .A2(W1724), .ZN(W2915));
  NANDX1 G32918 (.A1(W7472), .A2(W12543), .ZN(W21048));
  NANDX1 G32919 (.A1(W614), .A2(W3091), .ZN(O3337));
  NANDX1 G32920 (.A1(W1528), .A2(W436), .ZN(W2914));
  NANDX1 G32921 (.A1(W13425), .A2(W206), .ZN(O2140));
  NANDX1 G32922 (.A1(I826), .A2(W2271), .ZN(W2911));
  NANDX1 G32923 (.A1(W4114), .A2(W2555), .ZN(W12166));
  NANDX1 G32924 (.A1(W9966), .A2(W12418), .ZN(W21042));
  NANDX1 G32925 (.A1(W9220), .A2(W1804), .ZN(W12164));
  NANDX1 G32926 (.A1(W770), .A2(W19490), .ZN(W21056));
  NANDX1 G32927 (.A1(W1165), .A2(W260), .ZN(W21057));
  NANDX1 G32928 (.A1(W14704), .A2(W15306), .ZN(O2142));
  NANDX1 G32929 (.A1(I134), .A2(I135), .ZN(W67));
  NANDX1 G32930 (.A1(W9431), .A2(I1749), .ZN(O3334));
  NANDX1 G32931 (.A1(I136), .A2(I137), .ZN(W68));
  NANDX1 G32932 (.A1(W15958), .A2(I1386), .ZN(W21063));
  NANDX1 G32933 (.A1(W15176), .A2(W12785), .ZN(W21064));
  NANDX1 G32934 (.A1(W2144), .A2(I1002), .ZN(W2907));
  NANDX1 G32935 (.A1(W5022), .A2(W11759), .ZN(W12161));
  NANDX1 G32936 (.A1(W7510), .A2(W107), .ZN(W21067));
  NANDX1 G32937 (.A1(W6028), .A2(W10588), .ZN(W12160));
  NANDX1 G32938 (.A1(W4159), .A2(W1573), .ZN(W8871));
  NANDX1 G32939 (.A1(W20004), .A2(W11628), .ZN(O3340));
  NANDX1 G32940 (.A1(W2530), .A2(I376), .ZN(W2930));
  NANDX1 G32941 (.A1(W8956), .A2(W10828), .ZN(O574));
  NANDX1 G32942 (.A1(W5864), .A2(W7117), .ZN(W12183));
  NANDX1 G32943 (.A1(W4932), .A2(W5262), .ZN(W21018));
  NANDX1 G32944 (.A1(W7017), .A2(W19568), .ZN(W21020));
  NANDX1 G32945 (.A1(W14934), .A2(W5185), .ZN(W21021));
  NANDX1 G32946 (.A1(W4435), .A2(W10228), .ZN(W21023));
  NANDX1 G32947 (.A1(W15252), .A2(W1871), .ZN(O3341));
  NANDX1 G32948 (.A1(I1688), .A2(I1864), .ZN(W2926));
  NANDX1 G32949 (.A1(W3481), .A2(W7548), .ZN(W12179));
  NANDX1 G32950 (.A1(W10196), .A2(W17244), .ZN(W21026));
  NANDX1 G32951 (.A1(W7454), .A2(W10166), .ZN(W21027));
  NANDX1 G32952 (.A1(W473), .A2(W1758), .ZN(W2923));
  NANDX1 G32953 (.A1(W3508), .A2(W7516), .ZN(W21029));
  NANDX1 G32954 (.A1(W21084), .A2(W6415), .ZN(W22314));
  NANDX1 G32955 (.A1(W17500), .A2(W6032), .ZN(O2137));
  NANDX1 G32956 (.A1(W2319), .A2(W3398), .ZN(W21031));
  NANDX1 G32957 (.A1(W4597), .A2(W2558), .ZN(W12177));
  NANDX1 G32958 (.A1(W12139), .A2(W11862), .ZN(W12176));
  NANDX1 G32959 (.A1(W7800), .A2(W13119), .ZN(O2138));
  NANDX1 G32960 (.A1(W2563), .A2(W815), .ZN(W2922));
  NANDX1 G32961 (.A1(W4715), .A2(W7293), .ZN(W10242));
  NANDX1 G32962 (.A1(W8847), .A2(W18210), .ZN(W21035));
  NANDX1 G32963 (.A1(W8945), .A2(W8), .ZN(W25235));
  NANDX1 G32964 (.A1(W5462), .A2(W3077), .ZN(O573));
  NANDX1 G32965 (.A1(I1452), .A2(W5879), .ZN(W10245));
  NANDX1 G32966 (.A1(W17209), .A2(W17967), .ZN(W21039));
  NANDX1 G32967 (.A1(W18841), .A2(W8383), .ZN(W21041));
  NANDX1 G32968 (.A1(W9330), .A2(W9840), .ZN(W10246));
  NANDX1 G32969 (.A1(I1361), .A2(W1309), .ZN(W2175));
  NANDX1 G32970 (.A1(I501), .A2(W1110), .ZN(W11775));
  NANDX1 G32971 (.A1(W1549), .A2(I1979), .ZN(W2268));
  NANDX1 G32972 (.A1(W4130), .A2(W3714), .ZN(W11629));
  NANDX1 G32973 (.A1(W573), .A2(W8897), .ZN(O2444));
  NANDX1 G32974 (.A1(W9422), .A2(W10767), .ZN(W22136));
  NANDX1 G32975 (.A1(W6216), .A2(W10196), .ZN(W11704));
  NANDX1 G32976 (.A1(W8155), .A2(W5498), .ZN(O2372));
  NANDX1 G32977 (.A1(W59), .A2(W1854), .ZN(W11773));
  NANDX1 G32978 (.A1(W4566), .A2(W6026), .ZN(W11630));
  NANDX1 G32979 (.A1(W846), .A2(W6498), .ZN(W10054));
  NANDX1 G32980 (.A1(W1595), .A2(W2639), .ZN(W11772));
  NANDX1 G32981 (.A1(W8505), .A2(W7662), .ZN(W11626));
  NANDX1 G32982 (.A1(W1543), .A2(W179), .ZN(W2362));
  NANDX1 G32983 (.A1(W5308), .A2(W9068), .ZN(W22062));
  NANDX1 G32984 (.A1(W2886), .A2(W12350), .ZN(O2416));
  NANDX1 G32985 (.A1(W8834), .A2(W4273), .ZN(W24923));
  NANDX1 G32986 (.A1(W542), .A2(I26), .ZN(W2176));
  NANDX1 G32987 (.A1(W10175), .A2(W3581), .ZN(W11768));
  NANDX1 G32988 (.A1(W814), .A2(W739), .ZN(W2360));
  NANDX1 G32989 (.A1(W7644), .A2(W3128), .ZN(W11705));
  NANDX1 G32990 (.A1(W2309), .A2(I915), .ZN(W2358));
  NANDX1 G32991 (.A1(W10835), .A2(W973), .ZN(W11767));
  NANDX1 G32992 (.A1(W14655), .A2(W8229), .ZN(W22059));
  NANDX1 G32993 (.A1(W20468), .A2(W5242), .ZN(W21897));
  NANDX1 G32994 (.A1(W11074), .A2(W4579), .ZN(W11621));
  NANDX1 G32995 (.A1(W24295), .A2(W19090), .ZN(O3202));
  NANDX1 G32996 (.A1(W1307), .A2(W4749), .ZN(W11777));
  NANDX1 G32997 (.A1(W12130), .A2(W19204), .ZN(W21894));
  NANDX1 G32998 (.A1(I78), .A2(W1836), .ZN(W2368));
  NANDX1 G32999 (.A1(W6982), .A2(W8187), .ZN(O272));
  NANDX1 G33000 (.A1(I704), .A2(I705), .ZN(W352));
  NANDX1 G33001 (.A1(W5772), .A2(W8189), .ZN(W9227));
  NANDX1 G33002 (.A1(I564), .A2(I565), .ZN(W282));
  NANDX1 G33003 (.A1(W10589), .A2(W3460), .ZN(W21895));
  NANDX1 G33004 (.A1(W19024), .A2(W11433), .ZN(W21896));
  NANDX1 G33005 (.A1(W4200), .A2(W7408), .ZN(W11766));
  NANDX1 G33006 (.A1(I531), .A2(I1108), .ZN(W2367));
  NANDX1 G33007 (.A1(W20248), .A2(W16670), .ZN(W21898));
  NANDX1 G33008 (.A1(W7617), .A2(W3114), .ZN(W24925));
  NANDX1 G33009 (.A1(W10685), .A2(W6328), .ZN(W11623));
  NANDX1 G33010 (.A1(W1883), .A2(I1574), .ZN(W2216));
  NANDX1 G33011 (.A1(W4717), .A2(W3852), .ZN(W11624));
  NANDX1 G33012 (.A1(W10640), .A2(W18843), .ZN(O2370));
  NANDX1 G33013 (.A1(W2170), .A2(W137), .ZN(W2366));
  NANDX1 G33014 (.A1(W1099), .A2(W8727), .ZN(W22200));
  NANDX1 G33015 (.A1(W7473), .A2(W5710), .ZN(W24826));
  NANDX1 G33016 (.A1(I586), .A2(I587), .ZN(W293));
  NANDX1 G33017 (.A1(I580), .A2(I581), .ZN(W290));
  NANDX1 G33018 (.A1(W8874), .A2(I656), .ZN(W11761));
  NANDX1 G33019 (.A1(W4049), .A2(W12775), .ZN(W21920));
  NANDX1 G33020 (.A1(I816), .A2(I413), .ZN(W2182));
  NANDX1 G33021 (.A1(I799), .A2(W6224), .ZN(W9219));
  NANDX1 G33022 (.A1(W13699), .A2(W18808), .ZN(W21923));
  NANDX1 G33023 (.A1(W13152), .A2(W4800), .ZN(O2443));
  NANDX1 G33024 (.A1(W6161), .A2(W22863), .ZN(W24911));
  NANDX1 G33025 (.A1(W243), .A2(W1682), .ZN(W2186));
  NANDX1 G33026 (.A1(W993), .A2(W15871), .ZN(W24910));
  NANDX1 G33027 (.A1(W14029), .A2(W20333), .ZN(W21925));
  NANDX1 G33028 (.A1(W8909), .A2(W4149), .ZN(W9220));
  NANDX1 G33029 (.A1(W8011), .A2(W12511), .ZN(W24837));
  NANDX1 G33030 (.A1(W4390), .A2(I924), .ZN(W21926));
  NANDX1 G33031 (.A1(I692), .A2(I693), .ZN(W346));
  NANDX1 G33032 (.A1(W6476), .A2(I181), .ZN(W9216));
  NANDX1 G33033 (.A1(I1516), .A2(W530), .ZN(W2274));
  NANDX1 G33034 (.A1(I390), .A2(W2009), .ZN(W2348));
  NANDX1 G33035 (.A1(I622), .A2(I623), .ZN(W311));
  NANDX1 G33036 (.A1(W1321), .A2(I1860), .ZN(W2347));
  NANDX1 G33037 (.A1(W12119), .A2(W15197), .ZN(O2376));
  NANDX1 G33038 (.A1(W23181), .A2(W12420), .ZN(O3237));
  NANDX1 G33039 (.A1(W7796), .A2(W353), .ZN(W10396));
  NANDX1 G33040 (.A1(I574), .A2(I575), .ZN(W287));
  NANDX1 G33041 (.A1(W10763), .A2(I414), .ZN(W11631));
  NANDX1 G33042 (.A1(W3288), .A2(W1843), .ZN(W11632));
  NANDX1 G33043 (.A1(W50), .A2(W7974), .ZN(W11764));
  NANDX1 G33044 (.A1(I734), .A2(W11121), .ZN(W21913));
  NANDX1 G33045 (.A1(I666), .A2(W1455), .ZN(W2180));
  NANDX1 G33046 (.A1(W20498), .A2(W10062), .ZN(O2413));
  NANDX1 G33047 (.A1(W12486), .A2(W14939), .ZN(W21914));
  NANDX1 G33048 (.A1(W20584), .A2(W17712), .ZN(W24920));
  NANDX1 G33049 (.A1(W14080), .A2(W15999), .ZN(W24919));
  NANDX1 G33050 (.A1(I696), .A2(I697), .ZN(W348));
  NANDX1 G33051 (.A1(W22799), .A2(W2601), .ZN(W24868));
  NANDX1 G33052 (.A1(W24578), .A2(W747), .ZN(O3208));
  NANDX1 G33053 (.A1(W20027), .A2(W15303), .ZN(W21916));
  NANDX1 G33054 (.A1(W562), .A2(W895), .ZN(W11633));
  NANDX1 G33055 (.A1(W8327), .A2(W171), .ZN(O356));
  NANDX1 G33056 (.A1(W12858), .A2(W12045), .ZN(W22055));
  NANDX1 G33057 (.A1(I1434), .A2(W1195), .ZN(W2354));
  NANDX1 G33058 (.A1(W963), .A2(W3777), .ZN(W9130));
  NANDX1 G33059 (.A1(W1986), .A2(W1890), .ZN(W2272));
  NANDX1 G33060 (.A1(W17338), .A2(W9487), .ZN(W22191));
  NANDX1 G33061 (.A1(W7399), .A2(W5943), .ZN(O2431));
  NANDX1 G33062 (.A1(W1572), .A2(I583), .ZN(W10390));
  NANDX1 G33063 (.A1(W13776), .A2(W20547), .ZN(W24940));
  NANDX1 G33064 (.A1(W798), .A2(I1104), .ZN(W9119));
  NANDX1 G33065 (.A1(W6217), .A2(W521), .ZN(O354));
  NANDX1 G33066 (.A1(W2114), .A2(W10188), .ZN(W22076));
  NANDX1 G33067 (.A1(W12525), .A2(W5026), .ZN(O3221));
  NANDX1 G33068 (.A1(W15038), .A2(W10300), .ZN(W21859));
  NANDX1 G33069 (.A1(W7781), .A2(W5500), .ZN(W11794));
  NANDX1 G33070 (.A1(W8707), .A2(W8330), .ZN(W10026));
  NANDX1 G33071 (.A1(W17974), .A2(W11892), .ZN(W22219));
  NANDX1 G33072 (.A1(W3167), .A2(W10484), .ZN(W21860));
  NANDX1 G33073 (.A1(I916), .A2(I575), .ZN(W2263));
  NANDX1 G33074 (.A1(W11145), .A2(W8457), .ZN(W24818));
  NANDX1 G33075 (.A1(W599), .A2(W1893), .ZN(W2264));
  NANDX1 G33076 (.A1(W479), .A2(I594), .ZN(W2162));
  NANDX1 G33077 (.A1(W2273), .A2(W814), .ZN(W2386));
  NANDX1 G33078 (.A1(I718), .A2(I719), .ZN(W359));
  NANDX1 G33079 (.A1(W10228), .A2(I1886), .ZN(O525));
  NANDX1 G33080 (.A1(I532), .A2(I533), .ZN(W266));
  NANDX1 G33081 (.A1(I522), .A2(I1201), .ZN(W2385));
  NANDX1 G33082 (.A1(W9795), .A2(W4089), .ZN(W10027));
  NANDX1 G33083 (.A1(W7750), .A2(I176), .ZN(O537));
  NANDX1 G33084 (.A1(W3324), .A2(W5248), .ZN(W10435));
  NANDX1 G33085 (.A1(I534), .A2(I535), .ZN(W267));
  NANDX1 G33086 (.A1(W8065), .A2(W5930), .ZN(W9116));
  NANDX1 G33087 (.A1(I1982), .A2(I1584), .ZN(W2258));
  NANDX1 G33088 (.A1(W1021), .A2(W99), .ZN(W2156));
  NANDX1 G33089 (.A1(W4875), .A2(W8492), .ZN(O539));
  NANDX1 G33090 (.A1(W2395), .A2(I1684), .ZN(O266));
  NANDX1 G33091 (.A1(W8566), .A2(W4229), .ZN(W10388));
  NANDX1 G33092 (.A1(W5943), .A2(W9037), .ZN(O353));
  NANDX1 G33093 (.A1(W15023), .A2(W877), .ZN(W22223));
  NANDX1 G33094 (.A1(I660), .A2(I661), .ZN(O3));
  NANDX1 G33095 (.A1(I16), .A2(W650), .ZN(O538));
  NANDX1 G33096 (.A1(W6175), .A2(I670), .ZN(W11696));
  NANDX1 G33097 (.A1(I720), .A2(I721), .ZN(W360));
  NANDX1 G33098 (.A1(W6203), .A2(W1018), .ZN(W10434));
  NANDX1 G33099 (.A1(I1146), .A2(W2248), .ZN(W2259));
  NANDX1 G33100 (.A1(W2344), .A2(W4680), .ZN(W9117));
  NANDX1 G33101 (.A1(W523), .A2(W8326), .ZN(W9185));
  NANDX1 G33102 (.A1(W8386), .A2(W2017), .ZN(O357));
  NANDX1 G33103 (.A1(W3391), .A2(W9209), .ZN(W11670));
  NANDX1 G33104 (.A1(I550), .A2(W1306), .ZN(W2262));
  NANDX1 G33105 (.A1(I628), .A2(W7435), .ZN(W10060));
  NANDX1 G33106 (.A1(W7231), .A2(W5588), .ZN(W11798));
  NANDX1 G33107 (.A1(I953), .A2(W58), .ZN(W2218));
  NANDX1 G33108 (.A1(W7069), .A2(W2328), .ZN(W11796));
  NANDX1 G33109 (.A1(W14836), .A2(W5808), .ZN(O2365));
  NANDX1 G33110 (.A1(I1329), .A2(I1553), .ZN(W2265));
  NANDX1 G33111 (.A1(W2090), .A2(W865), .ZN(W2166));
  NANDX1 G33112 (.A1(W19339), .A2(W20429), .ZN(W22211));
  NANDX1 G33113 (.A1(W16776), .A2(W20327), .ZN(W22073));
  NANDX1 G33114 (.A1(W3989), .A2(W5349), .ZN(W11618));
  NANDX1 G33115 (.A1(W11127), .A2(W7545), .ZN(O2446));
  NANDX1 G33116 (.A1(W6028), .A2(W16492), .ZN(W22071));
  NANDX1 G33117 (.A1(W17347), .A2(W5475), .ZN(W22070));
  NANDX1 G33118 (.A1(W1216), .A2(W1989), .ZN(W2266));
  NANDX1 G33119 (.A1(W11992), .A2(I1209), .ZN(W21883));
  NANDX1 G33120 (.A1(W2774), .A2(W9349), .ZN(W10057));
  NANDX1 G33121 (.A1(W19636), .A2(W2423), .ZN(W21881));
  NANDX1 G33122 (.A1(W14266), .A2(W5241), .ZN(W22066));
  NANDX1 G33123 (.A1(W4059), .A2(W8571), .ZN(O2366));
  NANDX1 G33124 (.A1(I1459), .A2(W2061), .ZN(W10056));
  NANDX1 G33125 (.A1(W3422), .A2(W3374), .ZN(O2367));
  NANDX1 G33126 (.A1(W13245), .A2(W19775), .ZN(W22065));
  NANDX1 G33127 (.A1(W5963), .A2(W7023), .ZN(W11619));
  NANDX1 G33128 (.A1(I954), .A2(W411), .ZN(W2375));
  NANDX1 G33129 (.A1(W20587), .A2(W13911), .ZN(W24927));
  NANDX1 G33130 (.A1(W1992), .A2(I1497), .ZN(W2374));
  NANDX1 G33131 (.A1(W9312), .A2(W9438), .ZN(O2369));
  NANDX1 G33132 (.A1(I986), .A2(W3461), .ZN(W22215));
  NANDX1 G33133 (.A1(W7320), .A2(W10355), .ZN(O2357));
  NANDX1 G33134 (.A1(W6922), .A2(W850), .ZN(W11788));
  NANDX1 G33135 (.A1(I398), .A2(W8459), .ZN(W21870));
  NANDX1 G33136 (.A1(I1274), .A2(W1498), .ZN(W2383));
  NANDX1 G33137 (.A1(W19963), .A2(W13563), .ZN(W21872));
  NANDX1 G33138 (.A1(W11131), .A2(W586), .ZN(O3247));
  NANDX1 G33139 (.A1(W18541), .A2(W9944), .ZN(O2359));
  NANDX1 G33140 (.A1(I536), .A2(I537), .ZN(W268));
  NANDX1 G33141 (.A1(W1840), .A2(W3876), .ZN(O536));
  NANDX1 G33142 (.A1(I542), .A2(I543), .ZN(W271));
  NANDX1 G33143 (.A1(W18598), .A2(W8434), .ZN(O3222));
  NANDX1 G33144 (.A1(W4586), .A2(W162), .ZN(W11639));
  NANDX1 G33145 (.A1(W6703), .A2(W9813), .ZN(W10058));
  NANDX1 G33146 (.A1(I714), .A2(I715), .ZN(W357));
  NANDX1 G33147 (.A1(W121), .A2(W2159), .ZN(W2163));
  NANDX1 G33148 (.A1(W7934), .A2(W8625), .ZN(W21877));
  NANDX1 G33149 (.A1(W20915), .A2(W22837), .ZN(O3201));
  NANDX1 G33150 (.A1(W1912), .A2(I808), .ZN(W2381));
  NANDX1 G33151 (.A1(W1266), .A2(W19384), .ZN(W24933));
  NANDX1 G33152 (.A1(W4073), .A2(W3226), .ZN(W11781));
  NANDX1 G33153 (.A1(W3210), .A2(W2834), .ZN(W11780));
  NANDX1 G33154 (.A1(W2175), .A2(I1142), .ZN(W2378));
  NANDX1 G33155 (.A1(W11329), .A2(W17491), .ZN(W22009));
  NANDX1 G33156 (.A1(W18792), .A2(W4507), .ZN(W22048));
  NANDX1 G33157 (.A1(I1776), .A2(W1754), .ZN(W2199));
  NANDX1 G33158 (.A1(W9897), .A2(W8278), .ZN(W11734));
  NANDX1 G33159 (.A1(W2037), .A2(W8052), .ZN(W11733));
  NANDX1 G33160 (.A1(W14299), .A2(W11440), .ZN(W22004));
  NANDX1 G33161 (.A1(W2468), .A2(W7699), .ZN(O527));
  NANDX1 G33162 (.A1(W6996), .A2(W6807), .ZN(W10034));
  NANDX1 G33163 (.A1(W2267), .A2(I1243), .ZN(W2283));
  NANDX1 G33164 (.A1(W12792), .A2(W13256), .ZN(W24880));
  NANDX1 G33165 (.A1(W5380), .A2(W19039), .ZN(O2396));
  NANDX1 G33166 (.A1(W352), .A2(W1611), .ZN(W2201));
  NANDX1 G33167 (.A1(W6943), .A2(W10868), .ZN(O2411));
  NANDX1 G33168 (.A1(W10745), .A2(W14760), .ZN(O3227));
  NANDX1 G33169 (.A1(W79), .A2(I91), .ZN(W2310));
  NANDX1 G33170 (.A1(W6524), .A2(W1233), .ZN(W11664));
  NANDX1 G33171 (.A1(W1513), .A2(W4927), .ZN(W11729));
  NANDX1 G33172 (.A1(W545), .A2(W2484), .ZN(W9201));
  NANDX1 G33173 (.A1(W4399), .A2(W5219), .ZN(W11728));
  NANDX1 G33174 (.A1(W12426), .A2(W12269), .ZN(W22147));
  NANDX1 G33175 (.A1(W21026), .A2(W113), .ZN(O2398));
  NANDX1 G33176 (.A1(W1011), .A2(W19838), .ZN(W22150));
  NANDX1 G33177 (.A1(I477), .A2(W5274), .ZN(W22151));
  NANDX1 G33178 (.A1(I693), .A2(I1948), .ZN(O2399));
  NANDX1 G33179 (.A1(W9079), .A2(W19909), .ZN(W21998));
  NANDX1 G33180 (.A1(I292), .A2(W9614), .ZN(W21990));
  NANDX1 G33181 (.A1(W19194), .A2(W12655), .ZN(O3213));
  NANDX1 G33182 (.A1(I596), .A2(I597), .ZN(W298));
  NANDX1 G33183 (.A1(W366), .A2(W9887), .ZN(W24885));
  NANDX1 G33184 (.A1(I124), .A2(W808), .ZN(W2282));
  NANDX1 G33185 (.A1(W2797), .A2(I1051), .ZN(W9145));
  NANDX1 G33186 (.A1(I1409), .A2(W6523), .ZN(O268));
  NANDX1 G33187 (.A1(I277), .A2(W11702), .ZN(W21995));
  NANDX1 G33188 (.A1(W3527), .A2(W16629), .ZN(O3228));
  NANDX1 G33189 (.A1(I212), .A2(W1855), .ZN(W2321));
  NANDX1 G33190 (.A1(W13145), .A2(W12645), .ZN(W21996));
  NANDX1 G33191 (.A1(W2194), .A2(W9083), .ZN(W10412));
  NANDX1 G33192 (.A1(W6845), .A2(W9010), .ZN(W10409));
  NANDX1 G33193 (.A1(W49), .A2(I1617), .ZN(W2320));
  NANDX1 G33194 (.A1(W8533), .A2(W21862), .ZN(W21999));
  NANDX1 G33195 (.A1(I600), .A2(I601), .ZN(W300));
  NANDX1 G33196 (.A1(I270), .A2(W1250), .ZN(W2319));
  NANDX1 G33197 (.A1(W1823), .A2(I871), .ZN(O2394));
  NANDX1 G33198 (.A1(W2315), .A2(W1026), .ZN(W2318));
  NANDX1 G33199 (.A1(W12635), .A2(W4279), .ZN(W24882));
  NANDX1 G33200 (.A1(W718), .A2(W8299), .ZN(W9203));
  NANDX1 G33201 (.A1(W1622), .A2(W2256), .ZN(W2317));
  NANDX1 G33202 (.A1(W15599), .A2(W7634), .ZN(O2409));
  NANDX1 G33203 (.A1(W19854), .A2(W6777), .ZN(O2405));
  NANDX1 G33204 (.A1(I602), .A2(I603), .ZN(W301));
  NANDX1 G33205 (.A1(I604), .A2(I605), .ZN(W302));
  NANDX1 G33206 (.A1(W8318), .A2(W11572), .ZN(W22026));
  NANDX1 G33207 (.A1(W9757), .A2(W4317), .ZN(W22027));
  NANDX1 G33208 (.A1(W9190), .A2(W15064), .ZN(W22028));
  NANDX1 G33209 (.A1(W1843), .A2(I34), .ZN(W2298));
  NANDX1 G33210 (.A1(W9363), .A2(W9310), .ZN(W11724));
  NANDX1 G33211 (.A1(W15006), .A2(W219), .ZN(W22032));
  NANDX1 G33212 (.A1(W7640), .A2(W8244), .ZN(W9163));
  NANDX1 G33213 (.A1(W101), .A2(W558), .ZN(O270));
  NANDX1 G33214 (.A1(W11222), .A2(W1617), .ZN(W22023));
  NANDX1 G33215 (.A1(I401), .A2(I778), .ZN(W2297));
  NANDX1 G33216 (.A1(W393), .A2(I322), .ZN(W2208));
  NANDX1 G33217 (.A1(W1782), .A2(W1520), .ZN(W2209));
  NANDX1 G33218 (.A1(I608), .A2(I609), .ZN(W304));
  NANDX1 G33219 (.A1(I1600), .A2(W1250), .ZN(O533));
  NANDX1 G33220 (.A1(W11484), .A2(W21583), .ZN(W22153));
  NANDX1 G33221 (.A1(W10997), .A2(W11101), .ZN(W11719));
  NANDX1 G33222 (.A1(W6), .A2(W939), .ZN(W2292));
  NANDX1 G33223 (.A1(I500), .A2(I1582), .ZN(W2210));
  NANDX1 G33224 (.A1(W2067), .A2(I988), .ZN(W2294));
  NANDX1 G33225 (.A1(W4722), .A2(W14779), .ZN(O2401));
  NANDX1 G33226 (.A1(W728), .A2(W341), .ZN(W2305));
  NANDX1 G33227 (.A1(W3230), .A2(W2990), .ZN(W11667));
  NANDX1 G33228 (.A1(W652), .A2(W8860), .ZN(W9149));
  NANDX1 G33229 (.A1(W1859), .A2(I145), .ZN(W2303));
  NANDX1 G33230 (.A1(I592), .A2(W1046), .ZN(W2302));
  NANDX1 G33231 (.A1(W16686), .A2(W585), .ZN(W22045));
  NANDX1 G33232 (.A1(W3400), .A2(W6977), .ZN(W9166));
  NANDX1 G33233 (.A1(W313), .A2(I904), .ZN(W2212));
  NANDX1 G33234 (.A1(W703), .A2(I1874), .ZN(W2203));
  NANDX1 G33235 (.A1(W5817), .A2(I1156), .ZN(O2400));
  NANDX1 G33236 (.A1(W5206), .A2(I1963), .ZN(W24847));
  NANDX1 G33237 (.A1(W1668), .A2(W6168), .ZN(W21989));
  NANDX1 G33238 (.A1(W20698), .A2(I731), .ZN(W22159));
  NANDX1 G33239 (.A1(W1130), .A2(W14908), .ZN(O2402));
  NANDX1 G33240 (.A1(W1200), .A2(I1064), .ZN(W2300));
  NANDX1 G33241 (.A1(W9683), .A2(W5620), .ZN(W11716));
  NANDX1 G33242 (.A1(W1151), .A2(I1247), .ZN(W2289));
  NANDX1 G33243 (.A1(W6696), .A2(W4170), .ZN(W9199));
  NANDX1 G33244 (.A1(W873), .A2(W8325), .ZN(W10413));
  NANDX1 G33245 (.A1(I208), .A2(I1052), .ZN(W2299));
  NANDX1 G33246 (.A1(W531), .A2(W12752), .ZN(O2403));
  NANDX1 G33247 (.A1(W1194), .A2(W1257), .ZN(W2211));
  NANDX1 G33248 (.A1(W12540), .A2(W8034), .ZN(W21953));
  NANDX1 G33249 (.A1(I1329), .A2(W7674), .ZN(W11753));
  NANDX1 G33250 (.A1(I313), .A2(W7796), .ZN(W21947));
  NANDX1 G33251 (.A1(I698), .A2(W819), .ZN(W2340));
  NANDX1 G33252 (.A1(W3339), .A2(W22145), .ZN(O2440));
  NANDX1 G33253 (.A1(W7750), .A2(W2233), .ZN(W10404));
  NANDX1 G33254 (.A1(W16820), .A2(W4546), .ZN(O2383));
  NANDX1 G33255 (.A1(I4), .A2(W700), .ZN(W2339));
  NANDX1 G33256 (.A1(W16563), .A2(W4414), .ZN(W21951));
  NANDX1 G33257 (.A1(W3698), .A2(W9317), .ZN(W11752));
  NANDX1 G33258 (.A1(W14510), .A2(W12686), .ZN(W22144));
  NANDX1 G33259 (.A1(W2619), .A2(W11064), .ZN(W11714));
  NANDX1 G33260 (.A1(W112), .A2(W2106), .ZN(W2343));
  NANDX1 G33261 (.A1(W15666), .A2(W8301), .ZN(O3235));
  NANDX1 G33262 (.A1(I368), .A2(W8285), .ZN(W9209));
  NANDX1 G33263 (.A1(I838), .A2(W4159), .ZN(W11749));
  NANDX1 G33264 (.A1(W15207), .A2(W12178), .ZN(W21957));
  NANDX1 G33265 (.A1(W17914), .A2(W14275), .ZN(W21960));
  NANDX1 G33266 (.A1(W4793), .A2(W8154), .ZN(W22179));
  NANDX1 G33267 (.A1(W36), .A2(W2719), .ZN(W10033));
  NANDX1 G33268 (.A1(W4529), .A2(W9409), .ZN(W11747));
  NANDX1 G33269 (.A1(W559), .A2(W4939), .ZN(W22177));
  NANDX1 G33270 (.A1(W21459), .A2(W20837), .ZN(O2433));
  NANDX1 G33271 (.A1(W7653), .A2(W4855), .ZN(W21937));
  NANDX1 G33272 (.A1(W7997), .A2(I161), .ZN(W21931));
  NANDX1 G33273 (.A1(I690), .A2(I691), .ZN(W345));
  NANDX1 G33274 (.A1(W10048), .A2(W142), .ZN(W11711));
  NANDX1 G33275 (.A1(I124), .A2(W1425), .ZN(W2346));
  NANDX1 G33276 (.A1(W12618), .A2(W1970), .ZN(W22184));
  NANDX1 G33277 (.A1(W133), .A2(W6459), .ZN(W11759));
  NANDX1 G33278 (.A1(W19479), .A2(W13776), .ZN(W22183));
  NANDX1 G33279 (.A1(W8021), .A2(W18182), .ZN(O2378));
  NANDX1 G33280 (.A1(W11718), .A2(W16166), .ZN(W21935));
  NANDX1 G33281 (.A1(W2654), .A2(W21901), .ZN(O2379));
  NANDX1 G33282 (.A1(I1934), .A2(I1503), .ZN(W2345));
  NANDX1 G33283 (.A1(W7448), .A2(W8113), .ZN(W11743));
  NANDX1 G33284 (.A1(I1211), .A2(W10611), .ZN(W11713));
  NANDX1 G33285 (.A1(W9980), .A2(W19706), .ZN(W22143));
  NANDX1 G33286 (.A1(W13246), .A2(W6481), .ZN(W21938));
  NANDX1 G33287 (.A1(W1800), .A2(W2223), .ZN(W10048));
  NANDX1 G33288 (.A1(W4638), .A2(W4569), .ZN(W9213));
  NANDX1 G33289 (.A1(W2030), .A2(W2996), .ZN(W11757));
  NANDX1 G33290 (.A1(I664), .A2(I665), .ZN(W332));
  NANDX1 G33291 (.A1(W2490), .A2(W4947), .ZN(W10399));
  NANDX1 G33292 (.A1(W6650), .A2(W3937), .ZN(W9136));
  NANDX1 G33293 (.A1(I191), .A2(W7191), .ZN(W9212));
  NANDX1 G33294 (.A1(W6998), .A2(W7093), .ZN(W10416));
  NANDX1 G33295 (.A1(W14644), .A2(W24703), .ZN(W24893));
  NANDX1 G33296 (.A1(I196), .A2(I1425), .ZN(W2196));
  NANDX1 G33297 (.A1(I594), .A2(I595), .ZN(W297));
  NANDX1 G33298 (.A1(W10255), .A2(W6293), .ZN(W21980));
  NANDX1 G33299 (.A1(W24), .A2(W23545), .ZN(O3211));
  NANDX1 G33300 (.A1(W16638), .A2(W10629), .ZN(W22165));
  NANDX1 G33301 (.A1(I1714), .A2(I479), .ZN(W9206));
  NANDX1 G33302 (.A1(W7343), .A2(W1097), .ZN(W9142));
  NANDX1 G33303 (.A1(W60), .A2(W1751), .ZN(W2279));
  NANDX1 G33304 (.A1(I1919), .A2(W7833), .ZN(W24892));
  NANDX1 G33305 (.A1(W7814), .A2(W629), .ZN(W22050));
  NANDX1 G33306 (.A1(W1059), .A2(W16493), .ZN(W21977));
  NANDX1 G33307 (.A1(I684), .A2(I685), .ZN(W342));
  NANDX1 G33308 (.A1(W2593), .A2(W21008), .ZN(W24891));
  NANDX1 G33309 (.A1(W6957), .A2(W16620), .ZN(W21985));
  NANDX1 G33310 (.A1(W7003), .A2(I1738), .ZN(W11738));
  NANDX1 G33311 (.A1(W1950), .A2(I1003), .ZN(W2323));
  NANDX1 G33312 (.A1(W4130), .A2(W24712), .ZN(W24890));
  NANDX1 G33313 (.A1(W11616), .A2(W4916), .ZN(W22162));
  NANDX1 G33314 (.A1(W13365), .A2(W13730), .ZN(W21673));
  NANDX1 G33315 (.A1(W23436), .A2(W9442), .ZN(W24888));
  NANDX1 G33316 (.A1(W5975), .A2(W8914), .ZN(W9168));
  NANDX1 G33317 (.A1(W2544), .A2(I880), .ZN(O3231));
  NANDX1 G33318 (.A1(W21368), .A2(W8019), .ZN(W21965));
  NANDX1 G33319 (.A1(W7117), .A2(W21309), .ZN(O2439));
  NANDX1 G33320 (.A1(W10770), .A2(I1811), .ZN(W22052));
  NANDX1 G33321 (.A1(W13059), .A2(W6573), .ZN(O3232));
  NANDX1 G33322 (.A1(W4820), .A2(W6981), .ZN(W11650));
  NANDX1 G33323 (.A1(W24058), .A2(W19777), .ZN(W24839));
  NANDX1 G33324 (.A1(W7745), .A2(I718), .ZN(W11742));
  NANDX1 G33325 (.A1(W175), .A2(I434), .ZN(W11741));
  NANDX1 G33326 (.A1(W143), .A2(I1352), .ZN(O2390));
  NANDX1 G33327 (.A1(W9670), .A2(W8029), .ZN(W11654));
  NANDX1 G33328 (.A1(W4462), .A2(W798), .ZN(W9141));
  NANDX1 G33329 (.A1(W1517), .A2(I1557), .ZN(W2158));
  NANDX1 G33330 (.A1(I1042), .A2(I1604), .ZN(W21971));
  NANDX1 G33331 (.A1(W7584), .A2(I421), .ZN(W11655));
  NANDX1 G33332 (.A1(W15939), .A2(W24804), .ZN(W24894));
  NANDX1 G33333 (.A1(W5782), .A2(W19356), .ZN(W22171));
  NANDX1 G33334 (.A1(W19824), .A2(W6723), .ZN(W21972));
  NANDX1 G33335 (.A1(W5352), .A2(W15116), .ZN(O2391));
  NANDX1 G33336 (.A1(W1382), .A2(I1558), .ZN(W2328));
  NANDX1 G33337 (.A1(I686), .A2(I687), .ZN(W343));
  NANDX1 G33338 (.A1(W14891), .A2(W18872), .ZN(W24869));
  NANDX1 G33339 (.A1(W943), .A2(W1703), .ZN(W2327));
  NANDX1 G33340 (.A1(W1005), .A2(W725), .ZN(W2112));
  NANDX1 G33341 (.A1(W12047), .A2(W14944), .ZN(W21730));
  NANDX1 G33342 (.A1(W7959), .A2(W9083), .ZN(W10077));
  NANDX1 G33343 (.A1(W189), .A2(W2967), .ZN(W9194));
  NANDX1 G33344 (.A1(W21531), .A2(W1018), .ZN(W22102));
  NANDX1 G33345 (.A1(W10489), .A2(W6225), .ZN(W24800));
  NANDX1 G33346 (.A1(W12718), .A2(W11941), .ZN(W21731));
  NANDX1 G33347 (.A1(I782), .A2(W11698), .ZN(W24982));
  NANDX1 G33348 (.A1(W5811), .A2(W3379), .ZN(W22101));
  NANDX1 G33349 (.A1(W3876), .A2(W1573), .ZN(W24981));
  NANDX1 G33350 (.A1(W6192), .A2(W13108), .ZN(W21734));
  NANDX1 G33351 (.A1(I746), .A2(I747), .ZN(W373));
  NANDX1 G33352 (.A1(I1606), .A2(I82), .ZN(W2108));
  NANDX1 G33353 (.A1(W66), .A2(W393), .ZN(W2116));
  NANDX1 G33354 (.A1(W20111), .A2(W1193), .ZN(W21735));
  NANDX1 G33355 (.A1(W1025), .A2(I575), .ZN(W2480));
  NANDX1 G33356 (.A1(W8274), .A2(W12958), .ZN(W22099));
  NANDX1 G33357 (.A1(W4732), .A2(W6234), .ZN(W22098));
  NANDX1 G33358 (.A1(I1463), .A2(W7261), .ZN(W11597));
  NANDX1 G33359 (.A1(W24574), .A2(W24740), .ZN(W24979));
  NANDX1 G33360 (.A1(W9872), .A2(W13972), .ZN(W24859));
  NANDX1 G33361 (.A1(W5053), .A2(I1001), .ZN(W11892));
  NANDX1 G33362 (.A1(I459), .A2(W246), .ZN(W2119));
  NANDX1 G33363 (.A1(I1926), .A2(W675), .ZN(W2245));
  NANDX1 G33364 (.A1(W7796), .A2(W429), .ZN(W9256));
  NANDX1 G33365 (.A1(W7999), .A2(W9124), .ZN(W21719));
  NANDX1 G33366 (.A1(I1903), .A2(W17902), .ZN(W22291));
  NANDX1 G33367 (.A1(I456), .A2(I457), .ZN(W228));
  NANDX1 G33368 (.A1(W7320), .A2(W6990), .ZN(W22122));
  NANDX1 G33369 (.A1(W221), .A2(W903), .ZN(W2483));
  NANDX1 G33370 (.A1(W4680), .A2(W2808), .ZN(W21723));
  NANDX1 G33371 (.A1(W1883), .A2(I1552), .ZN(W2244));
  NANDX1 G33372 (.A1(W5066), .A2(W11203), .ZN(W11896));
  NANDX1 G33373 (.A1(W7531), .A2(I673), .ZN(W10373));
  NANDX1 G33374 (.A1(I1926), .A2(W10174), .ZN(W24794));
  NANDX1 G33375 (.A1(W2799), .A2(W8151), .ZN(O2321));
  NANDX1 G33376 (.A1(W8033), .A2(I920), .ZN(O2469));
  NANDX1 G33377 (.A1(W1904), .A2(W550), .ZN(W2107));
  NANDX1 G33378 (.A1(I1121), .A2(W7499), .ZN(W21725));
  NANDX1 G33379 (.A1(W20620), .A2(W20230), .ZN(W21726));
  NANDX1 G33380 (.A1(W4823), .A2(W19323), .ZN(W21727));
  NANDX1 G33381 (.A1(I595), .A2(W1958), .ZN(W2481));
  NANDX1 G33382 (.A1(W5825), .A2(W24180), .ZN(W24797));
  NANDX1 G33383 (.A1(W11421), .A2(W17962), .ZN(W22288));
  NANDX1 G33384 (.A1(W9936), .A2(W8362), .ZN(W21729));
  NANDX1 G33385 (.A1(I1102), .A2(I1092), .ZN(W2247));
  NANDX1 G33386 (.A1(I1051), .A2(W18676), .ZN(O3215));
  NANDX1 G33387 (.A1(W1987), .A2(I514), .ZN(W2228));
  NANDX1 G33388 (.A1(W19), .A2(W3385), .ZN(W10378));
  NANDX1 G33389 (.A1(W11358), .A2(W5773), .ZN(W11885));
  NANDX1 G33390 (.A1(W9208), .A2(W9068), .ZN(O2327));
  NANDX1 G33391 (.A1(I506), .A2(I370), .ZN(W2125));
  NANDX1 G33392 (.A1(W765), .A2(I877), .ZN(W2463));
  NANDX1 G33393 (.A1(W3142), .A2(W865), .ZN(W11883));
  NANDX1 G33394 (.A1(W544), .A2(W81), .ZN(W2460));
  NANDX1 G33395 (.A1(W6205), .A2(W13414), .ZN(W21762));
  NANDX1 G33396 (.A1(W3091), .A2(W12991), .ZN(W21763));
  NANDX1 G33397 (.A1(I878), .A2(W7871), .ZN(W10379));
  NANDX1 G33398 (.A1(I342), .A2(I998), .ZN(W2466));
  NANDX1 G33399 (.A1(W616), .A2(W1893), .ZN(W2458));
  NANDX1 G33400 (.A1(W8665), .A2(W6880), .ZN(O262));
  NANDX1 G33401 (.A1(I285), .A2(W3056), .ZN(W9189));
  NANDX1 G33402 (.A1(I346), .A2(W1988), .ZN(W9081));
  NANDX1 G33403 (.A1(W21400), .A2(W9288), .ZN(W24974));
  NANDX1 G33404 (.A1(W7583), .A2(I1380), .ZN(O276));
  NANDX1 G33405 (.A1(W10471), .A2(W10889), .ZN(W22273));
  NANDX1 G33406 (.A1(W4440), .A2(W12654), .ZN(W22271));
  NANDX1 G33407 (.A1(W7709), .A2(W9365), .ZN(W21767));
  NANDX1 G33408 (.A1(W14990), .A2(W20133), .ZN(W21768));
  NANDX1 G33409 (.A1(W66), .A2(I432), .ZN(W2472));
  NANDX1 G33410 (.A1(W14671), .A2(I176), .ZN(O2424));
  NANDX1 G33411 (.A1(W12160), .A2(W8557), .ZN(O2322));
  NANDX1 G33412 (.A1(I901), .A2(W695), .ZN(W2477));
  NANDX1 G33413 (.A1(W18208), .A2(W6974), .ZN(O2323));
  NANDX1 G33414 (.A1(W11327), .A2(W4635), .ZN(W22124));
  NANDX1 G33415 (.A1(W2421), .A2(W1631), .ZN(W2476));
  NANDX1 G33416 (.A1(I963), .A2(W464), .ZN(W10377));
  NANDX1 G33417 (.A1(W8980), .A2(W5411), .ZN(W9249));
  NANDX1 G33418 (.A1(I470), .A2(I471), .ZN(W235));
  NANDX1 G33419 (.A1(W14309), .A2(W16496), .ZN(W22277));
  NANDX1 G33420 (.A1(W21703), .A2(W9376), .ZN(W21748));
  NANDX1 G33421 (.A1(W1981), .A2(I1422), .ZN(W2484));
  NANDX1 G33422 (.A1(W8556), .A2(W4303), .ZN(W10074));
  NANDX1 G33423 (.A1(W9011), .A2(W9880), .ZN(W11889));
  NANDX1 G33424 (.A1(W10540), .A2(I236), .ZN(W21752));
  NANDX1 G33425 (.A1(I1135), .A2(W709), .ZN(W2469));
  NANDX1 G33426 (.A1(I1939), .A2(I1814), .ZN(W2468));
  NANDX1 G33427 (.A1(W1798), .A2(W3991), .ZN(O2325));
  NANDX1 G33428 (.A1(I474), .A2(I475), .ZN(O2));
  NANDX1 G33429 (.A1(W438), .A2(W895), .ZN(W2467));
  NANDX1 G33430 (.A1(I977), .A2(W19683), .ZN(W22275));
  NANDX1 G33431 (.A1(W5411), .A2(W7711), .ZN(W9190));
  NANDX1 G33432 (.A1(W9582), .A2(W9541), .ZN(W11586));
  NANDX1 G33433 (.A1(W197), .A2(W2086), .ZN(W2238));
  NANDX1 G33434 (.A1(W4406), .A2(W12058), .ZN(W22308));
  NANDX1 G33435 (.A1(I401), .A2(W2649), .ZN(W11686));
  NANDX1 G33436 (.A1(W589), .A2(I981), .ZN(W2508));
  NANDX1 G33437 (.A1(W4094), .A2(W20328), .ZN(O3194));
  NANDX1 G33438 (.A1(W1403), .A2(W1323), .ZN(W2239));
  NANDX1 G33439 (.A1(W1358), .A2(W654), .ZN(W2507));
  NANDX1 G33440 (.A1(W14160), .A2(W12386), .ZN(O2428));
  NANDX1 G33441 (.A1(W9397), .A2(W22505), .ZN(W24790));
  NANDX1 G33442 (.A1(I1032), .A2(I1229), .ZN(W2087));
  NANDX1 G33443 (.A1(I1441), .A2(W1049), .ZN(W2505));
  NANDX1 G33444 (.A1(I595), .A2(W12081), .ZN(W24996));
  NANDX1 G33445 (.A1(W6633), .A2(W15424), .ZN(O2473));
  NANDX1 G33446 (.A1(W18413), .A2(W11897), .ZN(O2312));
  NANDX1 G33447 (.A1(I357), .A2(I956), .ZN(W2241));
  NANDX1 G33448 (.A1(W3899), .A2(W4500), .ZN(W11901));
  NANDX1 G33449 (.A1(W8414), .A2(W6716), .ZN(W9073));
  NANDX1 G33450 (.A1(W22372), .A2(W18555), .ZN(W24791));
  NANDX1 G33451 (.A1(I1126), .A2(W11063), .ZN(W21696));
  NANDX1 G33452 (.A1(W16135), .A2(W10171), .ZN(O2472));
  NANDX1 G33453 (.A1(W101), .A2(W368), .ZN(W2088));
  NANDX1 G33454 (.A1(W7464), .A2(W6304), .ZN(W21697));
  NANDX1 G33455 (.A1(W2014), .A2(I813), .ZN(W2084));
  NANDX1 G33456 (.A1(I654), .A2(I655), .ZN(W327));
  NANDX1 G33457 (.A1(W240), .A2(I444), .ZN(W2511));
  NANDX1 G33458 (.A1(W5619), .A2(W4652), .ZN(W9193));
  NANDX1 G33459 (.A1(W7502), .A2(I78), .ZN(W10446));
  NANDX1 G33460 (.A1(I284), .A2(W14857), .ZN(W21675));
  NANDX1 G33461 (.A1(W2090), .A2(W2064), .ZN(O2426));
  NANDX1 G33462 (.A1(W3369), .A2(W21751), .ZN(O2478));
  NANDX1 G33463 (.A1(W12939), .A2(W21440), .ZN(W21676));
  NANDX1 G33464 (.A1(W14253), .A2(W89), .ZN(W21677));
  NANDX1 G33465 (.A1(W519), .A2(W7311), .ZN(W11581));
  NANDX1 G33466 (.A1(W9730), .A2(W2848), .ZN(O2308));
  NANDX1 G33467 (.A1(I1406), .A2(I1260), .ZN(W2504));
  NANDX1 G33468 (.A1(W1769), .A2(W20481), .ZN(W21681));
  NANDX1 G33469 (.A1(W15195), .A2(W17014), .ZN(W25000));
  NANDX1 G33470 (.A1(W7028), .A2(W5411), .ZN(W9262));
  NANDX1 G33471 (.A1(W11874), .A2(W7078), .ZN(W11902));
  NANDX1 G33472 (.A1(W15174), .A2(W21110), .ZN(W21684));
  NANDX1 G33473 (.A1(I137), .A2(I635), .ZN(W2085));
  NANDX1 G33474 (.A1(W1590), .A2(W1119), .ZN(W2086));
  NANDX1 G33475 (.A1(I480), .A2(W114), .ZN(W2509));
  NANDX1 G33476 (.A1(W21242), .A2(W10911), .ZN(W21689));
  NANDX1 G33477 (.A1(W15560), .A2(W14007), .ZN(W21693));
  NANDX1 G33478 (.A1(W2306), .A2(I1286), .ZN(W2494));
  NANDX1 G33479 (.A1(W4382), .A2(W7874), .ZN(O3265));
  NANDX1 G33480 (.A1(W2066), .A2(I1134), .ZN(W2099));
  NANDX1 G33481 (.A1(I1996), .A2(W9548), .ZN(W21705));
  NANDX1 G33482 (.A1(W9797), .A2(W6123), .ZN(W21708));
  NANDX1 G33483 (.A1(W778), .A2(W12423), .ZN(W22296));
  NANDX1 G33484 (.A1(W18240), .A2(W7829), .ZN(W21709));
  NANDX1 G33485 (.A1(W8837), .A2(W571), .ZN(W22295));
  NANDX1 G33486 (.A1(W2476), .A2(I638), .ZN(W2499));
  NANDX1 G33487 (.A1(W173), .A2(W676), .ZN(W2498));
  NANDX1 G33488 (.A1(W19051), .A2(W18274), .ZN(W21714));
  NANDX1 G33489 (.A1(W3871), .A2(W5926), .ZN(W9077));
  NANDX1 G33490 (.A1(W4109), .A2(I100), .ZN(W21704));
  NANDX1 G33491 (.A1(W200), .A2(W7509), .ZN(W11684));
  NANDX1 G33492 (.A1(I1068), .A2(W9050), .ZN(W11899));
  NANDX1 G33493 (.A1(W7569), .A2(W8917), .ZN(W10368));
  NANDX1 G33494 (.A1(W335), .A2(W2334), .ZN(W2492));
  NANDX1 G33495 (.A1(I619), .A2(I1087), .ZN(W2491));
  NANDX1 G33496 (.A1(I1648), .A2(W874), .ZN(W2490));
  NANDX1 G33497 (.A1(W879), .A2(W1861), .ZN(W22104));
  NANDX1 G33498 (.A1(W7666), .A2(W3089), .ZN(W10078));
  NANDX1 G33499 (.A1(W17326), .A2(W15179), .ZN(O2317));
  NANDX1 G33500 (.A1(W1355), .A2(I691), .ZN(W2103));
  NANDX1 G33501 (.A1(W1940), .A2(W953), .ZN(W2090));
  NANDX1 G33502 (.A1(W543), .A2(W1402), .ZN(W2502));
  NANDX1 G33503 (.A1(W14130), .A2(W5611), .ZN(W21699));
  NANDX1 G33504 (.A1(I1939), .A2(W15595), .ZN(W22301));
  NANDX1 G33505 (.A1(W1984), .A2(W299), .ZN(W2089));
  NANDX1 G33506 (.A1(I695), .A2(W1952), .ZN(W2501));
  NANDX1 G33507 (.A1(I450), .A2(I451), .ZN(W225));
  NANDX1 G33508 (.A1(W8624), .A2(W22027), .ZN(O3217));
  NANDX1 G33509 (.A1(W12486), .A2(W9641), .ZN(W22300));
  NANDX1 G33510 (.A1(I394), .A2(W2089), .ZN(W2500));
  NANDX1 G33511 (.A1(W11192), .A2(W11149), .ZN(O2471));
  NANDX1 G33512 (.A1(W447), .A2(W6198), .ZN(O384));
  NANDX1 G33513 (.A1(W4681), .A2(W1089), .ZN(W9084));
  NANDX1 G33514 (.A1(W12707), .A2(W21093), .ZN(W22106));
  NANDX1 G33515 (.A1(W1861), .A2(W3855), .ZN(W11688));
  NANDX1 G33516 (.A1(W6755), .A2(W1584), .ZN(W10079));
  NANDX1 G33517 (.A1(W82), .A2(I691), .ZN(W2094));
  NANDX1 G33518 (.A1(W17826), .A2(W18364), .ZN(O3195));
  NANDX1 G33519 (.A1(W11033), .A2(W3745), .ZN(W11685));
  NANDX1 G33520 (.A1(W4137), .A2(W137), .ZN(W9075));
  NANDX1 G33521 (.A1(W5020), .A2(W2904), .ZN(W9259));
  NANDX1 G33522 (.A1(I656), .A2(I657), .ZN(W328));
  NANDX1 G33523 (.A1(I1214), .A2(W19321), .ZN(W21703));
  NANDX1 G33524 (.A1(W8843), .A2(W4376), .ZN(W10429));
  NANDX1 G33525 (.A1(W487), .A2(W2413), .ZN(W9107));
  NANDX1 G33526 (.A1(W3948), .A2(W3648), .ZN(W22244));
  NANDX1 G33527 (.A1(I543), .A2(I370), .ZN(W2414));
  NANDX1 G33528 (.A1(W8216), .A2(W2298), .ZN(W9109));
  NANDX1 G33529 (.A1(I925), .A2(W460), .ZN(W10386));
  NANDX1 G33530 (.A1(I502), .A2(I503), .ZN(W251));
  NANDX1 G33531 (.A1(W22), .A2(W1605), .ZN(W2254));
  NANDX1 G33532 (.A1(W7659), .A2(I1686), .ZN(W9195));
  NANDX1 G33533 (.A1(W8110), .A2(W8144), .ZN(W9239));
  NANDX1 G33534 (.A1(W18580), .A2(W17582), .ZN(W24951));
  NANDX1 G33535 (.A1(W248), .A2(W20378), .ZN(W22242));
  NANDX1 G33536 (.A1(W7826), .A2(W10439), .ZN(W11836));
  NANDX1 G33537 (.A1(W16633), .A2(W17537), .ZN(W21832));
  NANDX1 G33538 (.A1(W8195), .A2(W14363), .ZN(W22239));
  NANDX1 G33539 (.A1(I1059), .A2(W1560), .ZN(W2227));
  NANDX1 G33540 (.A1(I1442), .A2(W990), .ZN(W9238));
  NANDX1 G33541 (.A1(W8147), .A2(W16928), .ZN(W22238));
  NANDX1 G33542 (.A1(W13873), .A2(W11742), .ZN(W24809));
  NANDX1 G33543 (.A1(I504), .A2(I505), .ZN(W252));
  NANDX1 G33544 (.A1(I220), .A2(W2128), .ZN(W2409));
  NANDX1 G33545 (.A1(W5657), .A2(W9724), .ZN(W10067));
  NANDX1 G33546 (.A1(W19072), .A2(W4400), .ZN(W21834));
  NANDX1 G33547 (.A1(W3759), .A2(W10250), .ZN(W11842));
  NANDX1 G33548 (.A1(I1703), .A2(W11273), .ZN(W11608));
  NANDX1 G33549 (.A1(W5390), .A2(I384), .ZN(W22248));
  NANDX1 G33550 (.A1(I498), .A2(I499), .ZN(W249));
  NANDX1 G33551 (.A1(W6865), .A2(W4999), .ZN(W11844));
  NANDX1 G33552 (.A1(I500), .A2(I501), .ZN(W250));
  NANDX1 G33553 (.A1(W8374), .A2(W12611), .ZN(O2338));
  NANDX1 G33554 (.A1(W11342), .A2(W13380), .ZN(O2462));
  NANDX1 G33555 (.A1(W1920), .A2(W13496), .ZN(W22129));
  NANDX1 G33556 (.A1(W8672), .A2(W9246), .ZN(O3254));
  NANDX1 G33557 (.A1(W9288), .A2(W11755), .ZN(W22247));
  NANDX1 G33558 (.A1(W847), .A2(I734), .ZN(W2422));
  NANDX1 G33559 (.A1(W19090), .A2(W19140), .ZN(W24811));
  NANDX1 G33560 (.A1(I328), .A2(W2286), .ZN(W2421));
  NANDX1 G33561 (.A1(W7252), .A2(W8847), .ZN(W9105));
  NANDX1 G33562 (.A1(W9316), .A2(W15437), .ZN(W21817));
  NANDX1 G33563 (.A1(I445), .A2(W767), .ZN(W2142));
  NANDX1 G33564 (.A1(W10480), .A2(I1326), .ZN(W11838));
  NANDX1 G33565 (.A1(W21265), .A2(W19), .ZN(O2344));
  NANDX1 G33566 (.A1(I1520), .A2(W18924), .ZN(O2345));
  NANDX1 G33567 (.A1(W533), .A2(W6823), .ZN(W21822));
  NANDX1 G33568 (.A1(W4179), .A2(W1169), .ZN(W21824));
  NANDX1 G33569 (.A1(W18501), .A2(W8480), .ZN(W21826));
  NANDX1 G33570 (.A1(W1725), .A2(W1965), .ZN(W2400));
  NANDX1 G33571 (.A1(W2840), .A2(W6989), .ZN(W21844));
  NANDX1 G33572 (.A1(I508), .A2(I509), .ZN(W254));
  NANDX1 G33573 (.A1(W1998), .A2(W6296), .ZN(O2351));
  NANDX1 G33574 (.A1(W2024), .A2(I741), .ZN(W2256));
  NANDX1 G33575 (.A1(W4038), .A2(W3769), .ZN(W22232));
  NANDX1 G33576 (.A1(W20770), .A2(W21193), .ZN(W22133));
  NANDX1 G33577 (.A1(W175), .A2(I1798), .ZN(W2401));
  NANDX1 G33578 (.A1(W19273), .A2(W2138), .ZN(O2456));
  NANDX1 G33579 (.A1(W19030), .A2(I1162), .ZN(W22083));
  NANDX1 G33580 (.A1(I444), .A2(W506), .ZN(W2152));
  NANDX1 G33581 (.A1(W6964), .A2(W6428), .ZN(W11672));
  NANDX1 G33582 (.A1(W1262), .A2(W2454), .ZN(O3252));
  NANDX1 G33583 (.A1(W1060), .A2(I1831), .ZN(W2399));
  NANDX1 G33584 (.A1(W22129), .A2(W12922), .ZN(W24815));
  NANDX1 G33585 (.A1(W16610), .A2(W6892), .ZN(W21850));
  NANDX1 G33586 (.A1(W6253), .A2(W2270), .ZN(W10423));
  NANDX1 G33587 (.A1(W11752), .A2(W7648), .ZN(O3249));
  NANDX1 G33588 (.A1(W5830), .A2(W6928), .ZN(W11611));
  NANDX1 G33589 (.A1(W17162), .A2(W13615), .ZN(W22227));
  NANDX1 G33590 (.A1(W13917), .A2(W20351), .ZN(W21851));
  NANDX1 G33591 (.A1(I368), .A2(I226), .ZN(W2398));
  NANDX1 G33592 (.A1(W19113), .A2(W3410), .ZN(O2454));
  NANDX1 G33593 (.A1(W10484), .A2(W11339), .ZN(W11674));
  NANDX1 G33594 (.A1(W11514), .A2(W5449), .ZN(W11691));
  NANDX1 G33595 (.A1(W11533), .A2(I708), .ZN(W22131));
  NANDX1 G33596 (.A1(W428), .A2(W7504), .ZN(W11823));
  NANDX1 G33597 (.A1(I734), .A2(I735), .ZN(W367));
  NANDX1 G33598 (.A1(W605), .A2(W23732), .ZN(W24812));
  NANDX1 G33599 (.A1(W1281), .A2(W17565), .ZN(O2347));
  NANDX1 G33600 (.A1(W20419), .A2(W9354), .ZN(O2421));
  NANDX1 G33601 (.A1(W15241), .A2(W9456), .ZN(W24862));
  NANDX1 G33602 (.A1(I1307), .A2(I1503), .ZN(W2147));
  NANDX1 G33603 (.A1(W4141), .A2(W5051), .ZN(W9235));
  NANDX1 G33604 (.A1(W18240), .A2(W1983), .ZN(O2348));
  NANDX1 G33605 (.A1(W11586), .A2(W129), .ZN(W22127));
  NANDX1 G33606 (.A1(W10852), .A2(I1894), .ZN(W22085));
  NANDX1 G33607 (.A1(W124), .A2(W633), .ZN(W2148));
  NANDX1 G33608 (.A1(W10131), .A2(W1209), .ZN(O3220));
  NANDX1 G33609 (.A1(I506), .A2(I507), .ZN(W253));
  NANDX1 G33610 (.A1(W5263), .A2(W1009), .ZN(W11610));
  NANDX1 G33611 (.A1(W7806), .A2(W550), .ZN(W11820));
  NANDX1 G33612 (.A1(I992), .A2(W7879), .ZN(W11816));
  NANDX1 G33613 (.A1(W297), .A2(W90), .ZN(W2402));
  NANDX1 G33614 (.A1(I603), .A2(W10941), .ZN(W11815));
  NANDX1 G33615 (.A1(W2415), .A2(W1329), .ZN(W11814));
  NANDX1 G33616 (.A1(W2295), .A2(W18697), .ZN(W24805));
  NANDX1 G33617 (.A1(W6686), .A2(W4777), .ZN(W22264));
  NANDX1 G33618 (.A1(W1168), .A2(W1310), .ZN(W2449));
  NANDX1 G33619 (.A1(W3227), .A2(W907), .ZN(W10382));
  NANDX1 G33620 (.A1(I1290), .A2(W6379), .ZN(W9089));
  NANDX1 G33621 (.A1(W7562), .A2(W6310), .ZN(O2422));
  NANDX1 G33622 (.A1(I1457), .A2(W535), .ZN(W2447));
  NANDX1 G33623 (.A1(I1864), .A2(W1068), .ZN(W11859));
  NANDX1 G33624 (.A1(I1156), .A2(W15133), .ZN(W24965));
  NANDX1 G33625 (.A1(W16936), .A2(W13470), .ZN(W22263));
  NANDX1 G33626 (.A1(I478), .A2(I479), .ZN(W239));
  NANDX1 G33627 (.A1(W5397), .A2(I443), .ZN(O3214));
  NANDX1 G33628 (.A1(W2771), .A2(W5704), .ZN(W11861));
  NANDX1 G33629 (.A1(W2622), .A2(W4142), .ZN(O2331));
  NANDX1 G33630 (.A1(W482), .A2(W1206), .ZN(W2131));
  NANDX1 G33631 (.A1(W455), .A2(W9693), .ZN(W21785));
  NANDX1 G33632 (.A1(W10328), .A2(W11441), .ZN(O524));
  NANDX1 G33633 (.A1(W9660), .A2(W5656), .ZN(W10071));
  NANDX1 G33634 (.A1(I740), .A2(I741), .ZN(W370));
  NANDX1 G33635 (.A1(W5439), .A2(W5612), .ZN(W22089));
  NANDX1 G33636 (.A1(W8660), .A2(W2547), .ZN(W10383));
  NANDX1 G33637 (.A1(W7506), .A2(W6925), .ZN(W9093));
  NANDX1 G33638 (.A1(W3798), .A2(W3567), .ZN(W11854));
  NANDX1 G33639 (.A1(W2764), .A2(I794), .ZN(O3262));
  NANDX1 G33640 (.A1(W6139), .A2(I158), .ZN(W11599));
  NANDX1 G33641 (.A1(W2077), .A2(I84), .ZN(W2453));
  NANDX1 G33642 (.A1(I730), .A2(W2971), .ZN(W10441));
  NANDX1 G33643 (.A1(W18736), .A2(W10430), .ZN(W24803));
  NANDX1 G33644 (.A1(I476), .A2(I477), .ZN(W238));
  NANDX1 G33645 (.A1(W5563), .A2(W4718), .ZN(W10380));
  NANDX1 G33646 (.A1(W21187), .A2(W12999), .ZN(W21769));
  NANDX1 G33647 (.A1(W7999), .A2(W10897), .ZN(W22092));
  NANDX1 G33648 (.A1(W4529), .A2(W10236), .ZN(W11868));
  NANDX1 G33649 (.A1(W11364), .A2(W7641), .ZN(W21772));
  NANDX1 G33650 (.A1(I482), .A2(I483), .ZN(W241));
  NANDX1 G33651 (.A1(I742), .A2(I743), .ZN(W371));
  NANDX1 G33652 (.A1(W18199), .A2(W8021), .ZN(W22091));
  NANDX1 G33653 (.A1(I693), .A2(W5431), .ZN(O3261));
  NANDX1 G33654 (.A1(W9930), .A2(W7458), .ZN(W11600));
  NANDX1 G33655 (.A1(W1628), .A2(W9760), .ZN(W21774));
  NANDX1 G33656 (.A1(W775), .A2(W9986), .ZN(W11865));
  NANDX1 G33657 (.A1(W5771), .A2(I1388), .ZN(W10381));
  NANDX1 G33658 (.A1(W2233), .A2(W871), .ZN(W11602));
  NANDX1 G33659 (.A1(I1760), .A2(W784), .ZN(W2130));
  NANDX1 G33660 (.A1(I642), .A2(I643), .ZN(W321));
  NANDX1 G33661 (.A1(W16481), .A2(W14229), .ZN(W21797));
  NANDX1 G33662 (.A1(W5999), .A2(W7076), .ZN(W11604));
  NANDX1 G33663 (.A1(W394), .A2(W2347), .ZN(W2433));
  NANDX1 G33664 (.A1(I308), .A2(W14752), .ZN(W21793));
  NANDX1 G33665 (.A1(W697), .A2(I200), .ZN(W2441));
  NANDX1 G33666 (.A1(W17458), .A2(W1956), .ZN(O2335));
  NANDX1 G33667 (.A1(W2587), .A2(W7195), .ZN(W9094));
  NANDX1 G33668 (.A1(W1624), .A2(W1788), .ZN(W2136));
  NANDX1 G33669 (.A1(W1355), .A2(W4575), .ZN(W11605));
  NANDX1 G33670 (.A1(W1415), .A2(W3606), .ZN(O359));
  NANDX1 G33671 (.A1(W15266), .A2(W7984), .ZN(W24959));
  NANDX1 G33672 (.A1(W6034), .A2(W19677), .ZN(W21796));
  NANDX1 G33673 (.A1(W1490), .A2(W1159), .ZN(W2135));
  NANDX1 G33674 (.A1(W13571), .A2(W15208), .ZN(W22252));
  NANDX1 G33675 (.A1(W510), .A2(W4594), .ZN(W11851));
  NANDX1 G33676 (.A1(W4154), .A2(W16037), .ZN(W22251));
  NANDX1 G33677 (.A1(W9803), .A2(W19083), .ZN(W21799));
  NANDX1 G33678 (.A1(W9833), .A2(W15176), .ZN(W24958));
  NANDX1 G33679 (.A1(W165), .A2(I582), .ZN(W9188));
  NANDX1 G33680 (.A1(W967), .A2(W7548), .ZN(W11850));
  NANDX1 G33681 (.A1(W783), .A2(W3375), .ZN(W11848));
  NANDX1 G33682 (.A1(W10139), .A2(W8596), .ZN(W11847));
  NANDX1 G33683 (.A1(I490), .A2(I491), .ZN(W245));
  NANDX1 G33684 (.A1(W2908), .A2(W74), .ZN(W10385));
  NANDX1 G33685 (.A1(I488), .A2(I489), .ZN(W244));
  NANDX1 G33686 (.A1(W41), .A2(I1748), .ZN(W2438));
  NANDX1 G33687 (.A1(W765), .A2(W1406), .ZN(W2440));
  NANDX1 G33688 (.A1(W10164), .A2(W2323), .ZN(O3257));
  NANDX1 G33689 (.A1(W11414), .A2(W16883), .ZN(W21789));
  NANDX1 G33690 (.A1(W5753), .A2(W1088), .ZN(W22259));
  NANDX1 G33691 (.A1(W4006), .A2(W21566), .ZN(W24807));
  NANDX1 G33692 (.A1(W3723), .A2(W13196), .ZN(W24961));
  NANDX1 G33693 (.A1(I16), .A2(I256), .ZN(W2133));
  NANDX1 G33694 (.A1(I637), .A2(W1703), .ZN(O2334));
  INVX1 G33695 (.I(W38412), .ZN(O11192));
  INVX1 G33696 (.I(W30910), .ZN(W43882));
  INVX1 G33697 (.I(W8108), .ZN(W10159));
  INVX1 G33698 (.I(W863), .ZN(W40902));
  INVX1 G33699 (.I(W31402), .ZN(O13461));
  INVX1 G33700 (.I(W2350), .ZN(O11227));
  INVX1 G33701 (.I(I1393), .ZN(W10155));
  INVX1 G33702 (.I(W2683), .ZN(W40712));
  INVX1 G33703 (.I(W1224), .ZN(W7396));
  INVX1 G33704 (.I(W3021), .ZN(O368));
  INVX1 G33705 (.I(W16015), .ZN(O13460));
  INVX1 G33706 (.I(I1850), .ZN(W7389));
  INVX1 G33707 (.I(W31351), .ZN(O11193));
  INVX1 G33708 (.I(I1136), .ZN(W7006));
  INVX1 G33709 (.I(W22364), .ZN(O13300));
  INVX1 G33710 (.I(W17291), .ZN(O11319));
  INVX1 G33711 (.I(W23322), .ZN(O13299));
  INVX1 G33712 (.I(W22634), .ZN(O13301));
  INVX1 G33713 (.I(W22834), .ZN(O13169));
  INVX1 G33714 (.I(W12914), .ZN(W41036));
  INVX1 G33715 (.I(I1091), .ZN(O11103));
  INVX1 G33716 (.I(W29366), .ZN(O13171));
  INVX1 G33717 (.I(W13148), .ZN(O11226));
  INVX1 G33718 (.I(W1776), .ZN(O13173));
  INVX1 G33719 (.I(W6646), .ZN(W9869));
  INVX1 G33720 (.I(W2377), .ZN(W7174));
  INVX1 G33721 (.I(W5650), .ZN(W7395));
  INVX1 G33722 (.I(W15458), .ZN(O11106));
  INVX1 G33723 (.I(W3752), .ZN(W9874));
  INVX1 G33724 (.I(W4416), .ZN(W9870));
  INVX1 G33725 (.I(W8656), .ZN(W41069));
  INVX1 G33726 (.I(W3515), .ZN(W7423));
  INVX1 G33727 (.I(W10090), .ZN(W10180));
  INVX1 G33728 (.I(W19906), .ZN(O11341));
  INVX1 G33729 (.I(W27137), .ZN(O11215));
  INVX1 G33730 (.I(W10219), .ZN(O13322));
  INVX1 G33731 (.I(W196), .ZN(W9832));
  INVX1 G33732 (.I(W39952), .ZN(O13310));
  INVX1 G33733 (.I(W2902), .ZN(W10023));
  INVX1 G33734 (.I(W1843), .ZN(W9831));
  INVX1 G33735 (.I(W7473), .ZN(W10179));
  INVX1 G33736 (.I(W1698), .ZN(W10014));
  INVX1 G33737 (.I(W29938), .ZN(O11213));
  INVX1 G33738 (.I(W37469), .ZN(O13151));
  INVX1 G33739 (.I(W3276), .ZN(W7425));
  INVX1 G33740 (.I(W8988), .ZN(W10181));
  INVX1 G33741 (.I(W14594), .ZN(W40881));
  INVX1 G33742 (.I(I1531), .ZN(W7199));
  INVX1 G33743 (.I(I975), .ZN(O13321));
  INVX1 G33744 (.I(W4690), .ZN(W10178));
  INVX1 G33745 (.I(W31629), .ZN(O11337));
  INVX1 G33746 (.I(W321), .ZN(W9835));
  INVX1 G33747 (.I(I937), .ZN(W7418));
  INVX1 G33748 (.I(W19376), .ZN(O11087));
  INVX1 G33749 (.I(I1265), .ZN(W7203));
  INVX1 G33750 (.I(W1782), .ZN(O170));
  INVX1 G33751 (.I(W34404), .ZN(O11339));
  INVX1 G33752 (.I(W4554), .ZN(W7419));
  INVX1 G33753 (.I(W3642), .ZN(W6993));
  INVX1 G33754 (.I(W39225), .ZN(O11082));
  INVX1 G33755 (.I(I1908), .ZN(W9834));
  INVX1 G33756 (.I(W3694), .ZN(W10011));
  INVX1 G33757 (.I(W9684), .ZN(W43477));
  INVX1 G33758 (.I(W9544), .ZN(W9833));
  INVX1 G33759 (.I(W4875), .ZN(W7422));
  INVX1 G33760 (.I(W6952), .ZN(W6992));
  INVX1 G33761 (.I(W31815), .ZN(O11202));
  INVX1 G33762 (.I(W26911), .ZN(W40704));
  INVX1 G33763 (.I(W1485), .ZN(W7430));
  INVX1 G33764 (.I(W13771), .ZN(O11206));
  INVX1 G33765 (.I(W30407), .ZN(W43914));
  INVX1 G33766 (.I(W11261), .ZN(O11208));
  INVX1 G33767 (.I(I160), .ZN(W7429));
  INVX1 G33768 (.I(W92), .ZN(W10022));
  INVX1 G33769 (.I(W1349), .ZN(W7187));
  INVX1 G33770 (.I(W3023), .ZN(O13485));
  INVX1 G33771 (.I(I1792), .ZN(W7188));
  INVX1 G33772 (.I(W35069), .ZN(O11078));
  INVX1 G33773 (.I(W38386), .ZN(O13484));
  INVX1 G33774 (.I(W1633), .ZN(O13143));
  INVX1 G33775 (.I(W5603), .ZN(W10020));
  INVX1 G33776 (.I(W4028), .ZN(W7190));
  INVX1 G33777 (.I(W1900), .ZN(O11346));
  INVX1 G33778 (.I(W8222), .ZN(W10185));
  INVX1 G33779 (.I(W1635), .ZN(W10187));
  INVX1 G33780 (.I(W6969), .ZN(W40875));
  INVX1 G33781 (.I(W5798), .ZN(O11076));
  INVX1 G33782 (.I(W5942), .ZN(W7196));
  INVX1 G33783 (.I(W40336), .ZN(O13481));
  INVX1 G33784 (.I(I1281), .ZN(O11204));
  INVX1 G33785 (.I(W16195), .ZN(W43910));
  INVX1 G33786 (.I(W24168), .ZN(O13482));
  INVX1 G33787 (.I(W17535), .ZN(O13148));
  INVX1 G33788 (.I(W33846), .ZN(O11211));
  INVX1 G33789 (.I(W28510), .ZN(O13320));
  INVX1 G33790 (.I(W22607), .ZN(O11080));
  INVX1 G33791 (.I(W32340), .ZN(O13311));
  INVX1 G33792 (.I(W23778), .ZN(O11216));
  INVX1 G33793 (.I(I1078), .ZN(W40696));
  INVX1 G33794 (.I(W26865), .ZN(W40871));
  INVX1 G33795 (.I(I1889), .ZN(O13146));
  INVX1 G33796 (.I(W19673), .ZN(O11205));
  INVX1 G33797 (.I(W7863), .ZN(W10017));
  INVX1 G33798 (.I(W19622), .ZN(O13145));
  INVX1 G33799 (.I(I886), .ZN(W7195));
  INVX1 G33800 (.I(W4379), .ZN(W7194));
  INVX1 G33801 (.I(W5247), .ZN(W10031));
  INVX1 G33802 (.I(W9002), .ZN(O11223));
  INVX1 G33803 (.I(W37516), .ZN(O13328));
  INVX1 G33804 (.I(W25625), .ZN(O13466));
  INVX1 G33805 (.I(W4502), .ZN(W7001));
  INVX1 G33806 (.I(W4799), .ZN(W7213));
  INVX1 G33807 (.I(W22972), .ZN(O13468));
  INVX1 G33808 (.I(W5326), .ZN(O13304));
  INVX1 G33809 (.I(W3359), .ZN(W9853));
  INVX1 G33810 (.I(I793), .ZN(W7000));
  INVX1 G33811 (.I(W39040), .ZN(O13465));
  INVX1 G33812 (.I(I479), .ZN(O11097));
  INVX1 G33813 (.I(W1957), .ZN(W7405));
  INVX1 G33814 (.I(W26838), .ZN(W43488));
  INVX1 G33815 (.I(W15834), .ZN(O11096));
  INVX1 G33816 (.I(W4123), .ZN(W6999));
  INVX1 G33817 (.I(W9748), .ZN(O351));
  INVX1 G33818 (.I(W14912), .ZN(W40720));
  INVX1 G33819 (.I(W41026), .ZN(W43896));
  INVX1 G33820 (.I(W21175), .ZN(O13330));
  INVX1 G33821 (.I(W5429), .ZN(W10001));
  INVX1 G33822 (.I(I398), .ZN(W10035));
  INVX1 G33823 (.I(W6771), .ZN(W7216));
  INVX1 G33824 (.I(I1140), .ZN(O180));
  INVX1 G33825 (.I(W1749), .ZN(W7177));
  INVX1 G33826 (.I(W9117), .ZN(W43886));
  INVX1 G33827 (.I(W38223), .ZN(O13303));
  INVX1 G33828 (.I(W4913), .ZN(W7004));
  INVX1 G33829 (.I(W7352), .ZN(W9867));
  INVX1 G33830 (.I(W9673), .ZN(W9849));
  INVX1 G33831 (.I(W305), .ZN(W7178));
  INVX1 G33832 (.I(W17077), .ZN(O13167));
  INVX1 G33833 (.I(W4842), .ZN(W9864));
  INVX1 G33834 (.I(W4738), .ZN(W7399));
  INVX1 G33835 (.I(W5081), .ZN(O11224));
  INVX1 G33836 (.I(W1154), .ZN(W9858));
  INVX1 G33837 (.I(W19994), .ZN(O13464));
  INVX1 G33838 (.I(W18892), .ZN(O11327));
  INVX1 G33839 (.I(W4834), .ZN(O13308));
  INVX1 G33840 (.I(W8103), .ZN(W9845));
  INVX1 G33841 (.I(W9218), .ZN(W10133));
  INVX1 G33842 (.I(I1616), .ZN(W41058));
  INVX1 G33843 (.I(W32473), .ZN(O13473));
  INVX1 G33844 (.I(W22815), .ZN(O13307));
  INVX1 G33845 (.I(W25727), .ZN(O11335));
  INVX1 G33846 (.I(W24622), .ZN(O13474));
  INVX1 G33847 (.I(W30670), .ZN(W40709));
  INVX1 G33848 (.I(W1334), .ZN(W7184));
  INVX1 G33849 (.I(W36539), .ZN(W40864));
  INVX1 G33850 (.I(W40156), .ZN(W43482));
  INVX1 G33851 (.I(W7632), .ZN(W10176));
  INVX1 G33852 (.I(W6456), .ZN(W43709));
  INVX1 G33853 (.I(W19047), .ZN(W43903));
  INVX1 G33854 (.I(W14935), .ZN(O11218));
  INVX1 G33855 (.I(I1608), .ZN(W7417));
  INVX1 G33856 (.I(I1332), .ZN(W6994));
  INVX1 G33857 (.I(W536), .ZN(W10009));
  INVX1 G33858 (.I(W835), .ZN(W6997));
  INVX1 G33859 (.I(W1094), .ZN(W7180));
  INVX1 G33860 (.I(W1702), .ZN(W7209));
  INVX1 G33861 (.I(W23536), .ZN(O11095));
  INVX1 G33862 (.I(W34302), .ZN(W40718));
  INVX1 G33863 (.I(I714), .ZN(W10030));
  INVX1 G33864 (.I(W4056), .ZN(W10029));
  INVX1 G33865 (.I(W2972), .ZN(O11199));
  INVX1 G33866 (.I(W28705), .ZN(W43685));
  INVX1 G33867 (.I(W11631), .ZN(O11100));
  INVX1 G33868 (.I(W1760), .ZN(W7412));
  INVX1 G33869 (.I(W619), .ZN(W7206));
  INVX1 G33870 (.I(I693), .ZN(W10028));
  INVX1 G33871 (.I(W1722), .ZN(W7204));
  INVX1 G33872 (.I(W20206), .ZN(W43898));
  INVX1 G33873 (.I(W3307), .ZN(W6996));
  INVX1 G33874 (.I(I1862), .ZN(W10171));
  INVX1 G33875 (.I(W2412), .ZN(W10172));
  INVX1 G33876 (.I(W5772), .ZN(W7323));
  INVX1 G33877 (.I(W44), .ZN(W7127));
  INVX1 G33878 (.I(W35876), .ZN(W40991));
  INVX1 G33879 (.I(W8080), .ZN(W10100));
  INVX1 G33880 (.I(W36336), .ZN(O13268));
  INVX1 G33881 (.I(W37712), .ZN(O11259));
  INVX1 G33882 (.I(W4772), .ZN(O13411));
  INVX1 G33883 (.I(W7226), .ZN(W10104));
  INVX1 G33884 (.I(I1915), .ZN(W7066));
  INVX1 G33885 (.I(W16853), .ZN(O13270));
  INVX1 G33886 (.I(W369), .ZN(W10108));
  INVX1 G33887 (.I(W410), .ZN(W7128));
  INVX1 G33888 (.I(W18968), .ZN(O13413));
  INVX1 G33889 (.I(I950), .ZN(W7126));
  INVX1 G33890 (.I(W5922), .ZN(W7064));
  INVX1 G33891 (.I(W7758), .ZN(W10109));
  INVX1 G33892 (.I(W41216), .ZN(O13225));
  INVX1 G33893 (.I(W19347), .ZN(O11257));
  INVX1 G33894 (.I(W10011), .ZN(W10111));
  INVX1 G33895 (.I(W6678), .ZN(W7063));
  INVX1 G33896 (.I(W21043), .ZN(O13271));
  INVX1 G33897 (.I(W4526), .ZN(W7130));
  INVX1 G33898 (.I(W5263), .ZN(W10113));
  INVX1 G33899 (.I(W6571), .ZN(W7271));
  INVX1 G33900 (.I(W5455), .ZN(W7268));
  INVX1 G33901 (.I(W3510), .ZN(O173));
  INVX1 G33902 (.I(W22883), .ZN(O11260));
  INVX1 G33903 (.I(W11521), .ZN(O11147));
  INVX1 G33904 (.I(W23913), .ZN(O13375));
  INVX1 G33905 (.I(W3329), .ZN(W7117));
  INVX1 G33906 (.I(W7410), .ZN(W43579));
  INVX1 G33907 (.I(W20902), .ZN(W40789));
  INVX1 G33908 (.I(W2077), .ZN(O345));
  INVX1 G33909 (.I(W20055), .ZN(W40788));
  INVX1 G33910 (.I(W8572), .ZN(W10095));
  INVX1 G33911 (.I(W40079), .ZN(O11261));
  INVX1 G33912 (.I(W14976), .ZN(W40785));
  INVX1 G33913 (.I(W47), .ZN(W7279));
  INVX1 G33914 (.I(W31939), .ZN(O13231));
  INVX1 G33915 (.I(I609), .ZN(W7328));
  INVX1 G33916 (.I(I772), .ZN(W7121));
  INVX1 G33917 (.I(W27783), .ZN(W40988));
  INVX1 G33918 (.I(W40798), .ZN(O13371));
  INVX1 G33919 (.I(W2481), .ZN(W7319));
  INVX1 G33920 (.I(W6193), .ZN(W7274));
  INVX1 G33921 (.I(W3092), .ZN(W7321));
  INVX1 G33922 (.I(W1016), .ZN(W9926));
  INVX1 G33923 (.I(W17410), .ZN(O13369));
  INVX1 G33924 (.I(I426), .ZN(O166));
  INVX1 G33925 (.I(W6942), .ZN(W7322));
  INVX1 G33926 (.I(W33551), .ZN(O13410));
  INVX1 G33927 (.I(W643), .ZN(W40936));
  INVX1 G33928 (.I(I1386), .ZN(W7335));
  INVX1 G33929 (.I(W3739), .ZN(W10062));
  INVX1 G33930 (.I(W4061), .ZN(W40995));
  INVX1 G33931 (.I(W43311), .ZN(O13217));
  INVX1 G33932 (.I(W8722), .ZN(W10117));
  INVX1 G33933 (.I(W1575), .ZN(W7337));
  INVX1 G33934 (.I(W2979), .ZN(W7058));
  INVX1 G33935 (.I(W6731), .ZN(W7258));
  INVX1 G33936 (.I(W18464), .ZN(W40938));
  INVX1 G33937 (.I(W24668), .ZN(O11253));
  INVX1 G33938 (.I(W10750), .ZN(O13214));
  INVX1 G33939 (.I(W20264), .ZN(W43831));
  INVX1 G33940 (.I(W2940), .ZN(O177));
  INVX1 G33941 (.I(W4915), .ZN(O164));
  INVX1 G33942 (.I(W33591), .ZN(O11167));
  INVX1 G33943 (.I(W12406), .ZN(W40768));
  INVX1 G33944 (.I(W9665), .ZN(W9922));
  INVX1 G33945 (.I(W5051), .ZN(W7251));
  INVX1 G33946 (.I(W3012), .ZN(W7138));
  INVX1 G33947 (.I(W24644), .ZN(O11297));
  INVX1 G33948 (.I(I531), .ZN(W7249));
  INVX1 G33949 (.I(W26513), .ZN(W43644));
  INVX1 G33950 (.I(W4275), .ZN(W43835));
  INVX1 G33951 (.I(W38922), .ZN(O11133));
  INVX1 G33952 (.I(W1998), .ZN(W9918));
  INVX1 G33953 (.I(I262), .ZN(W7263));
  INVX1 G33954 (.I(W5726), .ZN(W7061));
  INVX1 G33955 (.I(W26532), .ZN(O13273));
  INVX1 G33956 (.I(W17020), .ZN(O13363));
  INVX1 G33957 (.I(W2291), .ZN(W10065));
  INVX1 G33958 (.I(W6196), .ZN(W7330));
  INVX1 G33959 (.I(W12846), .ZN(O13416));
  INVX1 G33960 (.I(W12303), .ZN(O11294));
  INVX1 G33961 (.I(W34395), .ZN(O11137));
  INVX1 G33962 (.I(W29484), .ZN(O11136));
  INVX1 G33963 (.I(W1742), .ZN(W43633));
  INVX1 G33964 (.I(W448), .ZN(W7265));
  INVX1 G33965 (.I(W2405), .ZN(W7132));
  INVX1 G33966 (.I(W39415), .ZN(O11263));
  INVX1 G33967 (.I(W2794), .ZN(O165));
  INVX1 G33968 (.I(W14760), .ZN(O13275));
  INVX1 G33969 (.I(W8741), .ZN(W9965));
  INVX1 G33970 (.I(W16521), .ZN(W43566));
  INVX1 G33971 (.I(W16110), .ZN(O13362));
  INVX1 G33972 (.I(W7093), .ZN(W9966));
  INVX1 G33973 (.I(W184), .ZN(W7331));
  INVX1 G33974 (.I(W20343), .ZN(W43638));
  INVX1 G33975 (.I(W23508), .ZN(O13220));
  INVX1 G33976 (.I(W38739), .ZN(O13419));
  INVX1 G33977 (.I(W2958), .ZN(W9968));
  INVX1 G33978 (.I(W2313), .ZN(W7092));
  INVX1 G33979 (.I(W25633), .ZN(W40805));
  INVX1 G33980 (.I(W30193), .ZN(O11156));
  INVX1 G33981 (.I(W36148), .ZN(W43611));
  INVX1 G33982 (.I(W2382), .ZN(W9952));
  INVX1 G33983 (.I(W10973), .ZN(O11279));
  INVX1 G33984 (.I(W12417), .ZN(O13396));
  INVX1 G33985 (.I(W38215), .ZN(O13248));
  INVX1 G33986 (.I(W36294), .ZN(W40956));
  INVX1 G33987 (.I(W10410), .ZN(O11155));
  INVX1 G33988 (.I(W6270), .ZN(W7295));
  INVX1 G33989 (.I(W5718), .ZN(W10080));
  INVX1 G33990 (.I(W14006), .ZN(O11153));
  INVX1 G33991 (.I(W31689), .ZN(O13249));
  INVX1 G33992 (.I(W4071), .ZN(W7101));
  INVX1 G33993 (.I(W23586), .ZN(O11158));
  INVX1 G33994 (.I(W866), .ZN(W7089));
  INVX1 G33995 (.I(W36842), .ZN(W43801));
  INVX1 G33996 (.I(W6754), .ZN(W7284));
  INVX1 G33997 (.I(W4685), .ZN(W7088));
  INVX1 G33998 (.I(W18657), .ZN(O13259));
  INVX1 G33999 (.I(W40271), .ZN(O11280));
  INVX1 G34000 (.I(W28990), .ZN(O11281));
  INVX1 G34001 (.I(W8741), .ZN(O13244));
  INVX1 G34002 (.I(W42981), .ZN(O13388));
  INVX1 G34003 (.I(W2218), .ZN(W9939));
  INVX1 G34004 (.I(W18590), .ZN(O11269));
  INVX1 G34005 (.I(W11804), .ZN(W43604));
  INVX1 G34006 (.I(I408), .ZN(O13251));
  INVX1 G34007 (.I(W3869), .ZN(W9949));
  INVX1 G34008 (.I(W4786), .ZN(O342));
  INVX1 G34009 (.I(W34303), .ZN(O11272));
  INVX1 G34010 (.I(I368), .ZN(W9943));
  INVX1 G34011 (.I(W1374), .ZN(W7095));
  INVX1 G34012 (.I(I873), .ZN(W7094));
  INVX1 G34013 (.I(W23160), .ZN(O11271));
  INVX1 G34014 (.I(W11384), .ZN(W43793));
  INVX1 G34015 (.I(W5407), .ZN(W9950));
  INVX1 G34016 (.I(W7050), .ZN(W7294));
  INVX1 G34017 (.I(W21121), .ZN(W40799));
  INVX1 G34018 (.I(I1729), .ZN(O11268));
  INVX1 G34019 (.I(I185), .ZN(O13252));
  INVX1 G34020 (.I(W11567), .ZN(W40806));
  INVX1 G34021 (.I(W9081), .ZN(W9951));
  INVX1 G34022 (.I(W5454), .ZN(W7098));
  INVX1 G34023 (.I(W33273), .ZN(O13250));
  INVX1 G34024 (.I(W1225), .ZN(O11276));
  INVX1 G34025 (.I(W10831), .ZN(O11277));
  INVX1 G34026 (.I(W1644), .ZN(W9942));
  INVX1 G34027 (.I(I44), .ZN(W7289));
  INVX1 G34028 (.I(I1796), .ZN(W9940));
  INVX1 G34029 (.I(W1418), .ZN(W7282));
  INVX1 G34030 (.I(W14240), .ZN(O11152));
  INVX1 G34031 (.I(W31438), .ZN(O13383));
  INVX1 G34032 (.I(W10), .ZN(W7079));
  INVX1 G34033 (.I(W2313), .ZN(W9935));
  INVX1 G34034 (.I(W14779), .ZN(O13235));
  INVX1 G34035 (.I(W4601), .ZN(W9961));
  INVX1 G34036 (.I(W8341), .ZN(O13382));
  INVX1 G34037 (.I(W9224), .ZN(W10092));
  INVX1 G34038 (.I(W7685), .ZN(W10093));
  INVX1 G34039 (.I(W3876), .ZN(O13407));
  INVX1 G34040 (.I(W28285), .ZN(O13381));
  INVX1 G34041 (.I(W4905), .ZN(W7077));
  INVX1 G34042 (.I(W6554), .ZN(W7080));
  INVX1 G34043 (.I(W6399), .ZN(W7310));
  INVX1 G34044 (.I(I990), .ZN(W7110));
  INVX1 G34045 (.I(W13613), .ZN(O13233));
  INVX1 G34046 (.I(W13941), .ZN(O13379));
  INVX1 G34047 (.I(W15599), .ZN(O11288));
  INVX1 G34048 (.I(W10523), .ZN(O13376));
  INVX1 G34049 (.I(W1821), .ZN(W7281));
  INVX1 G34050 (.I(W1446), .ZN(O176));
  INVX1 G34051 (.I(W4638), .ZN(W7076));
  INVX1 G34052 (.I(W2974), .ZN(O11289));
  INVX1 G34053 (.I(W8165), .ZN(W9932));
  INVX1 G34054 (.I(W20725), .ZN(O11291));
  INVX1 G34055 (.I(W2103), .ZN(O11264));
  INVX1 G34056 (.I(W35941), .ZN(O13242));
  INVX1 G34057 (.I(W22554), .ZN(O13261));
  INVX1 G34058 (.I(W8433), .ZN(O13401));
  INVX1 G34059 (.I(W7070), .ZN(W7299));
  INVX1 G34060 (.I(W1595), .ZN(W10084));
  INVX1 G34061 (.I(I1580), .ZN(W7086));
  INVX1 G34062 (.I(I909), .ZN(W7085));
  INVX1 G34063 (.I(W1179), .ZN(W43807));
  INVX1 G34064 (.I(W1211), .ZN(W7102));
  INVX1 G34065 (.I(W8267), .ZN(W40976));
  INVX1 G34066 (.I(W923), .ZN(W43592));
  INVX1 G34067 (.I(W3938), .ZN(W7300));
  INVX1 G34068 (.I(W39220), .ZN(O13424));
  INVX1 G34069 (.I(W13472), .ZN(O13240));
  INVX1 G34070 (.I(W1171), .ZN(W7301));
  INVX1 G34071 (.I(W1968), .ZN(W7304));
  INVX1 G34072 (.I(W9981), .ZN(O13386));
  INVX1 G34073 (.I(W27026), .ZN(W43587));
  INVX1 G34074 (.I(W3423), .ZN(W7107));
  INVX1 G34075 (.I(W2109), .ZN(W7108));
  INVX1 G34076 (.I(W3339), .ZN(O11284));
  INVX1 G34077 (.I(W1821), .ZN(O344));
  INVX1 G34078 (.I(W5666), .ZN(O361));
  INVX1 G34079 (.I(W168), .ZN(W7082));
  INVX1 G34080 (.I(W37541), .ZN(O13190));
  INVX1 G34081 (.I(W527), .ZN(W7373));
  INVX1 G34082 (.I(W39641), .ZN(W41024));
  INVX1 G34083 (.I(W4181), .ZN(W7230));
  INVX1 G34084 (.I(W5431), .ZN(W7170));
  INVX1 G34085 (.I(W2338), .ZN(O11121));
  INVX1 G34086 (.I(I1022), .ZN(O11236));
  INVX1 G34087 (.I(W7065), .ZN(W9985));
  INVX1 G34088 (.I(W2174), .ZN(W9986));
  INVX1 G34089 (.I(I606), .ZN(W10140));
  INVX1 G34090 (.I(W28816), .ZN(O11184));
  INVX1 G34091 (.I(W8134), .ZN(O11312));
  INVX1 G34092 (.I(W12492), .ZN(O11119));
  INVX1 G34093 (.I(W6575), .ZN(O160));
  INVX1 G34094 (.I(W7540), .ZN(W10042));
  INVX1 G34095 (.I(W113), .ZN(O13189));
  INVX1 G34096 (.I(W1537), .ZN(O13188));
  INVX1 G34097 (.I(W3015), .ZN(W40844));
  INVX1 G34098 (.I(W244), .ZN(W7021));
  INVX1 G34099 (.I(W40479), .ZN(O11313));
  INVX1 G34100 (.I(W4036), .ZN(W9991));
  INVX1 G34101 (.I(W1733), .ZN(O13187));
  INVX1 G34102 (.I(W29961), .ZN(O11118));
  INVX1 G34103 (.I(W21553), .ZN(O13338));
  INVX1 G34104 (.I(W40815), .ZN(W40845));
  INVX1 G34105 (.I(I1497), .ZN(O366));
  INVX1 G34106 (.I(W39183), .ZN(O13197));
  INVX1 G34107 (.I(W32046), .ZN(O11182));
  INVX1 G34108 (.I(W37466), .ZN(O11125));
  INVX1 G34109 (.I(W4906), .ZN(W7369));
  INVX1 G34110 (.I(W480), .ZN(W10134));
  INVX1 G34111 (.I(W3472), .ZN(W7233));
  INVX1 G34112 (.I(W1210), .ZN(W9981));
  INVX1 G34113 (.I(W4424), .ZN(W10043));
  INVX1 G34114 (.I(W6042), .ZN(W10136));
  INVX1 G34115 (.I(W1938), .ZN(W41021));
  INVX1 G34116 (.I(W9273), .ZN(O11241));
  INVX1 G34117 (.I(W3793), .ZN(W9889));
  INVX1 G34118 (.I(I1161), .ZN(W10137));
  INVX1 G34119 (.I(I1323), .ZN(W10148));
  INVX1 G34120 (.I(W29550), .ZN(O13196));
  INVX1 G34121 (.I(W4171), .ZN(W10138));
  INVX1 G34122 (.I(W1476), .ZN(W9983));
  INVX1 G34123 (.I(W31395), .ZN(O11238));
  INVX1 G34124 (.I(W2731), .ZN(O13195));
  INVX1 G34125 (.I(W11538), .ZN(O13341));
  INVX1 G34126 (.I(W3703), .ZN(W7371));
  INVX1 G34127 (.I(I84), .ZN(O13193));
  INVX1 G34128 (.I(W3478), .ZN(W43526));
  INVX1 G34129 (.I(W3500), .ZN(W7372));
  INVX1 G34130 (.I(W3631), .ZN(O348));
  INVX1 G34131 (.I(W1735), .ZN(W7384));
  INVX1 G34132 (.I(W710), .ZN(W7378));
  INVX1 G34133 (.I(W7688), .ZN(W10039));
  INVX1 G34134 (.I(I364), .ZN(W10151));
  INVX1 G34135 (.I(W8599), .ZN(O13455));
  INVX1 G34136 (.I(W9351), .ZN(O355));
  INVX1 G34137 (.I(W20485), .ZN(O13182));
  INVX1 G34138 (.I(W1540), .ZN(W7013));
  INVX1 G34139 (.I(I1166), .ZN(O172));
  INVX1 G34140 (.I(W248), .ZN(W7220));
  INVX1 G34141 (.I(W22296), .ZN(O13181));
  INVX1 G34142 (.I(W23066), .ZN(O11318));
  INVX1 G34143 (.I(I380), .ZN(W7383));
  INVX1 G34144 (.I(W3318), .ZN(W7377));
  INVX1 G34145 (.I(W781), .ZN(W9996));
  INVX1 G34146 (.I(W35995), .ZN(O13298));
  INVX1 G34147 (.I(W2322), .ZN(W7011));
  INVX1 G34148 (.I(W13467), .ZN(O11229));
  INVX1 G34149 (.I(W7277), .ZN(W7387));
  INVX1 G34150 (.I(W3575), .ZN(W10152));
  INVX1 G34151 (.I(I656), .ZN(W7388));
  INVX1 G34152 (.I(W10035), .ZN(W10037));
  INVX1 G34153 (.I(W687), .ZN(W7010));
  INVX1 G34154 (.I(W12602), .ZN(O11190));
  INVX1 G34155 (.I(W25047), .ZN(O11191));
  INVX1 G34156 (.I(W8978), .ZN(O350));
  INVX1 G34157 (.I(W514), .ZN(W7015));
  INVX1 G34158 (.I(W984), .ZN(O13448));
  INVX1 G34159 (.I(W17122), .ZN(W43726));
  INVX1 G34160 (.I(I1698), .ZN(W7172));
  INVX1 G34161 (.I(W35946), .ZN(W43518));
  INVX1 G34162 (.I(W38310), .ZN(O11113));
  INVX1 G34163 (.I(W18935), .ZN(W40740));
  INVX1 G34164 (.I(W8294), .ZN(O11112));
  INVX1 G34165 (.I(W17899), .ZN(O13336));
  INVX1 G34166 (.I(W21657), .ZN(O13294));
  INVX1 G34167 (.I(W28433), .ZN(O13451));
  INVX1 G34168 (.I(W6730), .ZN(W10041));
  INVX1 G34169 (.I(I546), .ZN(W7225));
  INVX1 G34170 (.I(W22683), .ZN(O13443));
  INVX1 G34171 (.I(W39709), .ZN(O11187));
  INVX1 G34172 (.I(W10935), .ZN(W43516));
  INVX1 G34173 (.I(W7776), .ZN(W10150));
  INVX1 G34174 (.I(W10330), .ZN(O13186));
  INVX1 G34175 (.I(I614), .ZN(W7173));
  INVX1 G34176 (.I(W14414), .ZN(W41030));
  INVX1 G34177 (.I(W8733), .ZN(W9994));
  INVX1 G34178 (.I(W32340), .ZN(W43722));
  INVX1 G34179 (.I(W836), .ZN(W9995));
  INVX1 G34180 (.I(W3887), .ZN(W9879));
  INVX1 G34181 (.I(W38640), .ZN(O13453));
  INVX1 G34182 (.I(W1427), .ZN(W7044));
  INVX1 G34183 (.I(W5072), .ZN(W7350));
  INVX1 G34184 (.I(W5581), .ZN(W10055));
  INVX1 G34185 (.I(W6007), .ZN(W7151));
  INVX1 G34186 (.I(W20416), .ZN(W40934));
  INVX1 G34187 (.I(W12477), .ZN(W40826));
  INVX1 G34188 (.I(W1840), .ZN(W9903));
  INVX1 G34189 (.I(W21369), .ZN(O11251));
  INVX1 G34190 (.I(W18039), .ZN(O11303));
  INVX1 G34191 (.I(W23637), .ZN(O13208));
  INVX1 G34192 (.I(W1959), .ZN(O13207));
  INVX1 G34193 (.I(W1281), .ZN(W40932));
  INVX1 G34194 (.I(W1518), .ZN(O11250));
  INVX1 G34195 (.I(W4465), .ZN(W7045));
  INVX1 G34196 (.I(W808), .ZN(W7154));
  INVX1 G34197 (.I(W9197), .ZN(W10127));
  INVX1 G34198 (.I(W23344), .ZN(W43742));
  INVX1 G34199 (.I(W5830), .ZN(O11173));
  INVX1 G34200 (.I(W1715), .ZN(W10053));
  INVX1 G34201 (.I(W4473), .ZN(W9900));
  INVX1 G34202 (.I(W10941), .ZN(O11127));
  INVX1 G34203 (.I(W1453), .ZN(O163));
  INVX1 G34204 (.I(W6101), .ZN(W7351));
  INVX1 G34205 (.I(W25421), .ZN(W40759));
  INVX1 G34206 (.I(W9643), .ZN(W9898));
  INVX1 G34207 (.I(W1558), .ZN(W7353));
  INVX1 G34208 (.I(W1383), .ZN(O13280));
  INVX1 G34209 (.I(W6777), .ZN(W7144));
  INVX1 G34210 (.I(W2132), .ZN(W9915));
  INVX1 G34211 (.I(W2504), .ZN(W7145));
  INVX1 G34212 (.I(W22084), .ZN(W40822));
  INVX1 G34213 (.I(W7772), .ZN(W9914));
  INVX1 G34214 (.I(W1896), .ZN(W7338));
  INVX1 G34215 (.I(W4369), .ZN(W7247));
  INVX1 G34216 (.I(W5042), .ZN(W10118));
  INVX1 G34217 (.I(I428), .ZN(W7050));
  INVX1 G34218 (.I(W3897), .ZN(W7048));
  INVX1 G34219 (.I(W955), .ZN(W7148));
  INVX1 G34220 (.I(W3910), .ZN(O364));
  INVX1 G34221 (.I(W40888), .ZN(O13285));
  INVX1 G34222 (.I(W5176), .ZN(W7344));
  INVX1 G34223 (.I(I1803), .ZN(W10126));
  INVX1 G34224 (.I(W981), .ZN(W7245));
  INVX1 G34225 (.I(W23334), .ZN(W43746));
  INVX1 G34226 (.I(W1247), .ZN(W7345));
  INVX1 G34227 (.I(W743), .ZN(W9909));
  INVX1 G34228 (.I(W21778), .ZN(O13282));
  INVX1 G34229 (.I(W6333), .ZN(W7046));
  INVX1 G34230 (.I(I998), .ZN(W9907));
  INVX1 G34231 (.I(W18062), .ZN(W43842));
  INVX1 G34232 (.I(W20594), .ZN(O13210));
  INVX1 G34233 (.I(W5300), .ZN(W9892));
  INVX1 G34234 (.I(W580), .ZN(O11179));
  INVX1 G34235 (.I(W8988), .ZN(W10047));
  INVX1 G34236 (.I(W8385), .ZN(W10046));
  INVX1 G34237 (.I(W32470), .ZN(O13345));
  INVX1 G34238 (.I(W17441), .ZN(O11244));
  INVX1 G34239 (.I(W6087), .ZN(O13437));
  INVX1 G34240 (.I(W4190), .ZN(W10045));
  INVX1 G34241 (.I(W5672), .ZN(O161));
  INVX1 G34242 (.I(I684), .ZN(W7360));
  INVX1 G34243 (.I(W37170), .ZN(O11308));
  INVX1 G34244 (.I(W4668), .ZN(W9894));
  INVX1 G34245 (.I(W5703), .ZN(W7238));
  INVX1 G34246 (.I(W1145), .ZN(W7358));
  INVX1 G34247 (.I(W72), .ZN(W7164));
  INVX1 G34248 (.I(W5814), .ZN(O13439));
  INVX1 G34249 (.I(W39723), .ZN(O13440));
  INVX1 G34250 (.I(W5378), .ZN(W7030));
  INVX1 G34251 (.I(W3435), .ZN(W7237));
  INVX1 G34252 (.I(W695), .ZN(W7367));
  INVX1 G34253 (.I(W4370), .ZN(W7165));
  INVX1 G34254 (.I(W6433), .ZN(O13199));
  INVX1 G34255 (.I(W5798), .ZN(W9978));
  INVX1 G34256 (.I(I1418), .ZN(W7235));
  INVX1 G34257 (.I(I1754), .ZN(W9980));
  INVX1 G34258 (.I(W1335), .ZN(W10050));
  INVX1 G34259 (.I(W6922), .ZN(O13205));
  INVX1 G34260 (.I(W4802), .ZN(O11175));
  INVX1 G34261 (.I(W32656), .ZN(O11248));
  INVX1 G34262 (.I(W6497), .ZN(W7354));
  INVX1 G34263 (.I(W4071), .ZN(W7036));
  INVX1 G34264 (.I(I1060), .ZN(O13432));
  INVX1 G34265 (.I(W3546), .ZN(W7240));
  INVX1 G34266 (.I(W38270), .ZN(O13433));
  INVX1 G34267 (.I(W6771), .ZN(O11247));
  INVX1 G34268 (.I(W1621), .ZN(W7355));
  INVX1 G34269 (.I(W6272), .ZN(W43541));
  INVX1 G34270 (.I(W3695), .ZN(W7159));
  INVX1 G34271 (.I(W25941), .ZN(O11228));
  INVX1 G34272 (.I(W27828), .ZN(O13286));
  INVX1 G34273 (.I(I1727), .ZN(W10049));
  INVX1 G34274 (.I(W11221), .ZN(O11177));
  INVX1 G34275 (.I(W12232), .ZN(O13287));
  INVX1 G34276 (.I(W27072), .ZN(W41015));
  INVX1 G34277 (.I(W4164), .ZN(W7357));
  INVX1 G34278 (.I(W4831), .ZN(W7035));
  INVX1 G34279 (.I(W29751), .ZN(O11246));
  INVX1 G34280 (.I(W9509), .ZN(W10131));
  INVX1 G34281 (.I(W35054), .ZN(O13435));
  INVX1 G34282 (.I(W19757), .ZN(O13346));
  INVX1 G34283 (.I(W12048), .ZN(O12450));
  INVX1 G34284 (.I(W39349), .ZN(O11863));
  INVX1 G34285 (.I(W33387), .ZN(O11860));
  INVX1 G34286 (.I(W26791), .ZN(O12445));
  INVX1 G34287 (.I(W35805), .ZN(O11859));
  INVX1 G34288 (.I(W24934), .ZN(O11858));
  INVX1 G34289 (.I(W16376), .ZN(W41792));
  INVX1 G34290 (.I(W2266), .ZN(W9120));
  INVX1 G34291 (.I(W8925), .ZN(W9122));
  INVX1 G34292 (.I(W40200), .ZN(O11855));
  INVX1 G34293 (.I(W16389), .ZN(W42570));
  INVX1 G34294 (.I(W12715), .ZN(W41788));
  INVX1 G34295 (.I(W8311), .ZN(W8319));
  INVX1 G34296 (.I(W3535), .ZN(W8330));
  INVX1 G34297 (.I(W29557), .ZN(O11854));
  INVX1 G34298 (.I(W886), .ZN(W8317));
  INVX1 G34299 (.I(I246), .ZN(O11853));
  INVX1 G34300 (.I(W5272), .ZN(W8311));
  INVX1 G34301 (.I(W26135), .ZN(O12453));
  INVX1 G34302 (.I(W23215), .ZN(O11852));
  INVX1 G34303 (.I(W3201), .ZN(W41784));
  INVX1 G34304 (.I(W31707), .ZN(O11851));
  INVX1 G34305 (.I(W16430), .ZN(W42580));
  INVX1 G34306 (.I(W20385), .ZN(O11850));
  INVX1 G34307 (.I(W5144), .ZN(W8306));
  INVX1 G34308 (.I(W24590), .ZN(O12458));
  INVX1 G34309 (.I(W8999), .ZN(W9111));
  INVX1 G34310 (.I(I1421), .ZN(W9100));
  INVX1 G34311 (.I(W15282), .ZN(O12429));
  INVX1 G34312 (.I(W27162), .ZN(O12430));
  INVX1 G34313 (.I(W3008), .ZN(W9101));
  INVX1 G34314 (.I(W3244), .ZN(W9102));
  INVX1 G34315 (.I(W690), .ZN(O11871));
  INVX1 G34316 (.I(W2074), .ZN(W9104));
  INVX1 G34317 (.I(W34752), .ZN(O11869));
  INVX1 G34318 (.I(W6393), .ZN(O12431));
  INVX1 G34319 (.I(W36188), .ZN(W41808));
  INVX1 G34320 (.I(W2355), .ZN(W8338));
  INVX1 G34321 (.I(W7920), .ZN(O12433));
  INVX1 G34322 (.I(W8411), .ZN(W9123));
  INVX1 G34323 (.I(W6329), .ZN(O12435));
  INVX1 G34324 (.I(W6473), .ZN(W9113));
  INVX1 G34325 (.I(W2007), .ZN(O265));
  INVX1 G34326 (.I(W15338), .ZN(O12438));
  INVX1 G34327 (.I(W41005), .ZN(O11865));
  INVX1 G34328 (.I(W8717), .ZN(O12439));
  INVX1 G34329 (.I(W7803), .ZN(O11864));
  INVX1 G34330 (.I(W30084), .ZN(O12440));
  INVX1 G34331 (.I(W39304), .ZN(O12441));
  INVX1 G34332 (.I(W27548), .ZN(O12442));
  INVX1 G34333 (.I(W39962), .ZN(O12443));
  INVX1 G34334 (.I(W13492), .ZN(O12485));
  INVX1 G34335 (.I(W20935), .ZN(O12477));
  INVX1 G34336 (.I(W4680), .ZN(W9139));
  INVX1 G34337 (.I(W34166), .ZN(O11841));
  INVX1 G34338 (.I(W20094), .ZN(O11840));
  INVX1 G34339 (.I(W5561), .ZN(W8286));
  INVX1 G34340 (.I(W36448), .ZN(O12479));
  INVX1 G34341 (.I(W6732), .ZN(O11839));
  INVX1 G34342 (.I(W5027), .ZN(W9140));
  INVX1 G34343 (.I(W39671), .ZN(O11837));
  INVX1 G34344 (.I(W6767), .ZN(O221));
  INVX1 G34345 (.I(W40241), .ZN(O12481));
  INVX1 G34346 (.I(W24164), .ZN(O12483));
  INVX1 G34347 (.I(W11484), .ZN(O11844));
  INVX1 G34348 (.I(W252), .ZN(W8278));
  INVX1 G34349 (.I(W23316), .ZN(O12487));
  INVX1 G34350 (.I(W6301), .ZN(W9143));
  INVX1 G34351 (.I(W6855), .ZN(W9144));
  INVX1 G34352 (.I(W39921), .ZN(O12489));
  INVX1 G34353 (.I(W33485), .ZN(O12490));
  INVX1 G34354 (.I(W4650), .ZN(W8276));
  INVX1 G34355 (.I(W39379), .ZN(W42629));
  INVX1 G34356 (.I(W5271), .ZN(W8275));
  INVX1 G34357 (.I(W3009), .ZN(W8271));
  INVX1 G34358 (.I(W3688), .ZN(W8266));
  INVX1 G34359 (.I(W7918), .ZN(W9129));
  INVX1 G34360 (.I(I236), .ZN(W8303));
  INVX1 G34361 (.I(W6467), .ZN(W41780));
  INVX1 G34362 (.I(W29289), .ZN(O12462));
  INVX1 G34363 (.I(W31234), .ZN(O12463));
  INVX1 G34364 (.I(W24642), .ZN(O12465));
  INVX1 G34365 (.I(W32664), .ZN(W42594));
  INVX1 G34366 (.I(W5659), .ZN(W9125));
  INVX1 G34367 (.I(W20431), .ZN(W42595));
  INVX1 G34368 (.I(W10709), .ZN(O12466));
  INVX1 G34369 (.I(I1884), .ZN(W9127));
  INVX1 G34370 (.I(W6222), .ZN(W8299));
  INVX1 G34371 (.I(I431), .ZN(W8298));
  INVX1 G34372 (.I(W37621), .ZN(O12426));
  INVX1 G34373 (.I(W4191), .ZN(W8296));
  INVX1 G34374 (.I(W8957), .ZN(W9131));
  INVX1 G34375 (.I(I1993), .ZN(W9132));
  INVX1 G34376 (.I(W41864), .ZN(W42602));
  INVX1 G34377 (.I(W14040), .ZN(O12471));
  INVX1 G34378 (.I(W5915), .ZN(W9133));
  INVX1 G34379 (.I(W5629), .ZN(W9135));
  INVX1 G34380 (.I(W41869), .ZN(W42606));
  INVX1 G34381 (.I(W23216), .ZN(O12473));
  INVX1 G34382 (.I(W22066), .ZN(O12474));
  INVX1 G34383 (.I(W2076), .ZN(O12475));
  INVX1 G34384 (.I(W8528), .ZN(W9069));
  INVX1 G34385 (.I(W1289), .ZN(W42478));
  INVX1 G34386 (.I(W39572), .ZN(W41855));
  INVX1 G34387 (.I(W2), .ZN(W8411));
  INVX1 G34388 (.I(W7886), .ZN(W9063));
  INVX1 G34389 (.I(W4970), .ZN(O12375));
  INVX1 G34390 (.I(W1882), .ZN(W9066));
  INVX1 G34391 (.I(W34426), .ZN(O12376));
  INVX1 G34392 (.I(W21668), .ZN(O12377));
  INVX1 G34393 (.I(W12850), .ZN(W41851));
  INVX1 G34394 (.I(W6200), .ZN(O12378));
  INVX1 G34395 (.I(W33298), .ZN(O12379));
  INVX1 G34396 (.I(W29284), .ZN(O12381));
  INVX1 G34397 (.I(W20181), .ZN(W41856));
  INVX1 G34398 (.I(W29697), .ZN(O12383));
  INVX1 G34399 (.I(W252), .ZN(O12384));
  INVX1 G34400 (.I(W1907), .ZN(W9070));
  INVX1 G34401 (.I(I128), .ZN(W9071));
  INVX1 G34402 (.I(W1831), .ZN(W8399));
  INVX1 G34403 (.I(W33588), .ZN(O12388));
  INVX1 G34404 (.I(W9841), .ZN(O12389));
  INVX1 G34405 (.I(I1602), .ZN(W8398));
  INVX1 G34406 (.I(W3181), .ZN(W8397));
  INVX1 G34407 (.I(I1950), .ZN(W8394));
  INVX1 G34408 (.I(W36107), .ZN(O12393));
  INVX1 G34409 (.I(W1418), .ZN(W8416));
  INVX1 G34410 (.I(W5623), .ZN(O12358));
  INVX1 G34411 (.I(W7431), .ZN(W9045));
  INVX1 G34412 (.I(W15171), .ZN(O12359));
  INVX1 G34413 (.I(W11211), .ZN(O12360));
  INVX1 G34414 (.I(W5907), .ZN(W8424));
  INVX1 G34415 (.I(W8538), .ZN(W9047));
  INVX1 G34416 (.I(W8964), .ZN(W41866));
  INVX1 G34417 (.I(I535), .ZN(W9048));
  INVX1 G34418 (.I(I1338), .ZN(W9049));
  INVX1 G34419 (.I(W30), .ZN(W8419));
  INVX1 G34420 (.I(W4679), .ZN(W8418));
  INVX1 G34421 (.I(I1103), .ZN(W41861));
  INVX1 G34422 (.I(I1175), .ZN(W8393));
  INVX1 G34423 (.I(I639), .ZN(W9056));
  INVX1 G34424 (.I(W29626), .ZN(W42470));
  INVX1 G34425 (.I(I1005), .ZN(O12368));
  INVX1 G34426 (.I(W5396), .ZN(W9058));
  INVX1 G34427 (.I(W5610), .ZN(W8414));
  INVX1 G34428 (.I(I480), .ZN(O11903));
  INVX1 G34429 (.I(W10230), .ZN(O12371));
  INVX1 G34430 (.I(W8561), .ZN(W9060));
  INVX1 G34431 (.I(W98), .ZN(O12372));
  INVX1 G34432 (.I(W4932), .ZN(O12373));
  INVX1 G34433 (.I(W1776), .ZN(W8413));
  INVX1 G34434 (.I(W122), .ZN(W8361));
  INVX1 G34435 (.I(W34353), .ZN(W42527));
  INVX1 G34436 (.I(W7292), .ZN(W9085));
  INVX1 G34437 (.I(W5775), .ZN(W8367));
  INVX1 G34438 (.I(W33272), .ZN(W42529));
  INVX1 G34439 (.I(I337), .ZN(O12414));
  INVX1 G34440 (.I(W10568), .ZN(W41828));
  INVX1 G34441 (.I(W1013), .ZN(W41827));
  INVX1 G34442 (.I(W10134), .ZN(O11881));
  INVX1 G34443 (.I(W136), .ZN(W9086));
  INVX1 G34444 (.I(W27092), .ZN(O11880));
  INVX1 G34445 (.I(W41565), .ZN(O12417));
  INVX1 G34446 (.I(W12621), .ZN(O12418));
  INVX1 G34447 (.I(W4657), .ZN(W8369));
  INVX1 G34448 (.I(W23052), .ZN(O12419));
  INVX1 G34449 (.I(W4082), .ZN(W9090));
  INVX1 G34450 (.I(W41499), .ZN(O11878));
  INVX1 G34451 (.I(W35762), .ZN(W42540));
  INVX1 G34452 (.I(W7696), .ZN(W9092));
  INVX1 G34453 (.I(I198), .ZN(W8357));
  INVX1 G34454 (.I(W18420), .ZN(W42542));
  INVX1 G34455 (.I(W35036), .ZN(O12422));
  INVX1 G34456 (.I(W6100), .ZN(W8350));
  INVX1 G34457 (.I(W31783), .ZN(O11876));
  INVX1 G34458 (.I(W2922), .ZN(W9097));
  INVX1 G34459 (.I(W6512), .ZN(W8384));
  INVX1 G34460 (.I(W5089), .ZN(W9076));
  INVX1 G34461 (.I(W1934), .ZN(O12395));
  INVX1 G34462 (.I(I1394), .ZN(O12397));
  INVX1 G34463 (.I(W38259), .ZN(O12398));
  INVX1 G34464 (.I(I1991), .ZN(W9078));
  INVX1 G34465 (.I(W22349), .ZN(O12400));
  INVX1 G34466 (.I(W31929), .ZN(O11889));
  INVX1 G34467 (.I(W39313), .ZN(W42508));
  INVX1 G34468 (.I(W34267), .ZN(O12401));
  INVX1 G34469 (.I(W5209), .ZN(W8390));
  INVX1 G34470 (.I(W5479), .ZN(W8388));
  INVX1 G34471 (.I(W1286), .ZN(W8387));
  INVX1 G34472 (.I(W923), .ZN(W8265));
  INVX1 G34473 (.I(W6074), .ZN(W8383));
  INVX1 G34474 (.I(W37976), .ZN(O12407));
  INVX1 G34475 (.I(W3170), .ZN(W41839));
  INVX1 G34476 (.I(W22859), .ZN(W42518));
  INVX1 G34477 (.I(W13536), .ZN(O11888));
  INVX1 G34478 (.I(W15195), .ZN(O11887));
  INVX1 G34479 (.I(W9707), .ZN(O11886));
  INVX1 G34480 (.I(W41276), .ZN(W42521));
  INVX1 G34481 (.I(I1421), .ZN(W9079));
  INVX1 G34482 (.I(W26155), .ZN(O11885));
  INVX1 G34483 (.I(W36165), .ZN(W41833));
  INVX1 G34484 (.I(W9193), .ZN(W9274));
  INVX1 G34485 (.I(I909), .ZN(W8135));
  INVX1 G34486 (.I(W981), .ZN(W8134));
  INVX1 G34487 (.I(W8261), .ZN(O11770));
  INVX1 G34488 (.I(W6686), .ZN(W9265));
  INVX1 G34489 (.I(W6657), .ZN(W9266));
  INVX1 G34490 (.I(W21574), .ZN(O12590));
  INVX1 G34491 (.I(W6892), .ZN(W8131));
  INVX1 G34492 (.I(W4589), .ZN(O12592));
  INVX1 G34493 (.I(W9237), .ZN(W9269));
  INVX1 G34494 (.I(W8792), .ZN(O12593));
  INVX1 G34495 (.I(W1282), .ZN(W9273));
  INVX1 G34496 (.I(W21645), .ZN(O12594));
  INVX1 G34497 (.I(I1452), .ZN(W9263));
  INVX1 G34498 (.I(I919), .ZN(W8130));
  INVX1 G34499 (.I(W22811), .ZN(O11763));
  INVX1 G34500 (.I(W1137), .ZN(W9275));
  INVX1 G34501 (.I(W28461), .ZN(O12597));
  INVX1 G34502 (.I(W17207), .ZN(O12598));
  INVX1 G34503 (.I(W41160), .ZN(O12599));
  INVX1 G34504 (.I(W1152), .ZN(W9276));
  INVX1 G34505 (.I(W7652), .ZN(W8125));
  INVX1 G34506 (.I(W8103), .ZN(W8123));
  INVX1 G34507 (.I(W5331), .ZN(W8122));
  INVX1 G34508 (.I(W17856), .ZN(O11761));
  INVX1 G34509 (.I(I1146), .ZN(W9253));
  INVX1 G34510 (.I(W889), .ZN(W8169));
  INVX1 G34511 (.I(W8928), .ZN(W9243));
  INVX1 G34512 (.I(I1596), .ZN(W8166));
  INVX1 G34513 (.I(I1461), .ZN(W8165));
  INVX1 G34514 (.I(W5360), .ZN(W8163));
  INVX1 G34515 (.I(W5827), .ZN(W9245));
  INVX1 G34516 (.I(W1188), .ZN(W9246));
  INVX1 G34517 (.I(W19724), .ZN(O12574));
  INVX1 G34518 (.I(W6677), .ZN(W8157));
  INVX1 G34519 (.I(W3818), .ZN(W9251));
  INVX1 G34520 (.I(W84), .ZN(W9252));
  INVX1 G34521 (.I(I112), .ZN(W8154));
  INVX1 G34522 (.I(W2682), .ZN(O278));
  INVX1 G34523 (.I(I913), .ZN(W8151));
  INVX1 G34524 (.I(W1821), .ZN(W9258));
  INVX1 G34525 (.I(W36355), .ZN(O11772));
  INVX1 G34526 (.I(W27878), .ZN(O11771));
  INVX1 G34527 (.I(W1148), .ZN(W8147));
  INVX1 G34528 (.I(W17152), .ZN(O12582));
  INVX1 G34529 (.I(W14991), .ZN(W42745));
  INVX1 G34530 (.I(W8223), .ZN(W9260));
  INVX1 G34531 (.I(I113), .ZN(W8142));
  INVX1 G34532 (.I(W18948), .ZN(O12584));
  INVX1 G34533 (.I(W12146), .ZN(O12588));
  INVX1 G34534 (.I(W306), .ZN(W9321));
  INVX1 G34535 (.I(W7284), .ZN(W8098));
  INVX1 G34536 (.I(W6051), .ZN(W8096));
  INVX1 G34537 (.I(W6522), .ZN(W9309));
  INVX1 G34538 (.I(I989), .ZN(W9311));
  INVX1 G34539 (.I(W2548), .ZN(W9317));
  INVX1 G34540 (.I(W7518), .ZN(W8091));
  INVX1 G34541 (.I(W14581), .ZN(O12616));
  INVX1 G34542 (.I(W6263), .ZN(W41620));
  INVX1 G34543 (.I(W11664), .ZN(O11736));
  INVX1 G34544 (.I(W42510), .ZN(O12618));
  INVX1 G34545 (.I(W7740), .ZN(O211));
  INVX1 G34546 (.I(W2245), .ZN(W8084));
  INVX1 G34547 (.I(W14923), .ZN(W42788));
  INVX1 G34548 (.I(W29627), .ZN(W41616));
  INVX1 G34549 (.I(W26659), .ZN(O11733));
  INVX1 G34550 (.I(I488), .ZN(W8081));
  INVX1 G34551 (.I(W3906), .ZN(O11732));
  INVX1 G34552 (.I(W35281), .ZN(O12621));
  INVX1 G34553 (.I(I227), .ZN(W9323));
  INVX1 G34554 (.I(W30670), .ZN(O12623));
  INVX1 G34555 (.I(W6503), .ZN(W8075));
  INVX1 G34556 (.I(W21214), .ZN(O11729));
  INVX1 G34557 (.I(W5637), .ZN(W9329));
  INVX1 G34558 (.I(W7022), .ZN(W8072));
  INVX1 G34559 (.I(W2117), .ZN(W9295));
  INVX1 G34560 (.I(W3183), .ZN(W9280));
  INVX1 G34561 (.I(W7266), .ZN(W9281));
  INVX1 G34562 (.I(W29322), .ZN(W42771));
  INVX1 G34563 (.I(W13062), .ZN(W41647));
  INVX1 G34564 (.I(W3913), .ZN(W9283));
  INVX1 G34565 (.I(W9030), .ZN(W9285));
  INVX1 G34566 (.I(W28096), .ZN(W42772));
  INVX1 G34567 (.I(W31504), .ZN(W41643));
  INVX1 G34568 (.I(W5568), .ZN(W9290));
  INVX1 G34569 (.I(W25032), .ZN(O11754));
  INVX1 G34570 (.I(W4110), .ZN(W8114));
  INVX1 G34571 (.I(W13141), .ZN(O12607));
  INVX1 G34572 (.I(W7867), .ZN(W9242));
  INVX1 G34573 (.I(W2805), .ZN(W9297));
  INVX1 G34574 (.I(W39895), .ZN(O11750));
  INVX1 G34575 (.I(W15278), .ZN(O12609));
  INVX1 G34576 (.I(W2029), .ZN(W9300));
  INVX1 G34577 (.I(W3695), .ZN(W8108));
  INVX1 G34578 (.I(W7762), .ZN(W9301));
  INVX1 G34579 (.I(W39791), .ZN(O11747));
  INVX1 G34580 (.I(W19955), .ZN(W42783));
  INVX1 G34581 (.I(W27848), .ZN(O12611));
  INVX1 G34582 (.I(I1841), .ZN(O11746));
  INVX1 G34583 (.I(W1671), .ZN(W9302));
  INVX1 G34584 (.I(I1554), .ZN(W8224));
  INVX1 G34585 (.I(I1172), .ZN(W8241));
  INVX1 G34586 (.I(W1784), .ZN(W8239));
  INVX1 G34587 (.I(W6282), .ZN(W9187));
  INVX1 G34588 (.I(W3763), .ZN(W42658));
  INVX1 G34589 (.I(W17452), .ZN(O12513));
  INVX1 G34590 (.I(W14083), .ZN(O12514));
  INVX1 G34591 (.I(W6377), .ZN(O12515));
  INVX1 G34592 (.I(W7325), .ZN(W8235));
  INVX1 G34593 (.I(W2584), .ZN(W8234));
  INVX1 G34594 (.I(W35252), .ZN(O12518));
  INVX1 G34595 (.I(W5724), .ZN(O12520));
  INVX1 G34596 (.I(W5289), .ZN(O11814));
  INVX1 G34597 (.I(I990), .ZN(W9184));
  INVX1 G34598 (.I(W31534), .ZN(O12524));
  INVX1 G34599 (.I(W5097), .ZN(W9192));
  INVX1 G34600 (.I(W27608), .ZN(O11812));
  INVX1 G34601 (.I(W3104), .ZN(W8220));
  INVX1 G34602 (.I(W18537), .ZN(O11810));
  INVX1 G34603 (.I(W37198), .ZN(O11808));
  INVX1 G34604 (.I(W24594), .ZN(O12527));
  INVX1 G34605 (.I(W1137), .ZN(O11807));
  INVX1 G34606 (.I(W27083), .ZN(O12528));
  INVX1 G34607 (.I(W1219), .ZN(O11806));
  INVX1 G34608 (.I(W6639), .ZN(W9197));
  INVX1 G34609 (.I(W7036), .ZN(W9165));
  INVX1 G34610 (.I(W6355), .ZN(O269));
  INVX1 G34611 (.I(W22164), .ZN(O12497));
  INVX1 G34612 (.I(W22368), .ZN(O11832));
  INVX1 G34613 (.I(W8628), .ZN(O11831));
  INVX1 G34614 (.I(W250), .ZN(W8256));
  INVX1 G34615 (.I(W17825), .ZN(O11830));
  INVX1 G34616 (.I(W3836), .ZN(W8255));
  INVX1 G34617 (.I(W1828), .ZN(W9152));
  INVX1 G34618 (.I(W5075), .ZN(W9153));
  INVX1 G34619 (.I(I905), .ZN(W8254));
  INVX1 G34620 (.I(W5050), .ZN(W9157));
  INVX1 G34621 (.I(W5943), .ZN(W9159));
  INVX1 G34622 (.I(W5027), .ZN(W42681));
  INVX1 G34623 (.I(W2978), .ZN(W8248));
  INVX1 G34624 (.I(W27867), .ZN(W42648));
  INVX1 G34625 (.I(W8103), .ZN(W9171));
  INVX1 G34626 (.I(W1395), .ZN(W8246));
  INVX1 G34627 (.I(W12677), .ZN(O12507));
  INVX1 G34628 (.I(W3339), .ZN(W9176));
  INVX1 G34629 (.I(W8290), .ZN(W9179));
  INVX1 G34630 (.I(W35460), .ZN(O12509));
  INVX1 G34631 (.I(W6164), .ZN(W9182));
  INVX1 G34632 (.I(W3650), .ZN(W9183));
  INVX1 G34633 (.I(W15180), .ZN(O11818));
  INVX1 G34634 (.I(W31650), .ZN(O12559));
  INVX1 G34635 (.I(W1535), .ZN(W9225));
  INVX1 G34636 (.I(W932), .ZN(O11787));
  INVX1 G34637 (.I(W15347), .ZN(O12553));
  INVX1 G34638 (.I(I900), .ZN(W8186));
  INVX1 G34639 (.I(W32429), .ZN(O11786));
  INVX1 G34640 (.I(W1598), .ZN(W9229));
  INVX1 G34641 (.I(W20513), .ZN(O12555));
  INVX1 G34642 (.I(W8308), .ZN(W9231));
  INVX1 G34643 (.I(W5920), .ZN(W8181));
  INVX1 G34644 (.I(W15735), .ZN(O11784));
  INVX1 G34645 (.I(W15269), .ZN(O12558));
  INVX1 G34646 (.I(W9166), .ZN(W9233));
  INVX1 G34647 (.I(W5142), .ZN(W9222));
  INVX1 G34648 (.I(W37939), .ZN(O12560));
  INVX1 G34649 (.I(W27732), .ZN(O11782));
  INVX1 G34650 (.I(W5852), .ZN(W9234));
  INVX1 G34651 (.I(W22753), .ZN(O11781));
  INVX1 G34652 (.I(W2625), .ZN(W8178));
  INVX1 G34653 (.I(W24920), .ZN(W42719));
  INVX1 G34654 (.I(W25179), .ZN(O12563));
  INVX1 G34655 (.I(W6311), .ZN(W8177));
  INVX1 G34656 (.I(W32230), .ZN(O12565));
  INVX1 G34657 (.I(W2664), .ZN(O12566));
  INVX1 G34658 (.I(W7885), .ZN(W9241));
  INVX1 G34659 (.I(W2961), .ZN(W9207));
  INVX1 G34660 (.I(W2560), .ZN(O215));
  INVX1 G34661 (.I(W16907), .ZN(O11805));
  INVX1 G34662 (.I(W5620), .ZN(W9200));
  INVX1 G34663 (.I(W23168), .ZN(O12535));
  INVX1 G34664 (.I(W13640), .ZN(O12536));
  INVX1 G34665 (.I(W15361), .ZN(O12537));
  INVX1 G34666 (.I(W5585), .ZN(W9202));
  INVX1 G34667 (.I(W2654), .ZN(W8202));
  INVX1 G34668 (.I(W6920), .ZN(W9204));
  INVX1 G34669 (.I(I1734), .ZN(W8201));
  INVX1 G34670 (.I(W38831), .ZN(O11800));
  INVX1 G34671 (.I(W4921), .ZN(W42693));
  INVX1 G34672 (.I(W10945), .ZN(O12357));
  INVX1 G34673 (.I(W5499), .ZN(W8198));
  INVX1 G34674 (.I(W1536), .ZN(W9211));
  INVX1 G34675 (.I(I1913), .ZN(O11794));
  INVX1 G34676 (.I(W6262), .ZN(W9217));
  INVX1 G34677 (.I(I983), .ZN(W9218));
  INVX1 G34678 (.I(W7405), .ZN(O275));
  INVX1 G34679 (.I(W20613), .ZN(W41698));
  INVX1 G34680 (.I(W8914), .ZN(O11790));
  INVX1 G34681 (.I(W6048), .ZN(W8190));
  INVX1 G34682 (.I(W24597), .ZN(O12548));
  INVX1 G34683 (.I(W6322), .ZN(O12549));
  INVX1 G34684 (.I(W37073), .ZN(O12052));
  INVX1 G34685 (.I(W5440), .ZN(W8660));
  INVX1 G34686 (.I(W22564), .ZN(O12059));
  INVX1 G34687 (.I(I1034), .ZN(W8853));
  INVX1 G34688 (.I(W33884), .ZN(O12198));
  INVX1 G34689 (.I(W34419), .ZN(O12057));
  INVX1 G34690 (.I(W29850), .ZN(W42245));
  INVX1 G34691 (.I(I483), .ZN(W8855));
  INVX1 G34692 (.I(W19910), .ZN(O12055));
  INVX1 G34693 (.I(W7454), .ZN(W8651));
  INVX1 G34694 (.I(W5320), .ZN(O12054));
  INVX1 G34695 (.I(W9788), .ZN(W42251));
  INVX1 G34696 (.I(I1421), .ZN(W8860));
  INVX1 G34697 (.I(W6853), .ZN(W8661));
  INVX1 G34698 (.I(W3364), .ZN(W8644));
  INVX1 G34699 (.I(W2519), .ZN(W8642));
  INVX1 G34700 (.I(W3802), .ZN(W8862));
  INVX1 G34701 (.I(W8656), .ZN(O12209));
  INVX1 G34702 (.I(W3389), .ZN(W8863));
  INVX1 G34703 (.I(I1462), .ZN(W8638));
  INVX1 G34704 (.I(I815), .ZN(W8634));
  INVX1 G34705 (.I(W13385), .ZN(O12213));
  INVX1 G34706 (.I(I396), .ZN(W8865));
  INVX1 G34707 (.I(W6773), .ZN(W8866));
  INVX1 G34708 (.I(W26655), .ZN(O12214));
  INVX1 G34709 (.I(W7875), .ZN(W8867));
  INVX1 G34710 (.I(W2525), .ZN(W8668));
  INVX1 G34711 (.I(W1151), .ZN(O249));
  INVX1 G34712 (.I(W4413), .ZN(W8682));
  INVX1 G34713 (.I(W823), .ZN(W8835));
  INVX1 G34714 (.I(W3882), .ZN(O12070));
  INVX1 G34715 (.I(I1390), .ZN(W8840));
  INVX1 G34716 (.I(W17711), .ZN(O12184));
  INVX1 G34717 (.I(W2581), .ZN(W8843));
  INVX1 G34718 (.I(W10704), .ZN(O12186));
  INVX1 G34719 (.I(W1151), .ZN(W8676));
  INVX1 G34720 (.I(W5857), .ZN(W8675));
  INVX1 G34721 (.I(W4364), .ZN(W8674));
  INVX1 G34722 (.I(W6263), .ZN(W8672));
  INVX1 G34723 (.I(W32086), .ZN(W42044));
  INVX1 G34724 (.I(W12791), .ZN(O12193));
  INVX1 G34725 (.I(I888), .ZN(W8847));
  INVX1 G34726 (.I(I195), .ZN(W8848));
  INVX1 G34727 (.I(W34859), .ZN(O12062));
  INVX1 G34728 (.I(W18930), .ZN(W42237));
  INVX1 G34729 (.I(W22468), .ZN(W42065));
  INVX1 G34730 (.I(W3837), .ZN(W8852));
  INVX1 G34731 (.I(W9140), .ZN(W42063));
  INVX1 G34732 (.I(I1663), .ZN(W8664));
  INVX1 G34733 (.I(W37354), .ZN(O12061));
  INVX1 G34734 (.I(W35222), .ZN(O12060));
  INVX1 G34735 (.I(W8276), .ZN(W8889));
  INVX1 G34736 (.I(W2498), .ZN(O237));
  INVX1 G34737 (.I(W27824), .ZN(O12035));
  INVX1 G34738 (.I(I1392), .ZN(W8604));
  INVX1 G34739 (.I(W30437), .ZN(O12034));
  INVX1 G34740 (.I(W30319), .ZN(O12235));
  INVX1 G34741 (.I(W16171), .ZN(O12033));
  INVX1 G34742 (.I(W4153), .ZN(W8600));
  INVX1 G34743 (.I(W11538), .ZN(O12032));
  INVX1 G34744 (.I(W7766), .ZN(W8882));
  INVX1 G34745 (.I(W23048), .ZN(O12030));
  INVX1 G34746 (.I(W4954), .ZN(W8883));
  INVX1 G34747 (.I(W3433), .ZN(W8886));
  INVX1 G34748 (.I(W1387), .ZN(O12232));
  INVX1 G34749 (.I(W34449), .ZN(O12237));
  INVX1 G34750 (.I(W38362), .ZN(O12238));
  INVX1 G34751 (.I(W24122), .ZN(O12239));
  INVX1 G34752 (.I(W32997), .ZN(O12026));
  INVX1 G34753 (.I(W133), .ZN(W8893));
  INVX1 G34754 (.I(W4898), .ZN(O12024));
  INVX1 G34755 (.I(W30932), .ZN(O12023));
  INVX1 G34756 (.I(I576), .ZN(W8894));
  INVX1 G34757 (.I(W37226), .ZN(O12021));
  INVX1 G34758 (.I(W22805), .ZN(O12242));
  INVX1 G34759 (.I(W436), .ZN(W8897));
  INVX1 G34760 (.I(W6681), .ZN(O12043));
  INVX1 G34761 (.I(W4791), .ZN(W8868));
  INVX1 G34762 (.I(W32844), .ZN(W42042));
  INVX1 G34763 (.I(W22045), .ZN(O12217));
  INVX1 G34764 (.I(I1337), .ZN(W8624));
  INVX1 G34765 (.I(W361), .ZN(W8623));
  INVX1 G34766 (.I(W3755), .ZN(O12220));
  INVX1 G34767 (.I(W35443), .ZN(W42273));
  INVX1 G34768 (.I(W1564), .ZN(W8620));
  INVX1 G34769 (.I(W10869), .ZN(O12045));
  INVX1 G34770 (.I(I1490), .ZN(W8869));
  INVX1 G34771 (.I(W23819), .ZN(W42276));
  INVX1 G34772 (.I(W42242), .ZN(O12223));
  INVX1 G34773 (.I(W911), .ZN(O240));
  INVX1 G34774 (.I(W5295), .ZN(W8872));
  INVX1 G34775 (.I(W18185), .ZN(O12040));
  INVX1 G34776 (.I(I1769), .ZN(O238));
  INVX1 G34777 (.I(W5424), .ZN(O12039));
  INVX1 G34778 (.I(W6949), .ZN(W8873));
  INVX1 G34779 (.I(W5976), .ZN(W8875));
  INVX1 G34780 (.I(W20984), .ZN(O12037));
  INVX1 G34781 (.I(W8679), .ZN(W8876));
  INVX1 G34782 (.I(W3535), .ZN(W8879));
  INVX1 G34783 (.I(W308), .ZN(W8881));
  INVX1 G34784 (.I(W6584), .ZN(W8607));
  INVX1 G34785 (.I(I618), .ZN(W8744));
  INVX1 G34786 (.I(W8158), .ZN(O12097));
  INVX1 G34787 (.I(W1179), .ZN(W8753));
  INVX1 G34788 (.I(W7034), .ZN(W8751));
  INVX1 G34789 (.I(W4219), .ZN(W8750));
  INVX1 G34790 (.I(I698), .ZN(W8799));
  INVX1 G34791 (.I(W22726), .ZN(W42156));
  INVX1 G34792 (.I(W734), .ZN(W42111));
  INVX1 G34793 (.I(W15902), .ZN(O12095));
  INVX1 G34794 (.I(W8384), .ZN(W8800));
  INVX1 G34795 (.I(W7143), .ZN(W8745));
  INVX1 G34796 (.I(W6563), .ZN(O12136));
  INVX1 G34797 (.I(W32109), .ZN(W42106));
  INVX1 G34798 (.I(W20082), .ZN(O12128));
  INVX1 G34799 (.I(W18932), .ZN(O12138));
  INVX1 G34800 (.I(I1709), .ZN(W8742));
  INVX1 G34801 (.I(W2245), .ZN(W8741));
  INVX1 G34802 (.I(W7768), .ZN(W8740));
  INVX1 G34803 (.I(W31449), .ZN(O12142));
  INVX1 G34804 (.I(W2184), .ZN(O12143));
  INVX1 G34805 (.I(W40176), .ZN(O12144));
  INVX1 G34806 (.I(W8608), .ZN(W8806));
  INVX1 G34807 (.I(I1281), .ZN(W8807));
  INVX1 G34808 (.I(W7226), .ZN(W8734));
  INVX1 G34809 (.I(I966), .ZN(W8733));
  INVX1 G34810 (.I(W3906), .ZN(W8770));
  INVX1 G34811 (.I(W696), .ZN(W8785));
  INVX1 G34812 (.I(W5933), .ZN(W8786));
  INVX1 G34813 (.I(W1604), .ZN(W8779));
  INVX1 G34814 (.I(W38912), .ZN(O12106));
  INVX1 G34815 (.I(W7209), .ZN(O246));
  INVX1 G34816 (.I(W36021), .ZN(O12114));
  INVX1 G34817 (.I(W4752), .ZN(W8777));
  INVX1 G34818 (.I(W1022), .ZN(W8775));
  INVX1 G34819 (.I(W23088), .ZN(O12118));
  INVX1 G34820 (.I(I907), .ZN(W8773));
  INVX1 G34821 (.I(W4881), .ZN(W8789));
  INVX1 G34822 (.I(W7515), .ZN(O12120));
  INVX1 G34823 (.I(W7893), .ZN(O12147));
  INVX1 G34824 (.I(W8237), .ZN(W8769));
  INVX1 G34825 (.I(W2936), .ZN(W8791));
  INVX1 G34826 (.I(W376), .ZN(W8792));
  INVX1 G34827 (.I(W4544), .ZN(W8762));
  INVX1 G34828 (.I(W3605), .ZN(W8759));
  INVX1 G34829 (.I(W8191), .ZN(W8756));
  INVX1 G34830 (.I(W16977), .ZN(W42147));
  INVX1 G34831 (.I(W7442), .ZN(O12126));
  INVX1 G34832 (.I(W24477), .ZN(O12127));
  INVX1 G34833 (.I(W28760), .ZN(W42150));
  INVX1 G34834 (.I(W37253), .ZN(O12098));
  INVX1 G34835 (.I(W877), .ZN(W8697));
  INVX1 G34836 (.I(W33788), .ZN(W42089));
  INVX1 G34837 (.I(W1566), .ZN(O242));
  INVX1 G34838 (.I(W36595), .ZN(W42198));
  INVX1 G34839 (.I(I470), .ZN(W42199));
  INVX1 G34840 (.I(W4823), .ZN(W8708));
  INVX1 G34841 (.I(W41609), .ZN(O12167));
  INVX1 G34842 (.I(W7097), .ZN(W8707));
  INVX1 G34843 (.I(W542), .ZN(O12082));
  INVX1 G34844 (.I(W18085), .ZN(O12081));
  INVX1 G34845 (.I(W36733), .ZN(O12170));
  INVX1 G34846 (.I(W26289), .ZN(W42206));
  INVX1 G34847 (.I(W25413), .ZN(O12172));
  INVX1 G34848 (.I(W754), .ZN(W8710));
  INVX1 G34849 (.I(W4343), .ZN(W8696));
  INVX1 G34850 (.I(W2041), .ZN(O12175));
  INVX1 G34851 (.I(I1507), .ZN(W8830));
  INVX1 G34852 (.I(W42094), .ZN(O12176));
  INVX1 G34853 (.I(W13580), .ZN(O12076));
  INVX1 G34854 (.I(W5271), .ZN(W8832));
  INVX1 G34855 (.I(W19886), .ZN(W42080));
  INVX1 G34856 (.I(W710), .ZN(W8685));
  INVX1 G34857 (.I(W7980), .ZN(O12180));
  INVX1 G34858 (.I(W27077), .ZN(O12181));
  INVX1 G34859 (.I(W33186), .ZN(O12182));
  INVX1 G34860 (.I(W4906), .ZN(W8723));
  INVX1 G34861 (.I(W4909), .ZN(W8730));
  INVX1 G34862 (.I(W6834), .ZN(W42177));
  INVX1 G34863 (.I(W14199), .ZN(O12149));
  INVX1 G34864 (.I(W39618), .ZN(O12150));
  INVX1 G34865 (.I(W4004), .ZN(W42180));
  INVX1 G34866 (.I(W34370), .ZN(O12153));
  INVX1 G34867 (.I(W19286), .ZN(O12091));
  INVX1 G34868 (.I(W2222), .ZN(W8725));
  INVX1 G34869 (.I(I969), .ZN(O12155));
  INVX1 G34870 (.I(W6457), .ZN(O12156));
  INVX1 G34871 (.I(W4915), .ZN(W8813));
  INVX1 G34872 (.I(W3844), .ZN(W8724));
  INVX1 G34873 (.I(W1439), .ZN(W8593));
  INVX1 G34874 (.I(W3539), .ZN(W8814));
  INVX1 G34875 (.I(W7904), .ZN(O12158));
  INVX1 G34876 (.I(W6850), .ZN(W8722));
  INVX1 G34877 (.I(W246), .ZN(W8815));
  INVX1 G34878 (.I(W6727), .ZN(O12086));
  INVX1 G34879 (.I(W31118), .ZN(W42094));
  INVX1 G34880 (.I(W23206), .ZN(O12161));
  INVX1 G34881 (.I(W8146), .ZN(W8719));
  INVX1 G34882 (.I(I1599), .ZN(W8816));
  INVX1 G34883 (.I(W2726), .ZN(W8716));
  INVX1 G34884 (.I(I646), .ZN(W8820));
  INVX1 G34885 (.I(W7854), .ZN(O11945));
  INVX1 G34886 (.I(W4458), .ZN(O12311));
  INVX1 G34887 (.I(W1053), .ZN(W8481));
  INVX1 G34888 (.I(I115), .ZN(W8994));
  INVX1 G34889 (.I(I1003), .ZN(W8478));
  INVX1 G34890 (.I(W11901), .ZN(W42404));
  INVX1 G34891 (.I(I1010), .ZN(W8476));
  INVX1 G34892 (.I(W8723), .ZN(W8995));
  INVX1 G34893 (.I(W15185), .ZN(O12316));
  INVX1 G34894 (.I(W20285), .ZN(O12317));
  INVX1 G34895 (.I(W5483), .ZN(W8997));
  INVX1 G34896 (.I(W7757), .ZN(O12318));
  INVX1 G34897 (.I(W811), .ZN(W8998));
  INVX1 G34898 (.I(W15316), .ZN(O11951));
  INVX1 G34899 (.I(W670), .ZN(W8475));
  INVX1 G34900 (.I(W2635), .ZN(W8474));
  INVX1 G34901 (.I(W17322), .ZN(O11944));
  INVX1 G34902 (.I(W2924), .ZN(W8472));
  INVX1 G34903 (.I(W21511), .ZN(O12322));
  INVX1 G34904 (.I(W5025), .ZN(W8471));
  INVX1 G34905 (.I(W25096), .ZN(O11942));
  INVX1 G34906 (.I(W32359), .ZN(O11941));
  INVX1 G34907 (.I(W8682), .ZN(W9003));
  INVX1 G34908 (.I(W4419), .ZN(O232));
  INVX1 G34909 (.I(W38162), .ZN(O12326));
  INVX1 G34910 (.I(W7015), .ZN(O12302));
  INVX1 G34911 (.I(W1847), .ZN(W8979));
  INVX1 G34912 (.I(W5284), .ZN(W8500));
  INVX1 G34913 (.I(W4460), .ZN(O12295));
  INVX1 G34914 (.I(W39955), .ZN(O12296));
  INVX1 G34915 (.I(W8238), .ZN(W8980));
  INVX1 G34916 (.I(W2240), .ZN(W8982));
  INVX1 G34917 (.I(I598), .ZN(W8499));
  INVX1 G34918 (.I(W19141), .ZN(O12297));
  INVX1 G34919 (.I(W5321), .ZN(O11960));
  INVX1 G34920 (.I(W2056), .ZN(W8496));
  INVX1 G34921 (.I(W928), .ZN(W8984));
  INVX1 G34922 (.I(W7967), .ZN(W8494));
  INVX1 G34923 (.I(W31180), .ZN(W42419));
  INVX1 G34924 (.I(W479), .ZN(W8492));
  INVX1 G34925 (.I(W6926), .ZN(W8489));
  INVX1 G34926 (.I(W3295), .ZN(W8986));
  INVX1 G34927 (.I(W9395), .ZN(O12306));
  INVX1 G34928 (.I(W2066), .ZN(W8988));
  INVX1 G34929 (.I(W39556), .ZN(O12307));
  INVX1 G34930 (.I(I29), .ZN(O260));
  INVX1 G34931 (.I(I1086), .ZN(W8991));
  INVX1 G34932 (.I(W6615), .ZN(O11953));
  INVX1 G34933 (.I(W13478), .ZN(O12308));
  INVX1 G34934 (.I(W40307), .ZN(O12309));
  INVX1 G34935 (.I(W6836), .ZN(O227));
  INVX1 G34936 (.I(W3886), .ZN(O229));
  INVX1 G34937 (.I(W383), .ZN(W8443));
  INVX1 G34938 (.I(W38508), .ZN(O11923));
  INVX1 G34939 (.I(W33022), .ZN(O12344));
  INVX1 G34940 (.I(W41664), .ZN(O11920));
  INVX1 G34941 (.I(W5525), .ZN(O12347));
  INVX1 G34942 (.I(W5720), .ZN(O12349));
  INVX1 G34943 (.I(W6601), .ZN(W8436));
  INVX1 G34944 (.I(I1211), .ZN(W9030));
  INVX1 G34945 (.I(W7530), .ZN(W9031));
  INVX1 G34946 (.I(W2881), .ZN(W9033));
  INVX1 G34947 (.I(W5068), .ZN(W9035));
  INVX1 G34948 (.I(W2531), .ZN(W8445));
  INVX1 G34949 (.I(I578), .ZN(W8431));
  INVX1 G34950 (.I(W10912), .ZN(W42452));
  INVX1 G34951 (.I(W1423), .ZN(W9036));
  INVX1 G34952 (.I(W1684), .ZN(W9041));
  INVX1 G34953 (.I(W18376), .ZN(W42453));
  INVX1 G34954 (.I(W7265), .ZN(W42454));
  INVX1 G34955 (.I(W2012), .ZN(W9043));
  INVX1 G34956 (.I(W1370), .ZN(O11911));
  INVX1 G34957 (.I(W349), .ZN(W8429));
  INVX1 G34958 (.I(W32789), .ZN(W41870));
  INVX1 G34959 (.I(W20790), .ZN(O12356));
  INVX1 G34960 (.I(W3610), .ZN(O11931));
  INVX1 G34961 (.I(W11638), .ZN(O12328));
  INVX1 G34962 (.I(I638), .ZN(W9006));
  INVX1 G34963 (.I(I1467), .ZN(W8461));
  INVX1 G34964 (.I(W6638), .ZN(W9008));
  INVX1 G34965 (.I(W41316), .ZN(O11936));
  INVX1 G34966 (.I(W2235), .ZN(W9009));
  INVX1 G34967 (.I(W7284), .ZN(W9010));
  INVX1 G34968 (.I(W10093), .ZN(O12331));
  INVX1 G34969 (.I(W7768), .ZN(W8454));
  INVX1 G34970 (.I(W4382), .ZN(O11933));
  INVX1 G34971 (.I(W2508), .ZN(O261));
  INVX1 G34972 (.I(W36063), .ZN(O12333));
  INVX1 G34973 (.I(W5833), .ZN(W8976));
  INVX1 G34974 (.I(I1838), .ZN(W9016));
  INVX1 G34975 (.I(W38519), .ZN(W41894));
  INVX1 G34976 (.I(W6921), .ZN(W9017));
  INVX1 G34977 (.I(W6201), .ZN(O11928));
  INVX1 G34978 (.I(W5336), .ZN(O11927));
  INVX1 G34979 (.I(W908), .ZN(W9018));
  INVX1 G34980 (.I(W32087), .ZN(W42431));
  INVX1 G34981 (.I(W1830), .ZN(W8448));
  INVX1 G34982 (.I(W14829), .ZN(O12337));
  INVX1 G34983 (.I(W2349), .ZN(O12338));
  INVX1 G34984 (.I(I110), .ZN(W8446));
  INVX1 G34985 (.I(I1316), .ZN(W8927));
  INVX1 G34986 (.I(W6499), .ZN(W8910));
  INVX1 G34987 (.I(W13800), .ZN(O12256));
  INVX1 G34988 (.I(W8785), .ZN(W8912));
  INVX1 G34989 (.I(W37958), .ZN(W42322));
  INVX1 G34990 (.I(I1906), .ZN(W45809));
  INVX1 G34991 (.I(I671), .ZN(W41990));
  INVX1 G34992 (.I(W21183), .ZN(O12258));
  INVX1 G34993 (.I(W4714), .ZN(W42327));
  INVX1 G34994 (.I(W3469), .ZN(W41986));
  INVX1 G34995 (.I(W18356), .ZN(O12261));
  INVX1 G34996 (.I(W33377), .ZN(O12262));
  INVX1 G34997 (.I(W36725), .ZN(O12001));
  INVX1 G34998 (.I(W28527), .ZN(W42320));
  INVX1 G34999 (.I(I393), .ZN(W8928));
  INVX1 G35000 (.I(W6848), .ZN(O11998));
  INVX1 G35001 (.I(W18957), .ZN(O12263));
  INVX1 G35002 (.I(W463), .ZN(W8563));
  INVX1 G35003 (.I(I770), .ZN(W8929));
  INVX1 G35004 (.I(I844), .ZN(W8562));
  INVX1 G35005 (.I(W24626), .ZN(W41976));
  INVX1 G35006 (.I(W18402), .ZN(O12267));
  INVX1 G35007 (.I(W3952), .ZN(W8558));
  INVX1 G35008 (.I(W2177), .ZN(W8555));
  INVX1 G35009 (.I(W525), .ZN(W8553));
  INVX1 G35010 (.I(I597), .ZN(O12011));
  INVX1 G35011 (.I(W11139), .ZN(O12018));
  INVX1 G35012 (.I(W4317), .ZN(W8900));
  INVX1 G35013 (.I(W5672), .ZN(W8592));
  INVX1 G35014 (.I(W941), .ZN(W42006));
  INVX1 G35015 (.I(W5218), .ZN(W8590));
  INVX1 G35016 (.I(W12038), .ZN(O12245));
  INVX1 G35017 (.I(W41453), .ZN(W42305));
  INVX1 G35018 (.I(W5137), .ZN(W8587));
  INVX1 G35019 (.I(I1710), .ZN(W8903));
  INVX1 G35020 (.I(W22253), .ZN(O12247));
  INVX1 G35021 (.I(W409), .ZN(O12012));
  INVX1 G35022 (.I(W4780), .ZN(W42311));
  INVX1 G35023 (.I(W6590), .ZN(W8552));
  INVX1 G35024 (.I(I785), .ZN(W8577));
  INVX1 G35025 (.I(W37090), .ZN(W41998));
  INVX1 G35026 (.I(W6443), .ZN(W8907));
  INVX1 G35027 (.I(W21639), .ZN(O12009));
  INVX1 G35028 (.I(W8454), .ZN(O12251));
  INVX1 G35029 (.I(W15785), .ZN(O12252));
  INVX1 G35030 (.I(W27747), .ZN(O12253));
  INVX1 G35031 (.I(W4313), .ZN(W8909));
  INVX1 G35032 (.I(W2448), .ZN(O12254));
  INVX1 G35033 (.I(W22647), .ZN(O12007));
  INVX1 G35034 (.I(W10294), .ZN(O12255));
  INVX1 G35035 (.I(W6217), .ZN(W8516));
  INVX1 G35036 (.I(W7851), .ZN(W8958));
  INVX1 G35037 (.I(W21998), .ZN(W42359));
  INVX1 G35038 (.I(W1273), .ZN(W8959));
  INVX1 G35039 (.I(I494), .ZN(W8529));
  INVX1 G35040 (.I(I1158), .ZN(W8963));
  INVX1 G35041 (.I(W29820), .ZN(W42362));
  INVX1 G35042 (.I(W34322), .ZN(W42363));
  INVX1 G35043 (.I(I848), .ZN(W8964));
  INVX1 G35044 (.I(W41273), .ZN(W42366));
  INVX1 G35045 (.I(W365), .ZN(W42367));
  INVX1 G35046 (.I(W12821), .ZN(W42369));
  INVX1 G35047 (.I(W38582), .ZN(O11972));
  INVX1 G35048 (.I(W3221), .ZN(W8531));
  INVX1 G35049 (.I(W2324), .ZN(W8512));
  INVX1 G35050 (.I(I1633), .ZN(W8511));
  INVX1 G35051 (.I(W4122), .ZN(W8509));
  INVX1 G35052 (.I(W3994), .ZN(W8968));
  INVX1 G35053 (.I(I71), .ZN(W8969));
  INVX1 G35054 (.I(W7764), .ZN(W8970));
  INVX1 G35055 (.I(W7662), .ZN(O12290));
  INVX1 G35056 (.I(I253), .ZN(W8972));
  INVX1 G35057 (.I(I495), .ZN(W8974));
  INVX1 G35058 (.I(W7022), .ZN(W8975));
  INVX1 G35059 (.I(W8047), .ZN(W8505));
  INVX1 G35060 (.I(W3980), .ZN(W8539));
  INVX1 G35061 (.I(W24083), .ZN(O12273));
  INVX1 G35062 (.I(W4739), .ZN(W8935));
  INVX1 G35063 (.I(W5551), .ZN(O256));
  INVX1 G35064 (.I(I781), .ZN(W8547));
  INVX1 G35065 (.I(W2542), .ZN(O11993));
  INVX1 G35066 (.I(W1974), .ZN(W8939));
  INVX1 G35067 (.I(W22817), .ZN(W42346));
  INVX1 G35068 (.I(W32875), .ZN(O12275));
  INVX1 G35069 (.I(I1985), .ZN(W8542));
  INVX1 G35070 (.I(W8722), .ZN(W8940));
  INVX1 G35071 (.I(I54), .ZN(W8941));
  INVX1 G35072 (.I(W7950), .ZN(W8942));
  INVX1 G35073 (.I(W40243), .ZN(O11728));
  INVX1 G35074 (.I(W5147), .ZN(W8945));
  INVX1 G35075 (.I(W8499), .ZN(O11985));
  INVX1 G35076 (.I(W5188), .ZN(W8535));
  INVX1 G35077 (.I(W29858), .ZN(O12279));
  INVX1 G35078 (.I(W45), .ZN(W42354));
  INVX1 G35079 (.I(W37928), .ZN(O12280));
  INVX1 G35080 (.I(I418), .ZN(O11982));
  INVX1 G35081 (.I(W7004), .ZN(W8948));
  INVX1 G35082 (.I(W5646), .ZN(W8951));
  INVX1 G35083 (.I(W4347), .ZN(O258));
  INVX1 G35084 (.I(I1523), .ZN(W8954));
  INVX1 G35085 (.I(W18791), .ZN(O11455));
  INVX1 G35086 (.I(W6055), .ZN(O11460));
  INVX1 G35087 (.I(W21230), .ZN(O12978));
  INVX1 G35088 (.I(W14015), .ZN(O12979));
  INVX1 G35089 (.I(W19973), .ZN(O11459));
  INVX1 G35090 (.I(I791), .ZN(W9692));
  INVX1 G35091 (.I(W7594), .ZN(W9693));
  INVX1 G35092 (.I(W8330), .ZN(O12980));
  INVX1 G35093 (.I(W284), .ZN(W7630));
  INVX1 G35094 (.I(W13360), .ZN(O12981));
  INVX1 G35095 (.I(W34431), .ZN(O12982));
  INVX1 G35096 (.I(W33274), .ZN(O11457));
  INVX1 G35097 (.I(W35037), .ZN(O11456));
  INVX1 G35098 (.I(W427), .ZN(W7631));
  INVX1 G35099 (.I(W35452), .ZN(O12985));
  INVX1 G35100 (.I(W493), .ZN(W9700));
  INVX1 G35101 (.I(W7336), .ZN(W41221));
  INVX1 G35102 (.I(W42945), .ZN(O12986));
  INVX1 G35103 (.I(W3612), .ZN(O316));
  INVX1 G35104 (.I(W1463), .ZN(W7627));
  INVX1 G35105 (.I(W3591), .ZN(W9704));
  INVX1 G35106 (.I(W6725), .ZN(W7626));
  INVX1 G35107 (.I(W6372), .ZN(W7625));
  INVX1 G35108 (.I(W25144), .ZN(O11446));
  INVX1 G35109 (.I(W3417), .ZN(W7623));
  INVX1 G35110 (.I(W26645), .ZN(O11443));
  INVX1 G35111 (.I(W1459), .ZN(W9673));
  INVX1 G35112 (.I(W3939), .ZN(W7658));
  INVX1 G35113 (.I(W1726), .ZN(W7657));
  INVX1 G35114 (.I(I1574), .ZN(W7655));
  INVX1 G35115 (.I(W9953), .ZN(O12963));
  INVX1 G35116 (.I(W32402), .ZN(W41248));
  INVX1 G35117 (.I(W36814), .ZN(O12964));
  INVX1 G35118 (.I(W318), .ZN(W7651));
  INVX1 G35119 (.I(W4748), .ZN(W7650));
  INVX1 G35120 (.I(W21695), .ZN(O11468));
  INVX1 G35121 (.I(W6289), .ZN(W7649));
  INVX1 G35122 (.I(W26146), .ZN(O12967));
  INVX1 G35123 (.I(I1342), .ZN(O315));
  INVX1 G35124 (.I(W3296), .ZN(W41210));
  INVX1 G35125 (.I(W4158), .ZN(W9674));
  INVX1 G35126 (.I(W5695), .ZN(W9676));
  INVX1 G35127 (.I(W13225), .ZN(W41242));
  INVX1 G35128 (.I(W3908), .ZN(W41241));
  INVX1 G35129 (.I(I190), .ZN(W9677));
  INVX1 G35130 (.I(W31505), .ZN(O11462));
  INVX1 G35131 (.I(I1826), .ZN(W9682));
  INVX1 G35132 (.I(W16969), .ZN(W43251));
  INVX1 G35133 (.I(W2528), .ZN(W7641));
  INVX1 G35134 (.I(W7516), .ZN(W7637));
  INVX1 G35135 (.I(W6171), .ZN(W7636));
  INVX1 G35136 (.I(W20227), .ZN(W41194));
  INVX1 G35137 (.I(W3192), .ZN(O13013));
  INVX1 G35138 (.I(I1727), .ZN(W9726));
  INVX1 G35139 (.I(W2647), .ZN(W7596));
  INVX1 G35140 (.I(W25136), .ZN(O13019));
  INVX1 G35141 (.I(W6079), .ZN(W7593));
  INVX1 G35142 (.I(W42921), .ZN(O13021));
  INVX1 G35143 (.I(W18069), .ZN(O13023));
  INVX1 G35144 (.I(W17668), .ZN(O11435));
  INVX1 G35145 (.I(W12092), .ZN(W43311));
  INVX1 G35146 (.I(W36587), .ZN(W41196));
  INVX1 G35147 (.I(I90), .ZN(W7587));
  INVX1 G35148 (.I(W8497), .ZN(W9730));
  INVX1 G35149 (.I(W24642), .ZN(O13012));
  INVX1 G35150 (.I(W40440), .ZN(W41193));
  INVX1 G35151 (.I(W3989), .ZN(W7586));
  INVX1 G35152 (.I(W1673), .ZN(W9731));
  INVX1 G35153 (.I(W7781), .ZN(W9733));
  INVX1 G35154 (.I(I1066), .ZN(O13028));
  INVX1 G35155 (.I(W31643), .ZN(W41190));
  INVX1 G35156 (.I(W2979), .ZN(W41189));
  INVX1 G35157 (.I(I1445), .ZN(W7581));
  INVX1 G35158 (.I(W7617), .ZN(W9734));
  INVX1 G35159 (.I(W3763), .ZN(W41187));
  INVX1 G35160 (.I(W3321), .ZN(W7579));
  INVX1 G35161 (.I(W22796), .ZN(O13004));
  INVX1 G35162 (.I(W4834), .ZN(W7622));
  INVX1 G35163 (.I(W13681), .ZN(O12993));
  INVX1 G35164 (.I(W1538), .ZN(O12994));
  INVX1 G35165 (.I(W416), .ZN(W9715));
  INVX1 G35166 (.I(W39762), .ZN(O12995));
  INVX1 G35167 (.I(W6846), .ZN(W7617));
  INVX1 G35168 (.I(W30649), .ZN(O12997));
  INVX1 G35169 (.I(W14997), .ZN(O11442));
  INVX1 G35170 (.I(W360), .ZN(W9716));
  INVX1 G35171 (.I(W4057), .ZN(W9717));
  INVX1 G35172 (.I(I1686), .ZN(W7613));
  INVX1 G35173 (.I(W867), .ZN(W7612));
  INVX1 G35174 (.I(I477), .ZN(W7660));
  INVX1 G35175 (.I(W6613), .ZN(W7609));
  INVX1 G35176 (.I(W18848), .ZN(O13005));
  INVX1 G35177 (.I(W4682), .ZN(W9722));
  INVX1 G35178 (.I(W8851), .ZN(O13006));
  INVX1 G35179 (.I(W34258), .ZN(W43291));
  INVX1 G35180 (.I(W40992), .ZN(O13008));
  INVX1 G35181 (.I(W2269), .ZN(W7605));
  INVX1 G35182 (.I(W28921), .ZN(O13010));
  INVX1 G35183 (.I(W13225), .ZN(O11438));
  INVX1 G35184 (.I(I1501), .ZN(W7604));
  INVX1 G35185 (.I(W26250), .ZN(W41201));
  INVX1 G35186 (.I(W8129), .ZN(O12913));
  INVX1 G35187 (.I(I1628), .ZN(O11496));
  INVX1 G35188 (.I(W17218), .ZN(O11495));
  INVX1 G35189 (.I(W26529), .ZN(O12903));
  INVX1 G35190 (.I(W3147), .ZN(W7719));
  INVX1 G35191 (.I(I1772), .ZN(W7717));
  INVX1 G35192 (.I(W16703), .ZN(O11494));
  INVX1 G35193 (.I(W35778), .ZN(O12908));
  INVX1 G35194 (.I(W7978), .ZN(O12909));
  INVX1 G35195 (.I(W17143), .ZN(O12910));
  INVX1 G35196 (.I(W4194), .ZN(W9622));
  INVX1 G35197 (.I(W767), .ZN(W43178));
  INVX1 G35198 (.I(W10191), .ZN(O12912));
  INVX1 G35199 (.I(W19289), .ZN(W41300));
  INVX1 G35200 (.I(W4026), .ZN(W9625));
  INVX1 G35201 (.I(W804), .ZN(W7712));
  INVX1 G35202 (.I(W7945), .ZN(W9627));
  INVX1 G35203 (.I(I1409), .ZN(O307));
  INVX1 G35204 (.I(W26571), .ZN(O12915));
  INVX1 G35205 (.I(W4229), .ZN(W7711));
  INVX1 G35206 (.I(W40107), .ZN(W41284));
  INVX1 G35207 (.I(W3008), .ZN(W9629));
  INVX1 G35208 (.I(W2680), .ZN(O196));
  INVX1 G35209 (.I(I1514), .ZN(W7706));
  INVX1 G35210 (.I(W9545), .ZN(W41281));
  INVX1 G35211 (.I(W4820), .ZN(O12893));
  INVX1 G35212 (.I(W1923), .ZN(O12885));
  INVX1 G35213 (.I(W810), .ZN(W41316));
  INVX1 G35214 (.I(W15866), .ZN(O12887));
  INVX1 G35215 (.I(W28605), .ZN(O12888));
  INVX1 G35216 (.I(W8169), .ZN(W9605));
  INVX1 G35217 (.I(W29772), .ZN(O12889));
  INVX1 G35218 (.I(W36400), .ZN(W41314));
  INVX1 G35219 (.I(W5895), .ZN(W7735));
  INVX1 G35220 (.I(W455), .ZN(O11507));
  INVX1 G35221 (.I(W32689), .ZN(O11506));
  INVX1 G35222 (.I(W4080), .ZN(W7732));
  INVX1 G35223 (.I(W3522), .ZN(O11505));
  INVX1 G35224 (.I(W4741), .ZN(W9631));
  INVX1 G35225 (.I(I539), .ZN(O11504));
  INVX1 G35226 (.I(W4957), .ZN(W7729));
  INVX1 G35227 (.I(I1033), .ZN(W7727));
  INVX1 G35228 (.I(W41185), .ZN(O12897));
  INVX1 G35229 (.I(I172), .ZN(W9607));
  INVX1 G35230 (.I(W166), .ZN(W9610));
  INVX1 G35231 (.I(W39897), .ZN(O11501));
  INVX1 G35232 (.I(W25795), .ZN(W41305));
  INVX1 G35233 (.I(W6753), .ZN(W7725));
  INVX1 G35234 (.I(W20177), .ZN(O11500));
  INVX1 G35235 (.I(W20587), .ZN(W41302));
  INVX1 G35236 (.I(W41894), .ZN(W43221));
  INVX1 G35237 (.I(W4342), .ZN(W9651));
  INVX1 G35238 (.I(W7375), .ZN(W9652));
  INVX1 G35239 (.I(W5708), .ZN(W7687));
  INVX1 G35240 (.I(W9384), .ZN(O12942));
  INVX1 G35241 (.I(W3346), .ZN(W7681));
  INVX1 G35242 (.I(W2797), .ZN(W9657));
  INVX1 G35243 (.I(W33402), .ZN(O12944));
  INVX1 G35244 (.I(W6156), .ZN(O313));
  INVX1 G35245 (.I(W3999), .ZN(O12945));
  INVX1 G35246 (.I(W4812), .ZN(O11475));
  INVX1 G35247 (.I(W982), .ZN(O314));
  INVX1 G35248 (.I(W9413), .ZN(W41256));
  INVX1 G35249 (.I(W36929), .ZN(O12938));
  INVX1 G35250 (.I(I520), .ZN(W7677));
  INVX1 G35251 (.I(W9399), .ZN(W9663));
  INVX1 G35252 (.I(W7578), .ZN(O193));
  INVX1 G35253 (.I(W7249), .ZN(W9666));
  INVX1 G35254 (.I(W7396), .ZN(W7672));
  INVX1 G35255 (.I(W29958), .ZN(O12950));
  INVX1 G35256 (.I(W25550), .ZN(W41251));
  INVX1 G35257 (.I(W3823), .ZN(W7670));
  INVX1 G35258 (.I(I1580), .ZN(W7668));
  INVX1 G35259 (.I(W6570), .ZN(W7667));
  INVX1 G35260 (.I(W4307), .ZN(O192));
  INVX1 G35261 (.I(W10173), .ZN(O12927));
  INVX1 G35262 (.I(W8415), .ZN(W41279));
  INVX1 G35263 (.I(I386), .ZN(W7705));
  INVX1 G35264 (.I(W21065), .ZN(W41278));
  INVX1 G35265 (.I(W3217), .ZN(O12920));
  INVX1 G35266 (.I(W6769), .ZN(W9632));
  INVX1 G35267 (.I(W3059), .ZN(W9636));
  INVX1 G35268 (.I(W32351), .ZN(O12922));
  INVX1 G35269 (.I(W5494), .ZN(O12924));
  INVX1 G35270 (.I(W4635), .ZN(W41273));
  INVX1 G35271 (.I(W23810), .ZN(O11484));
  INVX1 G35272 (.I(I1575), .ZN(W9641));
  INVX1 G35273 (.I(W6720), .ZN(W9644));
  INVX1 G35274 (.I(W40830), .ZN(W41186));
  INVX1 G35275 (.I(W17335), .ZN(O12928));
  INVX1 G35276 (.I(W27367), .ZN(O11482));
  INVX1 G35277 (.I(W6483), .ZN(W9646));
  INVX1 G35278 (.I(W27460), .ZN(O12930));
  INVX1 G35279 (.I(I1014), .ZN(W43200));
  INVX1 G35280 (.I(W10960), .ZN(O12931));
  INVX1 G35281 (.I(I540), .ZN(W7692));
  INVX1 G35282 (.I(W35210), .ZN(O12935));
  INVX1 G35283 (.I(W1361), .ZN(O12936));
  INVX1 G35284 (.I(W361), .ZN(W9649));
  INVX1 G35285 (.I(W3923), .ZN(W7690));
  INVX1 G35286 (.I(W7794), .ZN(W9799));
  INVX1 G35287 (.I(W15192), .ZN(W41110));
  INVX1 G35288 (.I(W2744), .ZN(W7495));
  INVX1 G35289 (.I(W1663), .ZN(O13100));
  INVX1 G35290 (.I(W27769), .ZN(O13101));
  INVX1 G35291 (.I(W24030), .ZN(O13102));
  INVX1 G35292 (.I(W36071), .ZN(O13103));
  INVX1 G35293 (.I(W39022), .ZN(O11375));
  INVX1 G35294 (.I(I1122), .ZN(O11374));
  INVX1 G35295 (.I(W20447), .ZN(O11373));
  INVX1 G35296 (.I(W1645), .ZN(W7493));
  INVX1 G35297 (.I(W7102), .ZN(W7491));
  INVX1 G35298 (.I(W1993), .ZN(W41106));
  INVX1 G35299 (.I(W5821), .ZN(W7496));
  INVX1 G35300 (.I(W7066), .ZN(W7483));
  INVX1 G35301 (.I(I39), .ZN(W41104));
  INVX1 G35302 (.I(W11900), .ZN(O11371));
  INVX1 G35303 (.I(I1245), .ZN(W7480));
  INVX1 G35304 (.I(W7227), .ZN(W43417));
  INVX1 G35305 (.I(W6795), .ZN(O13109));
  INVX1 G35306 (.I(W2188), .ZN(W9800));
  INVX1 G35307 (.I(W3938), .ZN(W7476));
  INVX1 G35308 (.I(W6230), .ZN(O328));
  INVX1 G35309 (.I(W14067), .ZN(O11368));
  INVX1 G35310 (.I(I1880), .ZN(W7475));
  INVX1 G35311 (.I(W4534), .ZN(O11379));
  INVX1 G35312 (.I(W9669), .ZN(W9784));
  INVX1 G35313 (.I(W5538), .ZN(W9785));
  INVX1 G35314 (.I(W26462), .ZN(O11385));
  INVX1 G35315 (.I(I1562), .ZN(W9787));
  INVX1 G35316 (.I(W12219), .ZN(O11383));
  INVX1 G35317 (.I(W6159), .ZN(O324));
  INVX1 G35318 (.I(W114), .ZN(W7510));
  INVX1 G35319 (.I(W23512), .ZN(O11381));
  INVX1 G35320 (.I(I501), .ZN(O325));
  INVX1 G35321 (.I(W4622), .ZN(W7507));
  INVX1 G35322 (.I(I1856), .ZN(W9792));
  INVX1 G35323 (.I(W21582), .ZN(W43394));
  INVX1 G35324 (.I(W117), .ZN(W7474));
  INVX1 G35325 (.I(W3829), .ZN(W7504));
  INVX1 G35326 (.I(W5971), .ZN(W7503));
  INVX1 G35327 (.I(I166), .ZN(W7501));
  INVX1 G35328 (.I(W5558), .ZN(W7500));
  INVX1 G35329 (.I(W6151), .ZN(W9793));
  INVX1 G35330 (.I(W32942), .ZN(O13095));
  INVX1 G35331 (.I(W12604), .ZN(O13096));
  INVX1 G35332 (.I(W1459), .ZN(O11378));
  INVX1 G35333 (.I(W5987), .ZN(W9795));
  INVX1 G35334 (.I(W4840), .ZN(W7497));
  INVX1 G35335 (.I(W3609), .ZN(O13098));
  INVX1 G35336 (.I(I1663), .ZN(O11351));
  INVX1 G35337 (.I(W25012), .ZN(O11356));
  INVX1 G35338 (.I(W18098), .ZN(O13127));
  INVX1 G35339 (.I(W5352), .ZN(W7451));
  INVX1 G35340 (.I(W28429), .ZN(O11355));
  INVX1 G35341 (.I(W6067), .ZN(W9815));
  INVX1 G35342 (.I(W25470), .ZN(O11353));
  INVX1 G35343 (.I(W24633), .ZN(O13130));
  INVX1 G35344 (.I(W6943), .ZN(W7449));
  INVX1 G35345 (.I(W35732), .ZN(W43448));
  INVX1 G35346 (.I(I1461), .ZN(O11352));
  INVX1 G35347 (.I(W1257), .ZN(W7447));
  INVX1 G35348 (.I(W36579), .ZN(O13134));
  INVX1 G35349 (.I(W20986), .ZN(O13126));
  INVX1 G35350 (.I(W32882), .ZN(O13135));
  INVX1 G35351 (.I(W559), .ZN(W7446));
  INVX1 G35352 (.I(W6813), .ZN(W9816));
  INVX1 G35353 (.I(W2470), .ZN(W7444));
  INVX1 G35354 (.I(W2967), .ZN(W9819));
  INVX1 G35355 (.I(W18268), .ZN(O13138));
  INVX1 G35356 (.I(W6737), .ZN(W7441));
  INVX1 G35357 (.I(W33045), .ZN(O13140));
  INVX1 G35358 (.I(W6520), .ZN(W7439));
  INVX1 G35359 (.I(W5829), .ZN(O183));
  INVX1 G35360 (.I(W21723), .ZN(W41076));
  INVX1 G35361 (.I(W31633), .ZN(W43432));
  INVX1 G35362 (.I(W6282), .ZN(W9805));
  INVX1 G35363 (.I(W8454), .ZN(W9806));
  INVX1 G35364 (.I(W5956), .ZN(W7473));
  INVX1 G35365 (.I(I1435), .ZN(W7472));
  INVX1 G35366 (.I(W5603), .ZN(W7471));
  INVX1 G35367 (.I(W1184), .ZN(W7470));
  INVX1 G35368 (.I(W17687), .ZN(O11365));
  INVX1 G35369 (.I(I1156), .ZN(W7467));
  INVX1 G35370 (.I(W8157), .ZN(W41095));
  INVX1 G35371 (.I(W26597), .ZN(O11363));
  INVX1 G35372 (.I(W597), .ZN(O13119));
  INVX1 G35373 (.I(W23517), .ZN(W43431));
  INVX1 G35374 (.I(W3638), .ZN(W9783));
  INVX1 G35375 (.I(W4168), .ZN(W9811));
  INVX1 G35376 (.I(W5433), .ZN(W7464));
  INVX1 G35377 (.I(W28858), .ZN(O11361));
  INVX1 G35378 (.I(W5872), .ZN(W7463));
  INVX1 G35379 (.I(W17533), .ZN(W41091));
  INVX1 G35380 (.I(W2654), .ZN(W9812));
  INVX1 G35381 (.I(W31444), .ZN(O11359));
  INVX1 G35382 (.I(W983), .ZN(W7456));
  INVX1 G35383 (.I(W35199), .ZN(O11358));
  INVX1 G35384 (.I(W13346), .ZN(O11357));
  INVX1 G35385 (.I(W14257), .ZN(O13125));
  INVX1 G35386 (.I(W3410), .ZN(O13056));
  INVX1 G35387 (.I(W32164), .ZN(W41171));
  INVX1 G35388 (.I(W36241), .ZN(W41170));
  INVX1 G35389 (.I(W3585), .ZN(W7556));
  INVX1 G35390 (.I(W7000), .ZN(O11421));
  INVX1 G35391 (.I(W2143), .ZN(W7555));
  INVX1 G35392 (.I(W6238), .ZN(W7554));
  INVX1 G35393 (.I(W5100), .ZN(W7553));
  INVX1 G35394 (.I(W19636), .ZN(O11419));
  INVX1 G35395 (.I(W3930), .ZN(W7552));
  INVX1 G35396 (.I(W6082), .ZN(W9749));
  INVX1 G35397 (.I(W10625), .ZN(W41164));
  INVX1 G35398 (.I(W13985), .ZN(W43344));
  INVX1 G35399 (.I(W890), .ZN(W7558));
  INVX1 G35400 (.I(W20906), .ZN(O11416));
  INVX1 G35401 (.I(W2003), .ZN(W9751));
  INVX1 G35402 (.I(W33541), .ZN(O13057));
  INVX1 G35403 (.I(W18167), .ZN(O13058));
  INVX1 G35404 (.I(I1617), .ZN(W7548));
  INVX1 G35405 (.I(W20782), .ZN(W41160));
  INVX1 G35406 (.I(W1132), .ZN(O11414));
  INVX1 G35407 (.I(W1601), .ZN(W7547));
  INVX1 G35408 (.I(W40902), .ZN(O11412));
  INVX1 G35409 (.I(W10537), .ZN(W43352));
  INVX1 G35410 (.I(I544), .ZN(W7544));
  INVX1 G35411 (.I(W2521), .ZN(W7569));
  INVX1 G35412 (.I(W18095), .ZN(O13031));
  INVX1 G35413 (.I(W10130), .ZN(W41185));
  INVX1 G35414 (.I(W4425), .ZN(O321));
  INVX1 G35415 (.I(W3150), .ZN(W9736));
  INVX1 G35416 (.I(W36779), .ZN(W41182));
  INVX1 G35417 (.I(I1486), .ZN(W7574));
  INVX1 G35418 (.I(W28696), .ZN(O13035));
  INVX1 G35419 (.I(I91), .ZN(W7571));
  INVX1 G35420 (.I(W1314), .ZN(W9739));
  INVX1 G35421 (.I(W20416), .ZN(O11426));
  INVX1 G35422 (.I(W6609), .ZN(W9740));
  INVX1 G35423 (.I(W6101), .ZN(W9741));
  INVX1 G35424 (.I(W3034), .ZN(W9759));
  INVX1 G35425 (.I(W2908), .ZN(W9742));
  INVX1 G35426 (.I(W405), .ZN(W7567));
  INVX1 G35427 (.I(W10464), .ZN(O13040));
  INVX1 G35428 (.I(W6305), .ZN(W9744));
  INVX1 G35429 (.I(W6725), .ZN(W7565));
  INVX1 G35430 (.I(I1758), .ZN(W7564));
  INVX1 G35431 (.I(W7124), .ZN(W7562));
  INVX1 G35432 (.I(I1600), .ZN(O13045));
  INVX1 G35433 (.I(W1037), .ZN(W7561));
  INVX1 G35434 (.I(W15977), .ZN(O11422));
  INVX1 G35435 (.I(W10875), .ZN(O13047));
  INVX1 G35436 (.I(W29961), .ZN(O11395));
  INVX1 G35437 (.I(W30365), .ZN(O13080));
  INVX1 G35438 (.I(W5379), .ZN(W9764));
  INVX1 G35439 (.I(W9084), .ZN(W9765));
  INVX1 G35440 (.I(W4512), .ZN(W9766));
  INVX1 G35441 (.I(W1349), .ZN(W7524));
  INVX1 G35442 (.I(W16254), .ZN(O11400));
  INVX1 G35443 (.I(W34475), .ZN(O13081));
  INVX1 G35444 (.I(I1350), .ZN(O323));
  INVX1 G35445 (.I(W961), .ZN(W7520));
  INVX1 G35446 (.I(W8352), .ZN(O13084));
  INVX1 G35447 (.I(W16416), .ZN(O11397));
  INVX1 G35448 (.I(W28042), .ZN(O11396));
  INVX1 G35449 (.I(W4181), .ZN(W7525));
  INVX1 G35450 (.I(W33760), .ZN(O13086));
  INVX1 G35451 (.I(W1854), .ZN(W9772));
  INVX1 G35452 (.I(W56), .ZN(W7516));
  INVX1 G35453 (.I(W2921), .ZN(W9773));
  INVX1 G35454 (.I(W16930), .ZN(O11392));
  INVX1 G35455 (.I(W7900), .ZN(W9774));
  INVX1 G35456 (.I(W450), .ZN(W43386));
  INVX1 G35457 (.I(W5040), .ZN(W9780));
  INVX1 G35458 (.I(W22465), .ZN(W43389));
  INVX1 G35459 (.I(W6628), .ZN(W9782));
  INVX1 G35460 (.I(W20490), .ZN(W41127));
  INVX1 G35461 (.I(W14433), .ZN(O11405));
  INVX1 G35462 (.I(W6720), .ZN(W7543));
  INVX1 G35463 (.I(W1870), .ZN(W7542));
  INVX1 G35464 (.I(W11909), .ZN(O11409));
  INVX1 G35465 (.I(W13985), .ZN(W41152));
  INVX1 G35466 (.I(W34000), .ZN(O13066));
  INVX1 G35467 (.I(W5733), .ZN(W7539));
  INVX1 G35468 (.I(W24335), .ZN(O13068));
  INVX1 G35469 (.I(W2652), .ZN(O11407));
  INVX1 G35470 (.I(W5298), .ZN(W7537));
  INVX1 G35471 (.I(W6886), .ZN(W9761));
  INVX1 G35472 (.I(W11830), .ZN(O11406));
  INVX1 G35473 (.I(W4971), .ZN(W7536));
  INVX1 G35474 (.I(W6275), .ZN(W9602));
  INVX1 G35475 (.I(W24946), .ZN(W43365));
  INVX1 G35476 (.I(W36846), .ZN(O13072));
  INVX1 G35477 (.I(W5719), .ZN(W7533));
  INVX1 G35478 (.I(I1678), .ZN(W7532));
  INVX1 G35479 (.I(W17231), .ZN(W43369));
  INVX1 G35480 (.I(W15581), .ZN(O13075));
  INVX1 G35481 (.I(W32902), .ZN(O11404));
  INVX1 G35482 (.I(W3050), .ZN(W7530));
  INVX1 G35483 (.I(I17), .ZN(W7528));
  INVX1 G35484 (.I(I665), .ZN(W9763));
  INVX1 G35485 (.I(W2206), .ZN(W7526));
  INVX1 G35486 (.I(W9506), .ZN(W41517));
  INVX1 G35487 (.I(W6451), .ZN(O11664));
  INVX1 G35488 (.I(W11042), .ZN(O12706));
  INVX1 G35489 (.I(W3687), .ZN(W7976));
  INVX1 G35490 (.I(W34565), .ZN(O12708));
  INVX1 G35491 (.I(W23660), .ZN(O12709));
  INVX1 G35492 (.I(W19761), .ZN(O12710));
  INVX1 G35493 (.I(W15953), .ZN(W42918));
  INVX1 G35494 (.I(W3512), .ZN(O206));
  INVX1 G35495 (.I(W1908), .ZN(W7974));
  INVX1 G35496 (.I(W24923), .ZN(W42921));
  INVX1 G35497 (.I(W376), .ZN(W9411));
  INVX1 G35498 (.I(W3920), .ZN(O12713));
  INVX1 G35499 (.I(W109), .ZN(W9408));
  INVX1 G35500 (.I(W22065), .ZN(O11657));
  INVX1 G35501 (.I(W8062), .ZN(O11656));
  INVX1 G35502 (.I(W22555), .ZN(O11655));
  INVX1 G35503 (.I(W37964), .ZN(O12716));
  INVX1 G35504 (.I(W26180), .ZN(O12717));
  INVX1 G35505 (.I(W30070), .ZN(O12718));
  INVX1 G35506 (.I(W8248), .ZN(W9421));
  INVX1 G35507 (.I(I1367), .ZN(W7965));
  INVX1 G35508 (.I(W2330), .ZN(W9422));
  INVX1 G35509 (.I(W21773), .ZN(O12721));
  INVX1 G35510 (.I(W40266), .ZN(O12723));
  INVX1 G35511 (.I(W12677), .ZN(O11651));
  INVX1 G35512 (.I(W12), .ZN(W9394));
  INVX1 G35513 (.I(W2297), .ZN(W8000));
  INVX1 G35514 (.I(W8293), .ZN(W9386));
  INVX1 G35515 (.I(W39800), .ZN(O12692));
  INVX1 G35516 (.I(W2121), .ZN(O11680));
  INVX1 G35517 (.I(W3438), .ZN(W42895));
  INVX1 G35518 (.I(W1770), .ZN(W9387));
  INVX1 G35519 (.I(W30441), .ZN(O12693));
  INVX1 G35520 (.I(W495), .ZN(W9391));
  INVX1 G35521 (.I(W29409), .ZN(W42898));
  INVX1 G35522 (.I(I1681), .ZN(W9393));
  INVX1 G35523 (.I(W6172), .ZN(W7992));
  INVX1 G35524 (.I(W23158), .ZN(O11676));
  INVX1 G35525 (.I(W2110), .ZN(W7961));
  INVX1 G35526 (.I(W4741), .ZN(O11675));
  INVX1 G35527 (.I(W34569), .ZN(O12697));
  INVX1 G35528 (.I(W3649), .ZN(W9398));
  INVX1 G35529 (.I(W30743), .ZN(O11672));
  INVX1 G35530 (.I(W2716), .ZN(W7986));
  INVX1 G35531 (.I(W348), .ZN(W9403));
  INVX1 G35532 (.I(W9334), .ZN(O11669));
  INVX1 G35533 (.I(I1306), .ZN(O12702));
  INVX1 G35534 (.I(W2914), .ZN(W9404));
  INVX1 G35535 (.I(I172), .ZN(W41526));
  INVX1 G35536 (.I(W5069), .ZN(W7979));
  INVX1 G35537 (.I(W3015), .ZN(W7924));
  INVX1 G35538 (.I(W6585), .ZN(W7936));
  INVX1 G35539 (.I(W5301), .ZN(W9440));
  INVX1 G35540 (.I(W880), .ZN(W7934));
  INVX1 G35541 (.I(W2553), .ZN(W7933));
  INVX1 G35542 (.I(W29110), .ZN(O12744));
  INVX1 G35543 (.I(W30047), .ZN(O12745));
  INVX1 G35544 (.I(W33396), .ZN(W41485));
  INVX1 G35545 (.I(W2815), .ZN(W7931));
  INVX1 G35546 (.I(W32811), .ZN(O11635));
  INVX1 G35547 (.I(W7634), .ZN(W7928));
  INVX1 G35548 (.I(W327), .ZN(W7926));
  INVX1 G35549 (.I(W14599), .ZN(O12748));
  INVX1 G35550 (.I(W23114), .ZN(O12740));
  INVX1 G35551 (.I(W37898), .ZN(O12750));
  INVX1 G35552 (.I(W28499), .ZN(O12751));
  INVX1 G35553 (.I(I376), .ZN(W7923));
  INVX1 G35554 (.I(W753), .ZN(W9456));
  INVX1 G35555 (.I(W31022), .ZN(O12752));
  INVX1 G35556 (.I(W14754), .ZN(O12753));
  INVX1 G35557 (.I(W29363), .ZN(O12754));
  INVX1 G35558 (.I(W14716), .ZN(W41478));
  INVX1 G35559 (.I(I5), .ZN(W9457));
  INVX1 G35560 (.I(I1719), .ZN(O292));
  INVX1 G35561 (.I(W8795), .ZN(W9459));
  INVX1 G35562 (.I(W6309), .ZN(W42950));
  INVX1 G35563 (.I(W3812), .ZN(W9424));
  INVX1 G35564 (.I(W1704), .ZN(W7959));
  INVX1 G35565 (.I(W40128), .ZN(O12727));
  INVX1 G35566 (.I(W31881), .ZN(O12729));
  INVX1 G35567 (.I(W27340), .ZN(O11648));
  INVX1 G35568 (.I(W5554), .ZN(W7954));
  INVX1 G35569 (.I(W25635), .ZN(O11647));
  INVX1 G35570 (.I(W1664), .ZN(W42945));
  INVX1 G35571 (.I(W32242), .ZN(O11645));
  INVX1 G35572 (.I(W18277), .ZN(W41499));
  INVX1 G35573 (.I(W5275), .ZN(W7944));
  INVX1 G35574 (.I(W6268), .ZN(W9434));
  INVX1 G35575 (.I(W6918), .ZN(W8001));
  INVX1 G35576 (.I(W33101), .ZN(O12735));
  INVX1 G35577 (.I(W36381), .ZN(O12736));
  INVX1 G35578 (.I(W197), .ZN(O11643));
  INVX1 G35579 (.I(I1679), .ZN(W7942));
  INVX1 G35580 (.I(I1463), .ZN(W7940));
  INVX1 G35581 (.I(W2817), .ZN(W9436));
  INVX1 G35582 (.I(W8267), .ZN(W9438));
  INVX1 G35583 (.I(W34479), .ZN(O11640));
  INVX1 G35584 (.I(W39555), .ZN(W41492));
  INVX1 G35585 (.I(W39636), .ZN(O12739));
  INVX1 G35586 (.I(W8759), .ZN(W9439));
  INVX1 G35587 (.I(W2840), .ZN(W8041));
  INVX1 G35588 (.I(W31569), .ZN(W42833));
  INVX1 G35589 (.I(W25186), .ZN(O12648));
  INVX1 G35590 (.I(W2149), .ZN(W9344));
  INVX1 G35591 (.I(W24746), .ZN(O12649));
  INVX1 G35592 (.I(I992), .ZN(W8048));
  INVX1 G35593 (.I(W999), .ZN(W8047));
  INVX1 G35594 (.I(W21435), .ZN(W42841));
  INVX1 G35595 (.I(W7959), .ZN(W8045));
  INVX1 G35596 (.I(W688), .ZN(W8044));
  INVX1 G35597 (.I(W4260), .ZN(W9346));
  INVX1 G35598 (.I(W30063), .ZN(O11711));
  INVX1 G35599 (.I(I1053), .ZN(W8042));
  INVX1 G35600 (.I(W34207), .ZN(O11713));
  INVX1 G35601 (.I(W38771), .ZN(O11710));
  INVX1 G35602 (.I(W5313), .ZN(W9347));
  INVX1 G35603 (.I(W1658), .ZN(W9349));
  INVX1 G35604 (.I(W7222), .ZN(W42847));
  INVX1 G35605 (.I(W7438), .ZN(O12658));
  INVX1 G35606 (.I(W906), .ZN(W8039));
  INVX1 G35607 (.I(I301), .ZN(W9350));
  INVX1 G35608 (.I(W1987), .ZN(W9351));
  INVX1 G35609 (.I(W859), .ZN(W8038));
  INVX1 G35610 (.I(W4242), .ZN(W9353));
  INVX1 G35611 (.I(W8791), .ZN(W9354));
  INVX1 G35612 (.I(W13311), .ZN(O12637));
  INVX1 G35613 (.I(W37798), .ZN(O12629));
  INVX1 G35614 (.I(I1958), .ZN(W9330));
  INVX1 G35615 (.I(W136), .ZN(W9331));
  INVX1 G35616 (.I(W7719), .ZN(W9333));
  INVX1 G35617 (.I(W32783), .ZN(O12632));
  INVX1 G35618 (.I(W36318), .ZN(O11724));
  INVX1 G35619 (.I(W38389), .ZN(O12634));
  INVX1 G35620 (.I(I1213), .ZN(W8068));
  INVX1 G35621 (.I(W5064), .ZN(W41601));
  INVX1 G35622 (.I(I303), .ZN(O12636));
  INVX1 G35623 (.I(W1803), .ZN(W9335));
  INVX1 G35624 (.I(W2751), .ZN(O11722));
  INVX1 G35625 (.I(W6080), .ZN(W8035));
  INVX1 G35626 (.I(W2837), .ZN(W8065));
  INVX1 G35627 (.I(W1307), .ZN(W9336));
  INVX1 G35628 (.I(W3453), .ZN(W9339));
  INVX1 G35629 (.I(W17304), .ZN(O11717));
  INVX1 G35630 (.I(W5908), .ZN(W8061));
  INVX1 G35631 (.I(W3793), .ZN(W8060));
  INVX1 G35632 (.I(W2270), .ZN(O12643));
  INVX1 G35633 (.I(W3984), .ZN(W8054));
  INVX1 G35634 (.I(W1570), .ZN(W9342));
  INVX1 G35635 (.I(I1807), .ZN(W42831));
  INVX1 G35636 (.I(W1137), .ZN(O12647));
  INVX1 G35637 (.I(W473), .ZN(W8009));
  INVX1 G35638 (.I(W14181), .ZN(O12677));
  INVX1 G35639 (.I(I232), .ZN(W8016));
  INVX1 G35640 (.I(W8157), .ZN(W41565));
  INVX1 G35641 (.I(I1459), .ZN(W8015));
  INVX1 G35642 (.I(W5475), .ZN(W9368));
  INVX1 G35643 (.I(W744), .ZN(O11694));
  INVX1 G35644 (.I(W7002), .ZN(W9369));
  INVX1 G35645 (.I(W2696), .ZN(W8011));
  INVX1 G35646 (.I(W3875), .ZN(O11693));
  INVX1 G35647 (.I(W6194), .ZN(W9370));
  INVX1 G35648 (.I(W4328), .ZN(W9371));
  INVX1 G35649 (.I(W2862), .ZN(W9372));
  INVX1 G35650 (.I(W40552), .ZN(O12676));
  INVX1 G35651 (.I(W5146), .ZN(W8008));
  INVX1 G35652 (.I(W3453), .ZN(O11688));
  INVX1 G35653 (.I(W5767), .ZN(W8007));
  INVX1 G35654 (.I(W6609), .ZN(W9375));
  INVX1 G35655 (.I(I559), .ZN(O11686));
  INVX1 G35656 (.I(W5671), .ZN(W9377));
  INVX1 G35657 (.I(W28029), .ZN(O12687));
  INVX1 G35658 (.I(W8956), .ZN(W9382));
  INVX1 G35659 (.I(I941), .ZN(O11682));
  INVX1 G35660 (.I(W3851), .ZN(W8002));
  INVX1 G35661 (.I(W10300), .ZN(W42889));
  INVX1 G35662 (.I(W7314), .ZN(W8029));
  INVX1 G35663 (.I(W5479), .ZN(W8034));
  INVX1 G35664 (.I(W37620), .ZN(W42854));
  INVX1 G35665 (.I(I158), .ZN(W8032));
  INVX1 G35666 (.I(W23541), .ZN(O12665));
  INVX1 G35667 (.I(W2208), .ZN(W9355));
  INVX1 G35668 (.I(W6829), .ZN(O209));
  INVX1 G35669 (.I(W32573), .ZN(O12667));
  INVX1 G35670 (.I(W25960), .ZN(W42860));
  INVX1 G35671 (.I(W7701), .ZN(O12668));
  INVX1 G35672 (.I(W11036), .ZN(W41575));
  INVX1 G35673 (.I(W3835), .ZN(W9357));
  INVX1 G35674 (.I(W13394), .ZN(W42862));
  INVX1 G35675 (.I(W3236), .ZN(W7922));
  INVX1 G35676 (.I(W13973), .ZN(W41573));
  INVX1 G35677 (.I(W5839), .ZN(W8025));
  INVX1 G35678 (.I(W3224), .ZN(W9359));
  INVX1 G35679 (.I(W3209), .ZN(W9362));
  INVX1 G35680 (.I(W36790), .ZN(O12672));
  INVX1 G35681 (.I(I1181), .ZN(W9364));
  INVX1 G35682 (.I(W19140), .ZN(O12673));
  INVX1 G35683 (.I(W29259), .ZN(W42869));
  INVX1 G35684 (.I(W3846), .ZN(W8023));
  INVX1 G35685 (.I(W1462), .ZN(W8022));
  INVX1 G35686 (.I(W6847), .ZN(W8019));
  INVX1 G35687 (.I(W38920), .ZN(O12847));
  INVX1 G35688 (.I(W10965), .ZN(W41370));
  INVX1 G35689 (.I(W6871), .ZN(W7806));
  INVX1 G35690 (.I(W24627), .ZN(O11553));
  INVX1 G35691 (.I(W2125), .ZN(O12839));
  INVX1 G35692 (.I(W13579), .ZN(O12840));
  INVX1 G35693 (.I(W28145), .ZN(O11550));
  INVX1 G35694 (.I(W7015), .ZN(W7803));
  INVX1 G35695 (.I(W1716), .ZN(W41365));
  INVX1 G35696 (.I(W2418), .ZN(O11549));
  INVX1 G35697 (.I(W4549), .ZN(W7801));
  INVX1 G35698 (.I(W2733), .ZN(W7798));
  INVX1 G35699 (.I(W17747), .ZN(O12846));
  INVX1 G35700 (.I(W2957), .ZN(W7807));
  INVX1 G35701 (.I(W32211), .ZN(O11546));
  INVX1 G35702 (.I(W24110), .ZN(W41359));
  INVX1 G35703 (.I(W4945), .ZN(W7796));
  INVX1 G35704 (.I(W22126), .ZN(W43094));
  INVX1 G35705 (.I(W12048), .ZN(W43095));
  INVX1 G35706 (.I(W7273), .ZN(W7795));
  INVX1 G35707 (.I(W1394), .ZN(W7794));
  INVX1 G35708 (.I(W42108), .ZN(O12851));
  INVX1 G35709 (.I(W7314), .ZN(W9566));
  INVX1 G35710 (.I(W10703), .ZN(W41356));
  INVX1 G35711 (.I(I827), .ZN(O11543));
  INVX1 G35712 (.I(W7563), .ZN(O11560));
  INVX1 G35713 (.I(W3636), .ZN(O12817));
  INVX1 G35714 (.I(W5809), .ZN(W9540));
  INVX1 G35715 (.I(I1244), .ZN(W9541));
  INVX1 G35716 (.I(W6042), .ZN(W7828));
  INVX1 G35717 (.I(I165), .ZN(W9546));
  INVX1 G35718 (.I(W5306), .ZN(W7827));
  INVX1 G35719 (.I(W22779), .ZN(W43062));
  INVX1 G35720 (.I(I148), .ZN(W7826));
  INVX1 G35721 (.I(W2590), .ZN(W9547));
  INVX1 G35722 (.I(I1703), .ZN(O12822));
  INVX1 G35723 (.I(W19122), .ZN(O12823));
  INVX1 G35724 (.I(I872), .ZN(W9549));
  INVX1 G35725 (.I(W15215), .ZN(O12859));
  INVX1 G35726 (.I(W18414), .ZN(O11559));
  INVX1 G35727 (.I(W34251), .ZN(O12825));
  INVX1 G35728 (.I(W37015), .ZN(O12827));
  INVX1 G35729 (.I(W41280), .ZN(O11557));
  INVX1 G35730 (.I(W1856), .ZN(W9555));
  INVX1 G35731 (.I(I1963), .ZN(W7815));
  INVX1 G35732 (.I(W3161), .ZN(W9556));
  INVX1 G35733 (.I(W18084), .ZN(O11554));
  INVX1 G35734 (.I(W14015), .ZN(O12834));
  INVX1 G35735 (.I(W17), .ZN(W7808));
  INVX1 G35736 (.I(W17284), .ZN(O12836));
  INVX1 G35737 (.I(W24781), .ZN(W41329));
  INVX1 G35738 (.I(W6436), .ZN(W9588));
  INVX1 G35739 (.I(W39491), .ZN(O12872));
  INVX1 G35740 (.I(I741), .ZN(W7760));
  INVX1 G35741 (.I(I1416), .ZN(W7758));
  INVX1 G35742 (.I(W17884), .ZN(O12876));
  INVX1 G35743 (.I(W18289), .ZN(O11527));
  INVX1 G35744 (.I(W3420), .ZN(W7757));
  INVX1 G35745 (.I(W6094), .ZN(O11526));
  INVX1 G35746 (.I(W22050), .ZN(W43136));
  INVX1 G35747 (.I(W2377), .ZN(W9589));
  INVX1 G35748 (.I(W7911), .ZN(W9590));
  INVX1 G35749 (.I(W9397), .ZN(W9593));
  INVX1 G35750 (.I(I274), .ZN(W9587));
  INVX1 G35751 (.I(W8503), .ZN(O303));
  INVX1 G35752 (.I(I284), .ZN(W7754));
  INVX1 G35753 (.I(W924), .ZN(W9595));
  INVX1 G35754 (.I(W20938), .ZN(O12878));
  INVX1 G35755 (.I(W36938), .ZN(O11518));
  INVX1 G35756 (.I(I1739), .ZN(W9597));
  INVX1 G35757 (.I(W3556), .ZN(W7750));
  INVX1 G35758 (.I(W4118), .ZN(W9598));
  INVX1 G35759 (.I(W10942), .ZN(O11514));
  INVX1 G35760 (.I(W6030), .ZN(W7744));
  INVX1 G35761 (.I(W1197), .ZN(W7741));
  INVX1 G35762 (.I(W19804), .ZN(W43120));
  INVX1 G35763 (.I(W16140), .ZN(W43110));
  INVX1 G35764 (.I(W7551), .ZN(O12860));
  INVX1 G35765 (.I(W31076), .ZN(O11539));
  INVX1 G35766 (.I(W31751), .ZN(W41350));
  INVX1 G35767 (.I(W14973), .ZN(W41349));
  INVX1 G35768 (.I(W30859), .ZN(W43113));
  INVX1 G35769 (.I(I1494), .ZN(W9574));
  INVX1 G35770 (.I(W22691), .ZN(O12863));
  INVX1 G35771 (.I(I694), .ZN(W7772));
  INVX1 G35772 (.I(W8575), .ZN(W43117));
  INVX1 G35773 (.I(W6482), .ZN(W7771));
  INVX1 G35774 (.I(W613), .ZN(W7768));
  INVX1 G35775 (.I(W4934), .ZN(W9533));
  INVX1 G35776 (.I(W144), .ZN(W7766));
  INVX1 G35777 (.I(W9548), .ZN(W9577));
  INVX1 G35778 (.I(I631), .ZN(W9578));
  INVX1 G35779 (.I(W29743), .ZN(W41343));
  INVX1 G35780 (.I(I272), .ZN(W9580));
  INVX1 G35781 (.I(W5328), .ZN(O12867));
  INVX1 G35782 (.I(W16710), .ZN(O11532));
  INVX1 G35783 (.I(W9488), .ZN(W9583));
  INVX1 G35784 (.I(W2877), .ZN(W7762));
  INVX1 G35785 (.I(W34794), .ZN(O12871));
  INVX1 G35786 (.I(W35838), .ZN(W43128));
  INVX1 G35787 (.I(W18429), .ZN(O11610));
  INVX1 G35788 (.I(W3594), .ZN(W9475));
  INVX1 G35789 (.I(W40333), .ZN(O12768));
  INVX1 G35790 (.I(W34865), .ZN(W41452));
  INVX1 G35791 (.I(W21159), .ZN(O11614));
  INVX1 G35792 (.I(W16218), .ZN(W42999));
  INVX1 G35793 (.I(W40222), .ZN(W41450));
  INVX1 G35794 (.I(W1747), .ZN(W7890));
  INVX1 G35795 (.I(I1945), .ZN(W7887));
  INVX1 G35796 (.I(W25842), .ZN(W43004));
  INVX1 G35797 (.I(W7165), .ZN(O11612));
  INVX1 G35798 (.I(W29469), .ZN(O11611));
  INVX1 G35799 (.I(W9651), .ZN(W41446));
  INVX1 G35800 (.I(W33761), .ZN(W41456));
  INVX1 G35801 (.I(W19655), .ZN(O11606));
  INVX1 G35802 (.I(I239), .ZN(W9487));
  INVX1 G35803 (.I(W6524), .ZN(W7874));
  INVX1 G35804 (.I(W6719), .ZN(W9491));
  INVX1 G35805 (.I(W22494), .ZN(W43012));
  INVX1 G35806 (.I(W2107), .ZN(W7872));
  INVX1 G35807 (.I(W8720), .ZN(W9492));
  INVX1 G35808 (.I(I1012), .ZN(W9493));
  INVX1 G35809 (.I(W1702), .ZN(W7871));
  INVX1 G35810 (.I(W5117), .ZN(W7869));
  INVX1 G35811 (.I(W665), .ZN(W7867));
  INVX1 G35812 (.I(W38265), .ZN(O12763));
  INVX1 G35813 (.I(W9400), .ZN(W9461));
  INVX1 G35814 (.I(W35925), .ZN(O12755));
  INVX1 G35815 (.I(I1473), .ZN(W7916));
  INVX1 G35816 (.I(W6473), .ZN(W9462));
  INVX1 G35817 (.I(W679), .ZN(O11625));
  INVX1 G35818 (.I(W7026), .ZN(W7912));
  INVX1 G35819 (.I(W19943), .ZN(O11624));
  INVX1 G35820 (.I(W2689), .ZN(W7908));
  INVX1 G35821 (.I(W3358), .ZN(W7907));
  INVX1 G35822 (.I(W16098), .ZN(O12762));
  INVX1 G35823 (.I(W7629), .ZN(W9470));
  INVX1 G35824 (.I(W25915), .ZN(W41465));
  INVX1 G35825 (.I(W16403), .ZN(O11598));
  INVX1 G35826 (.I(W2172), .ZN(O11621));
  INVX1 G35827 (.I(I918), .ZN(W7906));
  INVX1 G35828 (.I(W2354), .ZN(W9472));
  INVX1 G35829 (.I(W6639), .ZN(O11619));
  INVX1 G35830 (.I(I863), .ZN(W7905));
  INVX1 G35831 (.I(I1156), .ZN(W7903));
  INVX1 G35832 (.I(W5908), .ZN(W42993));
  INVX1 G35833 (.I(W2573), .ZN(W7900));
  INVX1 G35834 (.I(W11169), .ZN(O11618));
  INVX1 G35835 (.I(I1884), .ZN(W9474));
  INVX1 G35836 (.I(W14571), .ZN(O11616));
  INVX1 G35837 (.I(I1669), .ZN(W9519));
  INVX1 G35838 (.I(W8341), .ZN(W9513));
  INVX1 G35839 (.I(W14630), .ZN(O11580));
  INVX1 G35840 (.I(W4313), .ZN(W7843));
  INVX1 G35841 (.I(W1228), .ZN(W7842));
  INVX1 G35842 (.I(W5640), .ZN(W7841));
  INVX1 G35843 (.I(W4607), .ZN(W7839));
  INVX1 G35844 (.I(W2449), .ZN(O12809));
  INVX1 G35845 (.I(W175), .ZN(O11578));
  INVX1 G35846 (.I(W3442), .ZN(W7838));
  INVX1 G35847 (.I(W10952), .ZN(O12812));
  INVX1 G35848 (.I(W38996), .ZN(O11575));
  INVX1 G35849 (.I(W9241), .ZN(O11574));
  INVX1 G35850 (.I(I1390), .ZN(W7844));
  INVX1 G35851 (.I(W17568), .ZN(W41401));
  INVX1 G35852 (.I(W3841), .ZN(W9522));
  INVX1 G35853 (.I(W5865), .ZN(O11571));
  INVX1 G35854 (.I(W6216), .ZN(W7833));
  INVX1 G35855 (.I(I414), .ZN(W7832));
  INVX1 G35856 (.I(W7623), .ZN(W9526));
  INVX1 G35857 (.I(W5905), .ZN(W9527));
  INVX1 G35858 (.I(I1750), .ZN(W7830));
  INVX1 G35859 (.I(W1464), .ZN(O297));
  INVX1 G35860 (.I(W10926), .ZN(O12816));
  INVX1 G35861 (.I(W24450), .ZN(W41392));
  INVX1 G35862 (.I(W5832), .ZN(W9503));
  INVX1 G35863 (.I(W2888), .ZN(W7866));
  INVX1 G35864 (.I(W6027), .ZN(W7862));
  INVX1 G35865 (.I(W20302), .ZN(O11596));
  INVX1 G35866 (.I(W5406), .ZN(W7859));
  INVX1 G35867 (.I(W6617), .ZN(W9496));
  INVX1 G35868 (.I(I1725), .ZN(O204));
  INVX1 G35869 (.I(I1160), .ZN(W7854));
  INVX1 G35870 (.I(W13729), .ZN(O12791));
  INVX1 G35871 (.I(W6375), .ZN(W7853));
  INVX1 G35872 (.I(W10714), .ZN(O12793));
  INVX1 G35873 (.I(W16054), .ZN(O11591));
  INVX1 G35874 (.I(W4445), .ZN(O12795));
  INVX1 G35875 (.I(W4658), .ZN(W9823));
  INVX1 G35876 (.I(W27605), .ZN(W41422));
  INVX1 G35877 (.I(W8595), .ZN(W9505));
  INVX1 G35878 (.I(W543), .ZN(O296));
  INVX1 G35879 (.I(W28872), .ZN(W43033));
  INVX1 G35880 (.I(W2332), .ZN(W7847));
  INVX1 G35881 (.I(W16594), .ZN(O12799));
  INVX1 G35882 (.I(W12254), .ZN(O12800));
  INVX1 G35883 (.I(W17179), .ZN(O12801));
  INVX1 G35884 (.I(W5611), .ZN(W9510));
  INVX1 G35885 (.I(W20848), .ZN(O12802));
  INVX1 G35886 (.I(W24578), .ZN(O11582));
  INVX1 G35887 (.I(W33494), .ZN(O17498));
  INVX1 G35888 (.I(I1710), .ZN(W2349));
  INVX1 G35889 (.I(W346), .ZN(W2350));
  INVX1 G35890 (.I(I1976), .ZN(W2351));
  INVX1 G35891 (.I(W2072), .ZN(W2353));
  INVX1 G35892 (.I(W29296), .ZN(O17503));
  INVX1 G35893 (.I(W19029), .ZN(O17502));
  INVX1 G35894 (.I(W7657), .ZN(O17501));
  INVX1 G35895 (.I(I504), .ZN(W2355));
  INVX1 G35896 (.I(I1092), .ZN(W2356));
  INVX1 G35897 (.I(W18548), .ZN(O17511));
  INVX1 G35898 (.I(W709), .ZN(W2361));
  INVX1 G35899 (.I(W835), .ZN(W2363));
  INVX1 G35900 (.I(I148), .ZN(O17492));
  INVX1 G35901 (.I(I1259), .ZN(W2364));
  INVX1 G35902 (.I(W20532), .ZN(O17490));
  INVX1 G35903 (.I(I1881), .ZN(W2365));
  INVX1 G35904 (.I(W16285), .ZN(O17486));
  INVX1 G35905 (.I(I1355), .ZN(W2369));
  INVX1 G35906 (.I(W15887), .ZN(O17524));
  INVX1 G35907 (.I(W48087), .ZN(O17531));
  INVX1 G35908 (.I(W1519), .ZN(W2329));
  INVX1 G35909 (.I(W1615), .ZN(W2330));
  INVX1 G35910 (.I(W10431), .ZN(W48663));
  INVX1 G35911 (.I(W1683), .ZN(W2331));
  INVX1 G35912 (.I(I910), .ZN(W2333));
  INVX1 G35913 (.I(I1881), .ZN(W2334));
  INVX1 G35914 (.I(I1542), .ZN(O17526));
  INVX1 G35915 (.I(I474), .ZN(W2335));
  INVX1 G35916 (.I(W1416), .ZN(W2376));
  INVX1 G35917 (.I(W1475), .ZN(W2336));
  INVX1 G35918 (.I(W904), .ZN(W2337));
  INVX1 G35919 (.I(I923), .ZN(W2341));
  INVX1 G35920 (.I(W40225), .ZN(O17517));
  INVX1 G35921 (.I(W8041), .ZN(O17516));
  INVX1 G35922 (.I(W47090), .ZN(O17515));
  INVX1 G35923 (.I(W27772), .ZN(O17513));
  INVX1 G35924 (.I(W44293), .ZN(O17512));
  INVX1 G35925 (.I(W33565), .ZN(O17447));
  INVX1 G35926 (.I(W2308), .ZN(W2391));
  INVX1 G35927 (.I(W31885), .ZN(O17458));
  INVX1 G35928 (.I(W20023), .ZN(O17457));
  INVX1 G35929 (.I(I874), .ZN(W2392));
  INVX1 G35930 (.I(W17165), .ZN(O17455));
  INVX1 G35931 (.I(W43344), .ZN(O17454));
  INVX1 G35932 (.I(I824), .ZN(W2393));
  INVX1 G35933 (.I(W1193), .ZN(W2396));
  INVX1 G35934 (.I(W19304), .ZN(O17448));
  INVX1 G35935 (.I(W40216), .ZN(O17460));
  INVX1 G35936 (.I(W32343), .ZN(O17446));
  INVX1 G35937 (.I(W25689), .ZN(O17444));
  INVX1 G35938 (.I(W2234), .ZN(W2403));
  INVX1 G35939 (.I(W2357), .ZN(W2405));
  INVX1 G35940 (.I(W15446), .ZN(W48569));
  INVX1 G35941 (.I(W114), .ZN(W2407));
  INVX1 G35942 (.I(I1337), .ZN(W2411));
  INVX1 G35943 (.I(I1145), .ZN(W2412));
  INVX1 G35944 (.I(W7714), .ZN(W48600));
  INVX1 G35945 (.I(W45426), .ZN(O17481));
  INVX1 G35946 (.I(I217), .ZN(O17480));
  INVX1 G35947 (.I(W43075), .ZN(O17478));
  INVX1 G35948 (.I(W35956), .ZN(O17477));
  INVX1 G35949 (.I(W185), .ZN(W2380));
  INVX1 G35950 (.I(W698), .ZN(W2382));
  INVX1 G35951 (.I(W36726), .ZN(O17473));
  INVX1 G35952 (.I(W46732), .ZN(O17472));
  INVX1 G35953 (.I(W19135), .ZN(O17471));
  INVX1 G35954 (.I(W46030), .ZN(O17532));
  INVX1 G35955 (.I(W468), .ZN(W2384));
  INVX1 G35956 (.I(W33256), .ZN(O17468));
  INVX1 G35957 (.I(W33238), .ZN(O17466));
  INVX1 G35958 (.I(I1044), .ZN(W2387));
  INVX1 G35959 (.I(I1463), .ZN(W2389));
  INVX1 G35960 (.I(W21310), .ZN(O17463));
  INVX1 G35961 (.I(W18050), .ZN(O17462));
  INVX1 G35962 (.I(W11176), .ZN(O17461));
  INVX1 G35963 (.I(W375), .ZN(W2253));
  INVX1 G35964 (.I(W2156), .ZN(W2229));
  INVX1 G35965 (.I(W1973), .ZN(W2230));
  INVX1 G35966 (.I(W1482), .ZN(W2233));
  INVX1 G35967 (.I(W1639), .ZN(W2237));
  INVX1 G35968 (.I(W31124), .ZN(O17612));
  INVX1 G35969 (.I(W3949), .ZN(O17610));
  INVX1 G35970 (.I(W727), .ZN(W2243));
  INVX1 G35971 (.I(W25386), .ZN(O17605));
  INVX1 G35972 (.I(W1502), .ZN(W2252));
  INVX1 G35973 (.I(W16183), .ZN(O17619));
  INVX1 G35974 (.I(W886), .ZN(W2255));
  INVX1 G35975 (.I(W26269), .ZN(O17599));
  INVX1 G35976 (.I(W8935), .ZN(O17597));
  INVX1 G35977 (.I(W2173), .ZN(W2260));
  INVX1 G35978 (.I(W45068), .ZN(O17594));
  INVX1 G35979 (.I(I250), .ZN(O17591));
  INVX1 G35980 (.I(W10519), .ZN(O17590));
  INVX1 G35981 (.I(I1887), .ZN(W2267));
  INVX1 G35982 (.I(W1291), .ZN(W2219));
  INVX1 G35983 (.I(W16960), .ZN(O17644));
  INVX1 G35984 (.I(I1000), .ZN(W2200));
  INVX1 G35985 (.I(W25523), .ZN(O17642));
  INVX1 G35986 (.I(I1815), .ZN(W2202));
  INVX1 G35987 (.I(W79), .ZN(O17641));
  INVX1 G35988 (.I(W196), .ZN(W2205));
  INVX1 G35989 (.I(I1374), .ZN(W2206));
  INVX1 G35990 (.I(I303), .ZN(W2207));
  INVX1 G35991 (.I(I1507), .ZN(W2217));
  INVX1 G35992 (.I(W27722), .ZN(O17586));
  INVX1 G35993 (.I(W2141), .ZN(W2220));
  INVX1 G35994 (.I(W5273), .ZN(O17628));
  INVX1 G35995 (.I(I1069), .ZN(W2224));
  INVX1 G35996 (.I(W34952), .ZN(O17625));
  INVX1 G35997 (.I(W37190), .ZN(O17624));
  INVX1 G35998 (.I(W10988), .ZN(O17622));
  INVX1 G35999 (.I(W25447), .ZN(O17621));
  INVX1 G36000 (.I(W1640), .ZN(O17620));
  INVX1 G36001 (.I(I1599), .ZN(W2314));
  INVX1 G36002 (.I(W16630), .ZN(O17562));
  INVX1 G36003 (.I(W10904), .ZN(O17560));
  INVX1 G36004 (.I(W4165), .ZN(O17559));
  INVX1 G36005 (.I(W1814), .ZN(W2301));
  INVX1 G36006 (.I(W977), .ZN(W2304));
  INVX1 G36007 (.I(W14648), .ZN(O17552));
  INVX1 G36008 (.I(I1254), .ZN(W2309));
  INVX1 G36009 (.I(W1231), .ZN(W2311));
  INVX1 G36010 (.I(W1350), .ZN(W2313));
  INVX1 G36011 (.I(W3576), .ZN(O17563));
  INVX1 G36012 (.I(W3995), .ZN(O17546));
  INVX1 G36013 (.I(W4266), .ZN(O17544));
  INVX1 G36014 (.I(W26690), .ZN(O17539));
  INVX1 G36015 (.I(I1875), .ZN(W2322));
  INVX1 G36016 (.I(I1736), .ZN(O17536));
  INVX1 G36017 (.I(I1498), .ZN(W2324));
  INVX1 G36018 (.I(W14548), .ZN(O17534));
  INVX1 G36019 (.I(W540), .ZN(W2326));
  INVX1 G36020 (.I(W918), .ZN(W2281));
  INVX1 G36021 (.I(W31957), .ZN(W48727));
  INVX1 G36022 (.I(I1048), .ZN(W2270));
  INVX1 G36023 (.I(W160), .ZN(W2271));
  INVX1 G36024 (.I(W1968), .ZN(W2275));
  INVX1 G36025 (.I(W1898), .ZN(W2277));
  INVX1 G36026 (.I(W38092), .ZN(O17578));
  INVX1 G36027 (.I(W34784), .ZN(O17577));
  INVX1 G36028 (.I(W3173), .ZN(O17576));
  INVX1 G36029 (.I(W21386), .ZN(O17438));
  INVX1 G36030 (.I(I85), .ZN(W2285));
  INVX1 G36031 (.I(W1153), .ZN(W2286));
  INVX1 G36032 (.I(W46817), .ZN(O17569));
  INVX1 G36033 (.I(W1902), .ZN(W2291));
  INVX1 G36034 (.I(I814), .ZN(W2296));
  INVX1 G36035 (.I(W44947), .ZN(W48705));
  INVX1 G36036 (.I(W33319), .ZN(O17566));
  INVX1 G36037 (.I(W27878), .ZN(O17565));
  INVX1 G36038 (.I(W17311), .ZN(O17291));
  INVX1 G36039 (.I(W4245), .ZN(O17303));
  INVX1 G36040 (.I(W17455), .ZN(O17302));
  INVX1 G36041 (.I(W2129), .ZN(W2559));
  INVX1 G36042 (.I(W1929), .ZN(W2560));
  INVX1 G36043 (.I(I422), .ZN(W2564));
  INVX1 G36044 (.I(W1808), .ZN(W2565));
  INVX1 G36045 (.I(W9646), .ZN(O17295));
  INVX1 G36046 (.I(W308), .ZN(W2566));
  INVX1 G36047 (.I(W695), .ZN(W2567));
  INVX1 G36048 (.I(W41800), .ZN(O17304));
  INVX1 G36049 (.I(W13104), .ZN(O17290));
  INVX1 G36050 (.I(W42203), .ZN(O17289));
  INVX1 G36051 (.I(W864), .ZN(W2577));
  INVX1 G36052 (.I(I776), .ZN(W2578));
  INVX1 G36053 (.I(I948), .ZN(W2579));
  INVX1 G36054 (.I(W37056), .ZN(W48389));
  INVX1 G36055 (.I(W1149), .ZN(W2580));
  INVX1 G36056 (.I(I1193), .ZN(W2582));
  INVX1 G36057 (.I(W10960), .ZN(O17318));
  INVX1 G36058 (.I(W43420), .ZN(O17330));
  INVX1 G36059 (.I(W2325), .ZN(O22));
  INVX1 G36060 (.I(W33069), .ZN(W48437));
  INVX1 G36061 (.I(W18795), .ZN(O17326));
  INVX1 G36062 (.I(W4074), .ZN(O17325));
  INVX1 G36063 (.I(W20528), .ZN(O17323));
  INVX1 G36064 (.I(W765), .ZN(W2539));
  INVX1 G36065 (.I(W26416), .ZN(O17321));
  INVX1 G36066 (.I(I1174), .ZN(W2540));
  INVX1 G36067 (.I(W599), .ZN(W2583));
  INVX1 G36068 (.I(W719), .ZN(W2544));
  INVX1 G36069 (.I(I1843), .ZN(W2545));
  INVX1 G36070 (.I(W144), .ZN(W2548));
  INVX1 G36071 (.I(W45049), .ZN(O17312));
  INVX1 G36072 (.I(W20165), .ZN(O17308));
  INVX1 G36073 (.I(W1662), .ZN(W2558));
  INVX1 G36074 (.I(W19723), .ZN(O17306));
  INVX1 G36075 (.I(W21762), .ZN(O17305));
  INVX1 G36076 (.I(I331), .ZN(W2635));
  INVX1 G36077 (.I(W8232), .ZN(O17248));
  INVX1 G36078 (.I(W21092), .ZN(O17247));
  INVX1 G36079 (.I(W35248), .ZN(O17242));
  INVX1 G36080 (.I(W15358), .ZN(O17240));
  INVX1 G36081 (.I(W1729), .ZN(O24));
  INVX1 G36082 (.I(I410), .ZN(W2633));
  INVX1 G36083 (.I(W28239), .ZN(O17236));
  INVX1 G36084 (.I(W9778), .ZN(O17235));
  INVX1 G36085 (.I(W1600), .ZN(W2634));
  INVX1 G36086 (.I(W676), .ZN(W2620));
  INVX1 G36087 (.I(I414), .ZN(W2638));
  INVX1 G36088 (.I(W1950), .ZN(W2641));
  INVX1 G36089 (.I(W22700), .ZN(O17226));
  INVX1 G36090 (.I(I1724), .ZN(W2648));
  INVX1 G36091 (.I(W41607), .ZN(O17223));
  INVX1 G36092 (.I(W11006), .ZN(O17221));
  INVX1 G36093 (.I(W2151), .ZN(W2653));
  INVX1 G36094 (.I(W10369), .ZN(O17218));
  INVX1 G36095 (.I(I634), .ZN(W2596));
  INVX1 G36096 (.I(W1505), .ZN(W2585));
  INVX1 G36097 (.I(W2038), .ZN(W2587));
  INVX1 G36098 (.I(I123), .ZN(O23));
  INVX1 G36099 (.I(I829), .ZN(W2589));
  INVX1 G36100 (.I(W23918), .ZN(O17272));
  INVX1 G36101 (.I(W35041), .ZN(O17271));
  INVX1 G36102 (.I(W1238), .ZN(W2593));
  INVX1 G36103 (.I(I410), .ZN(W2595));
  INVX1 G36104 (.I(W46914), .ZN(O17331));
  INVX1 G36105 (.I(I1341), .ZN(W2601));
  INVX1 G36106 (.I(W134), .ZN(W2606));
  INVX1 G36107 (.I(W1324), .ZN(W2611));
  INVX1 G36108 (.I(W317), .ZN(W2612));
  INVX1 G36109 (.I(W37338), .ZN(O17256));
  INVX1 G36110 (.I(W1673), .ZN(W2615));
  INVX1 G36111 (.I(W1610), .ZN(W2617));
  INVX1 G36112 (.I(W18737), .ZN(O17251));
  INVX1 G36113 (.I(W16174), .ZN(O17411));
  INVX1 G36114 (.I(W4382), .ZN(W48541));
  INVX1 G36115 (.I(W993), .ZN(W2444));
  INVX1 G36116 (.I(W2350), .ZN(W48535));
  INVX1 G36117 (.I(W2410), .ZN(W2446));
  INVX1 G36118 (.I(W4829), .ZN(O17418));
  INVX1 G36119 (.I(W16982), .ZN(O17417));
  INVX1 G36120 (.I(W16031), .ZN(O17416));
  INVX1 G36121 (.I(W18745), .ZN(O17414));
  INVX1 G36122 (.I(I1189), .ZN(W2450));
  INVX1 G36123 (.I(W1919), .ZN(W2432));
  INVX1 G36124 (.I(W23836), .ZN(O17410));
  INVX1 G36125 (.I(W11), .ZN(W2451));
  INVX1 G36126 (.I(W22365), .ZN(W48523));
  INVX1 G36127 (.I(W34128), .ZN(O17408));
  INVX1 G36128 (.I(W229), .ZN(W2452));
  INVX1 G36129 (.I(W33613), .ZN(O17406));
  INVX1 G36130 (.I(W20815), .ZN(O17404));
  INVX1 G36131 (.I(I625), .ZN(W2454));
  INVX1 G36132 (.I(W17725), .ZN(O17431));
  INVX1 G36133 (.I(W1134), .ZN(W2418));
  INVX1 G36134 (.I(I1308), .ZN(W2419));
  INVX1 G36135 (.I(W25158), .ZN(O17435));
  INVX1 G36136 (.I(W1011), .ZN(W2420));
  INVX1 G36137 (.I(W30943), .ZN(W48558));
  INVX1 G36138 (.I(W19101), .ZN(W48556));
  INVX1 G36139 (.I(W1500), .ZN(W48554));
  INVX1 G36140 (.I(W652), .ZN(W2424));
  INVX1 G36141 (.I(I135), .ZN(W2427));
  INVX1 G36142 (.I(W905), .ZN(W2455));
  INVX1 G36143 (.I(I1873), .ZN(W2428));
  INVX1 G36144 (.I(W17026), .ZN(O17429));
  INVX1 G36145 (.I(I635), .ZN(W2429));
  INVX1 G36146 (.I(W26473), .ZN(O17427));
  INVX1 G36147 (.I(W15353), .ZN(O17426));
  INVX1 G36148 (.I(W43862), .ZN(W48545));
  INVX1 G36149 (.I(I1142), .ZN(W2430));
  INVX1 G36150 (.I(I766), .ZN(W2431));
  INVX1 G36151 (.I(W2238), .ZN(W2519));
  INVX1 G36152 (.I(W26082), .ZN(O17364));
  INVX1 G36153 (.I(W36326), .ZN(O17359));
  INVX1 G36154 (.I(W26), .ZN(O17358));
  INVX1 G36155 (.I(I745), .ZN(O21));
  INVX1 G36156 (.I(I409), .ZN(W2512));
  INVX1 G36157 (.I(W2140), .ZN(W2513));
  INVX1 G36158 (.I(W16701), .ZN(O17348));
  INVX1 G36159 (.I(W1643), .ZN(W2518));
  INVX1 G36160 (.I(W1082), .ZN(O17347));
  INVX1 G36161 (.I(W32863), .ZN(W48478));
  INVX1 G36162 (.I(I1963), .ZN(W2520));
  INVX1 G36163 (.I(W18097), .ZN(O17344));
  INVX1 G36164 (.I(W1468), .ZN(W2525));
  INVX1 G36165 (.I(W70), .ZN(W2528));
  INVX1 G36166 (.I(W9141), .ZN(O17338));
  INVX1 G36167 (.I(W45923), .ZN(O17335));
  INVX1 G36168 (.I(W653), .ZN(W2534));
  INVX1 G36169 (.I(W1968), .ZN(O17332));
  INVX1 G36170 (.I(W2431), .ZN(O20));
  INVX1 G36171 (.I(W1277), .ZN(W2456));
  INVX1 G36172 (.I(W1201), .ZN(W2462));
  INVX1 G36173 (.I(W42790), .ZN(O17396));
  INVX1 G36174 (.I(W875), .ZN(O19));
  INVX1 G36175 (.I(I1800), .ZN(W2465));
  INVX1 G36176 (.I(W36541), .ZN(O17391));
  INVX1 G36177 (.I(W33779), .ZN(O17388));
  INVX1 G36178 (.I(W423), .ZN(W2473));
  INVX1 G36179 (.I(W18856), .ZN(O17646));
  INVX1 G36180 (.I(W33137), .ZN(O17384));
  INVX1 G36181 (.I(W998), .ZN(W2479));
  INVX1 G36182 (.I(W21323), .ZN(O17380));
  INVX1 G36183 (.I(W569), .ZN(W2482));
  INVX1 G36184 (.I(W23330), .ZN(O17375));
  INVX1 G36185 (.I(W2466), .ZN(W2485));
  INVX1 G36186 (.I(I1312), .ZN(W2493));
  INVX1 G36187 (.I(W1948), .ZN(W2496));
  INVX1 G36188 (.I(W46078), .ZN(W49078));
  INVX1 G36189 (.I(W1348), .ZN(W1902));
  INVX1 G36190 (.I(W23248), .ZN(O17918));
  INVX1 G36191 (.I(I1394), .ZN(O17917));
  INVX1 G36192 (.I(W17659), .ZN(O17916));
  INVX1 G36193 (.I(W1258), .ZN(W1905));
  INVX1 G36194 (.I(W204), .ZN(W1907));
  INVX1 G36195 (.I(W39786), .ZN(O17914));
  INVX1 G36196 (.I(I1355), .ZN(W1912));
  INVX1 G36197 (.I(W11696), .ZN(O17908));
  INVX1 G36198 (.I(I5), .ZN(W1898));
  INVX1 G36199 (.I(I590), .ZN(W1915));
  INVX1 G36200 (.I(W1326), .ZN(W1927));
  INVX1 G36201 (.I(W19077), .ZN(O17899));
  INVX1 G36202 (.I(W17636), .ZN(O17898));
  INVX1 G36203 (.I(W24183), .ZN(O17896));
  INVX1 G36204 (.I(I1580), .ZN(W1931));
  INVX1 G36205 (.I(I616), .ZN(W1933));
  INVX1 G36206 (.I(W635), .ZN(W1934));
  INVX1 G36207 (.I(W12197), .ZN(O17936));
  INVX1 G36208 (.I(W896), .ZN(W1865));
  INVX1 G36209 (.I(W40970), .ZN(O17949));
  INVX1 G36210 (.I(W30361), .ZN(O17948));
  INVX1 G36211 (.I(W555), .ZN(W1867));
  INVX1 G36212 (.I(W960), .ZN(W1870));
  INVX1 G36213 (.I(W5009), .ZN(O17943));
  INVX1 G36214 (.I(W24483), .ZN(O17942));
  INVX1 G36215 (.I(W29837), .ZN(O17941));
  INVX1 G36216 (.I(I1029), .ZN(W1874));
  INVX1 G36217 (.I(I1556), .ZN(W1937));
  INVX1 G36218 (.I(W44467), .ZN(O17935));
  INVX1 G36219 (.I(I1598), .ZN(W1883));
  INVX1 G36220 (.I(W1812), .ZN(W1885));
  INVX1 G36221 (.I(W33292), .ZN(O17929));
  INVX1 G36222 (.I(I1074), .ZN(W1890));
  INVX1 G36223 (.I(W588), .ZN(W1891));
  INVX1 G36224 (.I(W1115), .ZN(W1893));
  INVX1 G36225 (.I(W46617), .ZN(O17924));
  INVX1 G36226 (.I(W38084), .ZN(O17857));
  INVX1 G36227 (.I(W1364), .ZN(W1959));
  INVX1 G36228 (.I(W1162), .ZN(W1962));
  INVX1 G36229 (.I(W41192), .ZN(O17866));
  INVX1 G36230 (.I(W1956), .ZN(W1963));
  INVX1 G36231 (.I(W47067), .ZN(O17864));
  INVX1 G36232 (.I(W356), .ZN(W1965));
  INVX1 G36233 (.I(W615), .ZN(O17861));
  INVX1 G36234 (.I(W863), .ZN(W1968));
  INVX1 G36235 (.I(W289), .ZN(W1970));
  INVX1 G36236 (.I(W13046), .ZN(O17869));
  INVX1 G36237 (.I(W28161), .ZN(O17856));
  INVX1 G36238 (.I(W45265), .ZN(O17854));
  INVX1 G36239 (.I(W44386), .ZN(W49018));
  INVX1 G36240 (.I(W26108), .ZN(O17852));
  INVX1 G36241 (.I(W1963), .ZN(W1980));
  INVX1 G36242 (.I(W15903), .ZN(O17849));
  INVX1 G36243 (.I(W31541), .ZN(O17848));
  INVX1 G36244 (.I(W23132), .ZN(O17847));
  INVX1 G36245 (.I(W247), .ZN(W1947));
  INVX1 G36246 (.I(I495), .ZN(W1938));
  INVX1 G36247 (.I(W64), .ZN(W1939));
  INVX1 G36248 (.I(W1352), .ZN(W1940));
  INVX1 G36249 (.I(W1792), .ZN(W1942));
  INVX1 G36250 (.I(W11816), .ZN(O17885));
  INVX1 G36251 (.I(W1727), .ZN(W1946));
  INVX1 G36252 (.I(W16090), .ZN(O17883));
  INVX1 G36253 (.I(W44998), .ZN(O17882));
  INVX1 G36254 (.I(W306), .ZN(W1862));
  INVX1 G36255 (.I(W15302), .ZN(O17879));
  INVX1 G36256 (.I(W20464), .ZN(O17878));
  INVX1 G36257 (.I(W35879), .ZN(O17876));
  INVX1 G36258 (.I(I1431), .ZN(W1950));
  INVX1 G36259 (.I(W1224), .ZN(W1952));
  INVX1 G36260 (.I(W312), .ZN(W1955));
  INVX1 G36261 (.I(W47501), .ZN(O17870));
  INVX1 G36262 (.I(W45902), .ZN(W49037));
  INVX1 G36263 (.I(I452), .ZN(W1799));
  INVX1 G36264 (.I(W46858), .ZN(O18024));
  INVX1 G36265 (.I(W795), .ZN(W1792));
  INVX1 G36266 (.I(I1212), .ZN(W1793));
  INVX1 G36267 (.I(W32883), .ZN(O18020));
  INVX1 G36268 (.I(I1979), .ZN(W1796));
  INVX1 G36269 (.I(I976), .ZN(W1797));
  INVX1 G36270 (.I(W22288), .ZN(O18018));
  INVX1 G36271 (.I(W4633), .ZN(O18017));
  INVX1 G36272 (.I(W1759), .ZN(W1798));
  INVX1 G36273 (.I(W302), .ZN(W1791));
  INVX1 G36274 (.I(W642), .ZN(W1801));
  INVX1 G36275 (.I(W9226), .ZN(O18013));
  INVX1 G36276 (.I(W33903), .ZN(O18012));
  INVX1 G36277 (.I(W44686), .ZN(O18011));
  INVX1 G36278 (.I(W10220), .ZN(O18009));
  INVX1 G36279 (.I(W25086), .ZN(O18008));
  INVX1 G36280 (.I(W24311), .ZN(O18007));
  INVX1 G36281 (.I(W2634), .ZN(O18006));
  INVX1 G36282 (.I(W759), .ZN(W1783));
  INVX1 G36283 (.I(W13759), .ZN(O18046));
  INVX1 G36284 (.I(I60), .ZN(W1773));
  INVX1 G36285 (.I(W34859), .ZN(O18044));
  INVX1 G36286 (.I(W27907), .ZN(O18043));
  INVX1 G36287 (.I(W29458), .ZN(O18041));
  INVX1 G36288 (.I(W43262), .ZN(O18040));
  INVX1 G36289 (.I(W2353), .ZN(W49220));
  INVX1 G36290 (.I(W440), .ZN(W1780));
  INVX1 G36291 (.I(I1110), .ZN(W1781));
  INVX1 G36292 (.I(W20432), .ZN(O18005));
  INVX1 G36293 (.I(W14805), .ZN(O18033));
  INVX1 G36294 (.I(W19309), .ZN(O18031));
  INVX1 G36295 (.I(I1758), .ZN(W1786));
  INVX1 G36296 (.I(W5635), .ZN(O18029));
  INVX1 G36297 (.I(W1570), .ZN(W1788));
  INVX1 G36298 (.I(W31221), .ZN(O18028));
  INVX1 G36299 (.I(W1396), .ZN(W1789));
  INVX1 G36300 (.I(W1346), .ZN(W1790));
  INVX1 G36301 (.I(W10773), .ZN(O17965));
  INVX1 G36302 (.I(W15686), .ZN(O17981));
  INVX1 G36303 (.I(W10337), .ZN(O17980));
  INVX1 G36304 (.I(W1059), .ZN(W1835));
  INVX1 G36305 (.I(W18203), .ZN(O17977));
  INVX1 G36306 (.I(W32670), .ZN(O17976));
  INVX1 G36307 (.I(W31687), .ZN(O17974));
  INVX1 G36308 (.I(W1061), .ZN(W1839));
  INVX1 G36309 (.I(W48165), .ZN(O17971));
  INVX1 G36310 (.I(W1437), .ZN(O17968));
  INVX1 G36311 (.I(W21935), .ZN(O17982));
  INVX1 G36312 (.I(W1241), .ZN(W1847));
  INVX1 G36313 (.I(I1690), .ZN(W1853));
  INVX1 G36314 (.I(W44814), .ZN(O17961));
  INVX1 G36315 (.I(W24611), .ZN(O17960));
  INVX1 G36316 (.I(W7943), .ZN(W49133));
  INVX1 G36317 (.I(W317), .ZN(W1856));
  INVX1 G36318 (.I(W7896), .ZN(O17956));
  INVX1 G36319 (.I(I1667), .ZN(W1860));
  INVX1 G36320 (.I(I1808), .ZN(W1820));
  INVX1 G36321 (.I(W30135), .ZN(O18004));
  INVX1 G36322 (.I(I49), .ZN(W1805));
  INVX1 G36323 (.I(W16056), .ZN(O18002));
  INVX1 G36324 (.I(I996), .ZN(W1812));
  INVX1 G36325 (.I(W1208), .ZN(W1813));
  INVX1 G36326 (.I(W13589), .ZN(O18000));
  INVX1 G36327 (.I(W1778), .ZN(W1814));
  INVX1 G36328 (.I(W27793), .ZN(O17998));
  INVX1 G36329 (.I(W25848), .ZN(O17845));
  INVX1 G36330 (.I(W19057), .ZN(O17995));
  INVX1 G36331 (.I(W1230), .ZN(W1825));
  INVX1 G36332 (.I(I1180), .ZN(W1826));
  INVX1 G36333 (.I(W16256), .ZN(O17990));
  INVX1 G36334 (.I(I1116), .ZN(W1827));
  INVX1 G36335 (.I(W20413), .ZN(O17987));
  INVX1 G36336 (.I(W5082), .ZN(O17986));
  INVX1 G36337 (.I(I534), .ZN(W1832));
  INVX1 G36338 (.I(I1439), .ZN(W2153));
  INVX1 G36339 (.I(W591), .ZN(W2134));
  INVX1 G36340 (.I(W1803), .ZN(W2137));
  INVX1 G36341 (.I(I1181), .ZN(W2140));
  INVX1 G36342 (.I(W25955), .ZN(O17708));
  INVX1 G36343 (.I(W1769), .ZN(O17707));
  INVX1 G36344 (.I(W871), .ZN(W2143));
  INVX1 G36345 (.I(I637), .ZN(W2146));
  INVX1 G36346 (.I(W43937), .ZN(O17702));
  INVX1 G36347 (.I(I816), .ZN(W2150));
  INVX1 G36348 (.I(W18897), .ZN(O17714));
  INVX1 G36349 (.I(W12417), .ZN(O17697));
  INVX1 G36350 (.I(W1141), .ZN(W2157));
  INVX1 G36351 (.I(W10159), .ZN(O17694));
  INVX1 G36352 (.I(W2035), .ZN(W2160));
  INVX1 G36353 (.I(W29642), .ZN(O17691));
  INVX1 G36354 (.I(W38022), .ZN(O17690));
  INVX1 G36355 (.I(W27526), .ZN(O17689));
  INVX1 G36356 (.I(W18769), .ZN(O17688));
  INVX1 G36357 (.I(I1442), .ZN(W2118));
  INVX1 G36358 (.I(W6897), .ZN(O17744));
  INVX1 G36359 (.I(I758), .ZN(W2091));
  INVX1 G36360 (.I(W39354), .ZN(O17739));
  INVX1 G36361 (.I(I495), .ZN(W2097));
  INVX1 G36362 (.I(I630), .ZN(W2101));
  INVX1 G36363 (.I(W48535), .ZN(O17734));
  INVX1 G36364 (.I(W1919), .ZN(O17732));
  INVX1 G36365 (.I(W3074), .ZN(O17730));
  INVX1 G36366 (.I(W871), .ZN(W2109));
  INVX1 G36367 (.I(W1781), .ZN(W2165));
  INVX1 G36368 (.I(W1058), .ZN(W2120));
  INVX1 G36369 (.I(W1167), .ZN(W2124));
  INVX1 G36370 (.I(W31877), .ZN(O17722));
  INVX1 G36371 (.I(W12840), .ZN(O17721));
  INVX1 G36372 (.I(W1502), .ZN(W2128));
  INVX1 G36373 (.I(I1036), .ZN(W2129));
  INVX1 G36374 (.I(W31612), .ZN(W48872));
  INVX1 G36375 (.I(W9487), .ZN(O17717));
  INVX1 G36376 (.I(I1646), .ZN(W2190));
  INVX1 G36377 (.I(W45373), .ZN(O17666));
  INVX1 G36378 (.I(W2134), .ZN(W2183));
  INVX1 G36379 (.I(W23778), .ZN(O17662));
  INVX1 G36380 (.I(I1749), .ZN(W2187));
  INVX1 G36381 (.I(W28886), .ZN(O17660));
  INVX1 G36382 (.I(W25431), .ZN(O17659));
  INVX1 G36383 (.I(I467), .ZN(W2188));
  INVX1 G36384 (.I(W38761), .ZN(O17657));
  INVX1 G36385 (.I(W7629), .ZN(O17656));
  INVX1 G36386 (.I(W31023), .ZN(O17667));
  INVX1 G36387 (.I(W1215), .ZN(W2192));
  INVX1 G36388 (.I(W570), .ZN(W2193));
  INVX1 G36389 (.I(I793), .ZN(W2194));
  INVX1 G36390 (.I(W2355), .ZN(O17652));
  INVX1 G36391 (.I(I822), .ZN(W2195));
  INVX1 G36392 (.I(W675), .ZN(W2197));
  INVX1 G36393 (.I(I1289), .ZN(W2198));
  INVX1 G36394 (.I(W33246), .ZN(O17647));
  INVX1 G36395 (.I(W13379), .ZN(W48828));
  INVX1 G36396 (.I(I1820), .ZN(W2167));
  INVX1 G36397 (.I(W26705), .ZN(O17684));
  INVX1 G36398 (.I(W39745), .ZN(O17683));
  INVX1 G36399 (.I(W1438), .ZN(W2170));
  INVX1 G36400 (.I(W36843), .ZN(O17681));
  INVX1 G36401 (.I(W22594), .ZN(O17680));
  INVX1 G36402 (.I(W982), .ZN(W2171));
  INVX1 G36403 (.I(W17370), .ZN(O17678));
  INVX1 G36404 (.I(W45124), .ZN(O17746));
  INVX1 G36405 (.I(W1613), .ZN(W2172));
  INVX1 G36406 (.I(W15643), .ZN(O17676));
  INVX1 G36407 (.I(I1092), .ZN(W2173));
  INVX1 G36408 (.I(W22926), .ZN(O17672));
  INVX1 G36409 (.I(I459), .ZN(W2178));
  INVX1 G36410 (.I(W36402), .ZN(O17669));
  INVX1 G36411 (.I(W9101), .ZN(W48818));
  INVX1 G36412 (.I(I1572), .ZN(W2181));
  INVX1 G36413 (.I(W121), .ZN(W2023));
  INVX1 G36414 (.I(W461), .ZN(W2009));
  INVX1 G36415 (.I(W3618), .ZN(O17815));
  INVX1 G36416 (.I(W14591), .ZN(O17813));
  INVX1 G36417 (.I(W1912), .ZN(W2014));
  INVX1 G36418 (.I(W24804), .ZN(O17810));
  INVX1 G36419 (.I(W1540), .ZN(O17809));
  INVX1 G36420 (.I(W1058), .ZN(W2019));
  INVX1 G36421 (.I(W7), .ZN(W2021));
  INVX1 G36422 (.I(W44053), .ZN(O17803));
  INVX1 G36423 (.I(W7077), .ZN(O17819));
  INVX1 G36424 (.I(I1692), .ZN(W2024));
  INVX1 G36425 (.I(I809), .ZN(W2028));
  INVX1 G36426 (.I(W31197), .ZN(O17798));
  INVX1 G36427 (.I(W23943), .ZN(O17797));
  INVX1 G36428 (.I(W1010), .ZN(O17796));
  INVX1 G36429 (.I(I1684), .ZN(W2030));
  INVX1 G36430 (.I(W39), .ZN(W2033));
  INVX1 G36431 (.I(W1763), .ZN(W2038));
  INVX1 G36432 (.I(W7549), .ZN(O17831));
  INVX1 G36433 (.I(W7817), .ZN(O17844));
  INVX1 G36434 (.I(W39589), .ZN(O17843));
  INVX1 G36435 (.I(W514), .ZN(W1984));
  INVX1 G36436 (.I(I486), .ZN(W1985));
  INVX1 G36437 (.I(W656), .ZN(W1989));
  INVX1 G36438 (.I(W21086), .ZN(O17838));
  INVX1 G36439 (.I(W25874), .ZN(O17835));
  INVX1 G36440 (.I(W359), .ZN(W1993));
  INVX1 G36441 (.I(I690), .ZN(O17833));
  INVX1 G36442 (.I(I256), .ZN(W2039));
  INVX1 G36443 (.I(W3432), .ZN(O17830));
  INVX1 G36444 (.I(W23443), .ZN(O17829));
  INVX1 G36445 (.I(W135), .ZN(W1995));
  INVX1 G36446 (.I(W22073), .ZN(O17827));
  INVX1 G36447 (.I(W28072), .ZN(O17824));
  INVX1 G36448 (.I(I14), .ZN(W1998));
  INVX1 G36449 (.I(W531), .ZN(W2004));
  INVX1 G36450 (.I(W17695), .ZN(O17820));
  INVX1 G36451 (.I(W31831), .ZN(O17758));
  INVX1 G36452 (.I(W48537), .ZN(O17767));
  INVX1 G36453 (.I(W2010), .ZN(W2062));
  INVX1 G36454 (.I(W1572), .ZN(W2063));
  INVX1 G36455 (.I(W222), .ZN(W2064));
  INVX1 G36456 (.I(W957), .ZN(W2065));
  INVX1 G36457 (.I(W1780), .ZN(W2066));
  INVX1 G36458 (.I(W26168), .ZN(O17761));
  INVX1 G36459 (.I(I590), .ZN(W2068));
  INVX1 G36460 (.I(W31327), .ZN(O17759));
  INVX1 G36461 (.I(W18078), .ZN(O17770));
  INVX1 G36462 (.I(W44166), .ZN(O17757));
  INVX1 G36463 (.I(W1233), .ZN(W2069));
  INVX1 G36464 (.I(I1516), .ZN(W2070));
  INVX1 G36465 (.I(W1509), .ZN(W2071));
  INVX1 G36466 (.I(I825), .ZN(W2072));
  INVX1 G36467 (.I(I1546), .ZN(W2080));
  INVX1 G36468 (.I(W1832), .ZN(W2083));
  INVX1 G36469 (.I(W31735), .ZN(O17749));
  INVX1 G36470 (.I(W1060), .ZN(W2052));
  INVX1 G36471 (.I(W23841), .ZN(O17789));
  INVX1 G36472 (.I(W580), .ZN(W2042));
  INVX1 G36473 (.I(I1926), .ZN(W2044));
  INVX1 G36474 (.I(I1078), .ZN(W2045));
  INVX1 G36475 (.I(I1277), .ZN(W2046));
  INVX1 G36476 (.I(I1248), .ZN(W2048));
  INVX1 G36477 (.I(I1732), .ZN(W2050));
  INVX1 G36478 (.I(W36017), .ZN(O17781));
  INVX1 G36479 (.I(W1480), .ZN(W2659));
  INVX1 G36480 (.I(W28058), .ZN(O17779));
  INVX1 G36481 (.I(W637), .ZN(W2054));
  INVX1 G36482 (.I(I48), .ZN(W2057));
  INVX1 G36483 (.I(I1088), .ZN(W2058));
  INVX1 G36484 (.I(W22114), .ZN(O17774));
  INVX1 G36485 (.I(W11944), .ZN(O17773));
  INVX1 G36486 (.I(W4787), .ZN(O17772));
  INVX1 G36487 (.I(W943), .ZN(W2059));
  INVX1 G36488 (.I(W23300), .ZN(O16693));
  INVX1 G36489 (.I(I502), .ZN(W3202));
  INVX1 G36490 (.I(W33315), .ZN(O16701));
  INVX1 G36491 (.I(W44718), .ZN(W47758));
  INVX1 G36492 (.I(W11430), .ZN(O16700));
  INVX1 G36493 (.I(W41978), .ZN(O16699));
  INVX1 G36494 (.I(W33), .ZN(W3203));
  INVX1 G36495 (.I(W43516), .ZN(O16697));
  INVX1 G36496 (.I(W1273), .ZN(O16696));
  INVX1 G36497 (.I(W15441), .ZN(O16694));
  INVX1 G36498 (.I(W45890), .ZN(O16703));
  INVX1 G36499 (.I(W34916), .ZN(O16691));
  INVX1 G36500 (.I(W22250), .ZN(O16689));
  INVX1 G36501 (.I(W10136), .ZN(O16688));
  INVX1 G36502 (.I(W1171), .ZN(W3209));
  INVX1 G36503 (.I(W11999), .ZN(O16685));
  INVX1 G36504 (.I(W12201), .ZN(O16682));
  INVX1 G36505 (.I(W11687), .ZN(O16681));
  INVX1 G36506 (.I(W41064), .ZN(O16679));
  INVX1 G36507 (.I(W46299), .ZN(O16716));
  INVX1 G36508 (.I(I882), .ZN(O16727));
  INVX1 G36509 (.I(W975), .ZN(O16726));
  INVX1 G36510 (.I(W8391), .ZN(W47787));
  INVX1 G36511 (.I(I1586), .ZN(W3178));
  INVX1 G36512 (.I(W18268), .ZN(O16724));
  INVX1 G36513 (.I(W46210), .ZN(O16723));
  INVX1 G36514 (.I(W10525), .ZN(O16719));
  INVX1 G36515 (.I(I1066), .ZN(O16718));
  INVX1 G36516 (.I(I242), .ZN(W3186));
  INVX1 G36517 (.I(W11394), .ZN(O16675));
  INVX1 G36518 (.I(I710), .ZN(W3189));
  INVX1 G36519 (.I(W45525), .ZN(O16711));
  INVX1 G36520 (.I(I644), .ZN(W3194));
  INVX1 G36521 (.I(W24035), .ZN(O16707));
  INVX1 G36522 (.I(I1800), .ZN(W3198));
  INVX1 G36523 (.I(I798), .ZN(W3199));
  INVX1 G36524 (.I(W1779), .ZN(W3200));
  INVX1 G36525 (.I(I799), .ZN(W3201));
  INVX1 G36526 (.I(W248), .ZN(W3265));
  INVX1 G36527 (.I(W2097), .ZN(W3250));
  INVX1 G36528 (.I(I466), .ZN(W3252));
  INVX1 G36529 (.I(W19355), .ZN(O16646));
  INVX1 G36530 (.I(W40601), .ZN(O16645));
  INVX1 G36531 (.I(W1225), .ZN(W3257));
  INVX1 G36532 (.I(W2043), .ZN(W3259));
  INVX1 G36533 (.I(W36266), .ZN(O16640));
  INVX1 G36534 (.I(I445), .ZN(O31));
  INVX1 G36535 (.I(W25064), .ZN(O16636));
  INVX1 G36536 (.I(I368), .ZN(W3244));
  INVX1 G36537 (.I(W2324), .ZN(W3274));
  INVX1 G36538 (.I(I417), .ZN(W3276));
  INVX1 G36539 (.I(W1272), .ZN(W3277));
  INVX1 G36540 (.I(W1042), .ZN(W3279));
  INVX1 G36541 (.I(W32306), .ZN(O16626));
  INVX1 G36542 (.I(W47105), .ZN(O16625));
  INVX1 G36543 (.I(W831), .ZN(O16624));
  INVX1 G36544 (.I(W34708), .ZN(O16622));
  INVX1 G36545 (.I(I1633), .ZN(W3238));
  INVX1 G36546 (.I(W37330), .ZN(O16674));
  INVX1 G36547 (.I(I5), .ZN(O16671));
  INVX1 G36548 (.I(W1117), .ZN(W3229));
  INVX1 G36549 (.I(W9997), .ZN(O16668));
  INVX1 G36550 (.I(I56), .ZN(W3232));
  INVX1 G36551 (.I(W1761), .ZN(W3234));
  INVX1 G36552 (.I(I1739), .ZN(W3235));
  INVX1 G36553 (.I(I1142), .ZN(O16663));
  INVX1 G36554 (.I(W2441), .ZN(W3176));
  INVX1 G36555 (.I(W2722), .ZN(O16661));
  INVX1 G36556 (.I(W17970), .ZN(O16660));
  INVX1 G36557 (.I(W7185), .ZN(O16659));
  INVX1 G36558 (.I(I36), .ZN(W3239));
  INVX1 G36559 (.I(W1834), .ZN(W3240));
  INVX1 G36560 (.I(W37566), .ZN(O16656));
  INVX1 G36561 (.I(W557), .ZN(W3242));
  INVX1 G36562 (.I(I121), .ZN(W3243));
  INVX1 G36563 (.I(W15073), .ZN(O16783));
  INVX1 G36564 (.I(W1562), .ZN(W3115));
  INVX1 G36565 (.I(W790), .ZN(W3116));
  INVX1 G36566 (.I(W851), .ZN(O16791));
  INVX1 G36567 (.I(I171), .ZN(W3120));
  INVX1 G36568 (.I(W457), .ZN(W3121));
  INVX1 G36569 (.I(I1446), .ZN(W3126));
  INVX1 G36570 (.I(W47338), .ZN(W47853));
  INVX1 G36571 (.I(W8773), .ZN(O16786));
  INVX1 G36572 (.I(W17657), .ZN(O16785));
  INVX1 G36573 (.I(W2710), .ZN(W3112));
  INVX1 G36574 (.I(W15807), .ZN(O16782));
  INVX1 G36575 (.I(W30420), .ZN(O16781));
  INVX1 G36576 (.I(W28487), .ZN(O16780));
  INVX1 G36577 (.I(W1039), .ZN(O16779));
  INVX1 G36578 (.I(W9745), .ZN(O16777));
  INVX1 G36579 (.I(W8179), .ZN(O16776));
  INVX1 G36580 (.I(I1265), .ZN(W3130));
  INVX1 G36581 (.I(I1808), .ZN(W3132));
  INVX1 G36582 (.I(W23245), .ZN(O16806));
  INVX1 G36583 (.I(W678), .ZN(W3089));
  INVX1 G36584 (.I(W734), .ZN(W3091));
  INVX1 G36585 (.I(W28476), .ZN(W47886));
  INVX1 G36586 (.I(W17608), .ZN(O16815));
  INVX1 G36587 (.I(W29721), .ZN(W47884));
  INVX1 G36588 (.I(I1754), .ZN(W3092));
  INVX1 G36589 (.I(W32698), .ZN(O16812));
  INVX1 G36590 (.I(W1144), .ZN(W3096));
  INVX1 G36591 (.I(I1281), .ZN(W3098));
  INVX1 G36592 (.I(W578), .ZN(W3136));
  INVX1 G36593 (.I(W1636), .ZN(W3101));
  INVX1 G36594 (.I(W46928), .ZN(O16804));
  INVX1 G36595 (.I(I860), .ZN(O16802));
  INVX1 G36596 (.I(I1793), .ZN(W3109));
  INVX1 G36597 (.I(W39206), .ZN(O16799));
  INVX1 G36598 (.I(W754), .ZN(W3110));
  INVX1 G36599 (.I(W20454), .ZN(O16796));
  INVX1 G36600 (.I(W20142), .ZN(O16795));
  INVX1 G36601 (.I(W167), .ZN(W3171));
  INVX1 G36602 (.I(W41018), .ZN(O16750));
  INVX1 G36603 (.I(W4135), .ZN(O16749));
  INVX1 G36604 (.I(W39618), .ZN(O16748));
  INVX1 G36605 (.I(I694), .ZN(W3163));
  INVX1 G36606 (.I(W32500), .ZN(O16745));
  INVX1 G36607 (.I(W1054), .ZN(W3164));
  INVX1 G36608 (.I(W1532), .ZN(W3166));
  INVX1 G36609 (.I(I1199), .ZN(W3168));
  INVX1 G36610 (.I(W34117), .ZN(O16740));
  INVX1 G36611 (.I(W18963), .ZN(O16751));
  INVX1 G36612 (.I(W13527), .ZN(O16738));
  INVX1 G36613 (.I(W38115), .ZN(O16737));
  INVX1 G36614 (.I(W10165), .ZN(O16736));
  INVX1 G36615 (.I(W39271), .ZN(O16734));
  INVX1 G36616 (.I(I1563), .ZN(O16733));
  INVX1 G36617 (.I(W2338), .ZN(W3173));
  INVX1 G36618 (.I(I1321), .ZN(W3174));
  INVX1 G36619 (.I(W42541), .ZN(O16730));
  INVX1 G36620 (.I(W10884), .ZN(O16760));
  INVX1 G36621 (.I(W2615), .ZN(O16772));
  INVX1 G36622 (.I(W2716), .ZN(W3137));
  INVX1 G36623 (.I(W1428), .ZN(W3141));
  INVX1 G36624 (.I(W5838), .ZN(O16768));
  INVX1 G36625 (.I(W43950), .ZN(O16767));
  INVX1 G36626 (.I(I1685), .ZN(O16766));
  INVX1 G36627 (.I(W15983), .ZN(O16765));
  INVX1 G36628 (.I(W45269), .ZN(O16762));
  INVX1 G36629 (.I(W41207), .ZN(O16621));
  INVX1 G36630 (.I(W11), .ZN(W3149));
  INVX1 G36631 (.I(W1222), .ZN(W3151));
  INVX1 G36632 (.I(I536), .ZN(W3153));
  INVX1 G36633 (.I(W1867), .ZN(W3154));
  INVX1 G36634 (.I(W1992), .ZN(W3156));
  INVX1 G36635 (.I(W24809), .ZN(O16755));
  INVX1 G36636 (.I(W1107), .ZN(W3157));
  INVX1 G36637 (.I(W45570), .ZN(O16752));
  INVX1 G36638 (.I(W1597), .ZN(W47518));
  INVX1 G36639 (.I(W2135), .ZN(W3439));
  INVX1 G36640 (.I(I747), .ZN(W3442));
  INVX1 G36641 (.I(W2453), .ZN(W3443));
  INVX1 G36642 (.I(W37718), .ZN(O16492));
  INVX1 G36643 (.I(W1977), .ZN(W3446));
  INVX1 G36644 (.I(W9044), .ZN(O16489));
  INVX1 G36645 (.I(W2042), .ZN(W3452));
  INVX1 G36646 (.I(W762), .ZN(O16485));
  INVX1 G36647 (.I(W1851), .ZN(W3455));
  INVX1 G36648 (.I(W1320), .ZN(O16497));
  INVX1 G36649 (.I(W374), .ZN(W3458));
  INVX1 G36650 (.I(W38056), .ZN(O16478));
  INVX1 G36651 (.I(W1947), .ZN(W3464));
  INVX1 G36652 (.I(W22477), .ZN(O16476));
  INVX1 G36653 (.I(W2525), .ZN(W3468));
  INVX1 G36654 (.I(W37715), .ZN(O16472));
  INVX1 G36655 (.I(W26480), .ZN(W47504));
  INVX1 G36656 (.I(W15712), .ZN(W47501));
  INVX1 G36657 (.I(W22411), .ZN(O16510));
  INVX1 G36658 (.I(I1884), .ZN(W3406));
  INVX1 G36659 (.I(W2432), .ZN(W3408));
  INVX1 G36660 (.I(W25450), .ZN(O16517));
  INVX1 G36661 (.I(I1988), .ZN(W3410));
  INVX1 G36662 (.I(W710), .ZN(W3413));
  INVX1 G36663 (.I(W38025), .ZN(O16515));
  INVX1 G36664 (.I(I1389), .ZN(W3415));
  INVX1 G36665 (.I(W2807), .ZN(W3419));
  INVX1 G36666 (.I(W21469), .ZN(O16511));
  INVX1 G36667 (.I(W2078), .ZN(W3477));
  INVX1 G36668 (.I(W24833), .ZN(O16509));
  INVX1 G36669 (.I(W12878), .ZN(W47547));
  INVX1 G36670 (.I(I1585), .ZN(W3426));
  INVX1 G36671 (.I(W12615), .ZN(O16503));
  INVX1 G36672 (.I(W35522), .ZN(O16500));
  INVX1 G36673 (.I(I1215), .ZN(W3438));
  INVX1 G36674 (.I(W29155), .ZN(O16499));
  INVX1 G36675 (.I(W9589), .ZN(O16498));
  INVX1 G36676 (.I(W2651), .ZN(W3506));
  INVX1 G36677 (.I(W14007), .ZN(O16444));
  INVX1 G36678 (.I(W951), .ZN(W3500));
  INVX1 G36679 (.I(W4110), .ZN(O16441));
  INVX1 G36680 (.I(W250), .ZN(W3501));
  INVX1 G36681 (.I(I608), .ZN(W3502));
  INVX1 G36682 (.I(W377), .ZN(W3504));
  INVX1 G36683 (.I(W44249), .ZN(O16436));
  INVX1 G36684 (.I(W17495), .ZN(O16435));
  INVX1 G36685 (.I(W36850), .ZN(O16434));
  INVX1 G36686 (.I(W603), .ZN(W3498));
  INVX1 G36687 (.I(W561), .ZN(W3508));
  INVX1 G36688 (.I(W2523), .ZN(O16430));
  INVX1 G36689 (.I(W25523), .ZN(O16428));
  INVX1 G36690 (.I(I1924), .ZN(W3511));
  INVX1 G36691 (.I(W2305), .ZN(W3514));
  INVX1 G36692 (.I(W33254), .ZN(O16424));
  INVX1 G36693 (.I(W1689), .ZN(W3516));
  INVX1 G36694 (.I(W2185), .ZN(W3519));
  INVX1 G36695 (.I(W31074), .ZN(O16456));
  INVX1 G36696 (.I(W1551), .ZN(W3478));
  INVX1 G36697 (.I(W2101), .ZN(W3480));
  INVX1 G36698 (.I(W10756), .ZN(O16463));
  INVX1 G36699 (.I(W14577), .ZN(O16462));
  INVX1 G36700 (.I(W18796), .ZN(O16461));
  INVX1 G36701 (.I(W28164), .ZN(O16460));
  INVX1 G36702 (.I(W1960), .ZN(O16458));
  INVX1 G36703 (.I(W2013), .ZN(O16457));
  INVX1 G36704 (.I(W3212), .ZN(W3405));
  INVX1 G36705 (.I(W39406), .ZN(O16455));
  INVX1 G36706 (.I(I746), .ZN(O36));
  INVX1 G36707 (.I(W10581), .ZN(O16451));
  INVX1 G36708 (.I(I1851), .ZN(O37));
  INVX1 G36709 (.I(W14644), .ZN(O16449));
  INVX1 G36710 (.I(W554), .ZN(W3495));
  INVX1 G36711 (.I(W2466), .ZN(W3497));
  INVX1 G36712 (.I(W33292), .ZN(O16446));
  INVX1 G36713 (.I(W2598), .ZN(W3334));
  INVX1 G36714 (.I(W6190), .ZN(O16596));
  INVX1 G36715 (.I(I1852), .ZN(W3314));
  INVX1 G36716 (.I(I655), .ZN(W3316));
  INVX1 G36717 (.I(W44824), .ZN(O16593));
  INVX1 G36718 (.I(W19101), .ZN(O16590));
  INVX1 G36719 (.I(W230), .ZN(W3327));
  INVX1 G36720 (.I(W27667), .ZN(O16584));
  INVX1 G36721 (.I(W45656), .ZN(O16582));
  INVX1 G36722 (.I(I830), .ZN(W47632));
  INVX1 G36723 (.I(W1907), .ZN(W3311));
  INVX1 G36724 (.I(W3184), .ZN(W3336));
  INVX1 G36725 (.I(I1380), .ZN(W3339));
  INVX1 G36726 (.I(W1887), .ZN(W3340));
  INVX1 G36727 (.I(W38085), .ZN(W47624));
  INVX1 G36728 (.I(W802), .ZN(W3344));
  INVX1 G36729 (.I(W14754), .ZN(O16574));
  INVX1 G36730 (.I(W15093), .ZN(O16572));
  INVX1 G36731 (.I(W883), .ZN(W3350));
  INVX1 G36732 (.I(W26088), .ZN(O16611));
  INVX1 G36733 (.I(W6904), .ZN(W47675));
  INVX1 G36734 (.I(W2180), .ZN(W3282));
  INVX1 G36735 (.I(W2707), .ZN(W3283));
  INVX1 G36736 (.I(I1044), .ZN(W3284));
  INVX1 G36737 (.I(W2232), .ZN(W3288));
  INVX1 G36738 (.I(W764), .ZN(W3291));
  INVX1 G36739 (.I(W33280), .ZN(O16613));
  INVX1 G36740 (.I(I1029), .ZN(W3292));
  INVX1 G36741 (.I(W1476), .ZN(W3293));
  INVX1 G36742 (.I(I1730), .ZN(W3352));
  INVX1 G36743 (.I(W47057), .ZN(O16609));
  INVX1 G36744 (.I(W3008), .ZN(W3295));
  INVX1 G36745 (.I(I1339), .ZN(W3297));
  INVX1 G36746 (.I(W1702), .ZN(W3299));
  INVX1 G36747 (.I(W910), .ZN(W3303));
  INVX1 G36748 (.I(W555), .ZN(W3306));
  INVX1 G36749 (.I(W548), .ZN(W3307));
  INVX1 G36750 (.I(W31524), .ZN(O16599));
  INVX1 G36751 (.I(W1034), .ZN(W3388));
  INVX1 G36752 (.I(W1706), .ZN(O16546));
  INVX1 G36753 (.I(W17303), .ZN(O16545));
  INVX1 G36754 (.I(W46193), .ZN(O16544));
  INVX1 G36755 (.I(I316), .ZN(W3380));
  INVX1 G36756 (.I(I895), .ZN(W3381));
  INVX1 G36757 (.I(W1381), .ZN(W3385));
  INVX1 G36758 (.I(W38857), .ZN(O16536));
  INVX1 G36759 (.I(W31811), .ZN(O16535));
  INVX1 G36760 (.I(W24514), .ZN(O16534));
  INVX1 G36761 (.I(W538), .ZN(W3376));
  INVX1 G36762 (.I(I1367), .ZN(W3390));
  INVX1 G36763 (.I(W18459), .ZN(O16531));
  INVX1 G36764 (.I(I1120), .ZN(W3392));
  INVX1 G36765 (.I(W215), .ZN(W3396));
  INVX1 G36766 (.I(W2870), .ZN(W3398));
  INVX1 G36767 (.I(W2348), .ZN(W3400));
  INVX1 G36768 (.I(W10897), .ZN(O16523));
  INVX1 G36769 (.I(W2521), .ZN(W3403));
  INVX1 G36770 (.I(W30125), .ZN(O16562));
  INVX1 G36771 (.I(W11196), .ZN(O16569));
  INVX1 G36772 (.I(W386), .ZN(W3354));
  INVX1 G36773 (.I(W36959), .ZN(O16567));
  INVX1 G36774 (.I(W37144), .ZN(O16566));
  INVX1 G36775 (.I(W1678), .ZN(W3356));
  INVX1 G36776 (.I(I1240), .ZN(W3357));
  INVX1 G36777 (.I(W1430), .ZN(W3358));
  INVX1 G36778 (.I(W34273), .ZN(O16563));
  INVX1 G36779 (.I(W35206), .ZN(O16819));
  INVX1 G36780 (.I(I196), .ZN(W3359));
  INVX1 G36781 (.I(W26074), .ZN(O16560));
  INVX1 G36782 (.I(W2937), .ZN(W3364));
  INVX1 G36783 (.I(W3364), .ZN(W3365));
  INVX1 G36784 (.I(W46005), .ZN(O16552));
  INVX1 G36785 (.I(W956), .ZN(W3375));
  INVX1 G36786 (.I(W25981), .ZN(O16549));
  INVX1 G36787 (.I(W16296), .ZN(O16548));
  INVX1 G36788 (.I(I190), .ZN(W2791));
  INVX1 G36789 (.I(I502), .ZN(W2778));
  INVX1 G36790 (.I(W34189), .ZN(O17098));
  INVX1 G36791 (.I(W13298), .ZN(O17097));
  INVX1 G36792 (.I(I91), .ZN(W2781));
  INVX1 G36793 (.I(I492), .ZN(W2783));
  INVX1 G36794 (.I(W1985), .ZN(W2784));
  INVX1 G36795 (.I(W31205), .ZN(O17090));
  INVX1 G36796 (.I(W1139), .ZN(W2785));
  INVX1 G36797 (.I(W41422), .ZN(W48181));
  INVX1 G36798 (.I(W14631), .ZN(O17100));
  INVX1 G36799 (.I(I1949), .ZN(W2792));
  INVX1 G36800 (.I(W2437), .ZN(O17083));
  INVX1 G36801 (.I(W30199), .ZN(O17079));
  INVX1 G36802 (.I(W52), .ZN(W2797));
  INVX1 G36803 (.I(W45225), .ZN(O17077));
  INVX1 G36804 (.I(W2074), .ZN(W2801));
  INVX1 G36805 (.I(I1966), .ZN(W2806));
  INVX1 G36806 (.I(W629), .ZN(W2807));
  INVX1 G36807 (.I(W1812), .ZN(W2768));
  INVX1 G36808 (.I(W48181), .ZN(O17120));
  INVX1 G36809 (.I(I1644), .ZN(W2763));
  INVX1 G36810 (.I(I483), .ZN(W2764));
  INVX1 G36811 (.I(W44666), .ZN(O17116));
  INVX1 G36812 (.I(W30867), .ZN(O17115));
  INVX1 G36813 (.I(I1260), .ZN(W2767));
  INVX1 G36814 (.I(W10247), .ZN(O17113));
  INVX1 G36815 (.I(W40500), .ZN(O17112));
  INVX1 G36816 (.I(W37280), .ZN(W48207));
  INVX1 G36817 (.I(W16305), .ZN(O17070));
  INVX1 G36818 (.I(W6176), .ZN(O17110));
  INVX1 G36819 (.I(W12152), .ZN(O17109));
  INVX1 G36820 (.I(W841), .ZN(W2769));
  INVX1 G36821 (.I(I1720), .ZN(W2772));
  INVX1 G36822 (.I(W1889), .ZN(W2773));
  INVX1 G36823 (.I(W9592), .ZN(O17104));
  INVX1 G36824 (.I(W979), .ZN(W2774));
  INVX1 G36825 (.I(W888), .ZN(W2775));
  INVX1 G36826 (.I(W40408), .ZN(O17031));
  INVX1 G36827 (.I(W15961), .ZN(O17046));
  INVX1 G36828 (.I(W2446), .ZN(W2835));
  INVX1 G36829 (.I(W1769), .ZN(W2836));
  INVX1 G36830 (.I(I1284), .ZN(O17043));
  INVX1 G36831 (.I(W37770), .ZN(O17042));
  INVX1 G36832 (.I(I1021), .ZN(W2849));
  INVX1 G36833 (.I(I779), .ZN(W2850));
  INVX1 G36834 (.I(I1238), .ZN(W2854));
  INVX1 G36835 (.I(W1045), .ZN(W2858));
  INVX1 G36836 (.I(W132), .ZN(W2834));
  INVX1 G36837 (.I(W47226), .ZN(O17030));
  INVX1 G36838 (.I(W16869), .ZN(O17029));
  INVX1 G36839 (.I(W46357), .ZN(O17028));
  INVX1 G36840 (.I(W42), .ZN(W2859));
  INVX1 G36841 (.I(W990), .ZN(O17027));
  INVX1 G36842 (.I(I1988), .ZN(W2863));
  INVX1 G36843 (.I(W30526), .ZN(O17022));
  INVX1 G36844 (.I(W11721), .ZN(O17021));
  INVX1 G36845 (.I(W2203), .ZN(W2823));
  INVX1 G36846 (.I(W36131), .ZN(O17068));
  INVX1 G36847 (.I(W13824), .ZN(O17067));
  INVX1 G36848 (.I(W35229), .ZN(O17066));
  INVX1 G36849 (.I(W1554), .ZN(W2815));
  INVX1 G36850 (.I(W2473), .ZN(W2817));
  INVX1 G36851 (.I(I132), .ZN(W2818));
  INVX1 G36852 (.I(W10332), .ZN(O17060));
  INVX1 G36853 (.I(I1259), .ZN(W2822));
  INVX1 G36854 (.I(W39566), .ZN(O17121));
  INVX1 G36855 (.I(W14539), .ZN(O17056));
  INVX1 G36856 (.I(W16394), .ZN(O17055));
  INVX1 G36857 (.I(W35908), .ZN(O17054));
  INVX1 G36858 (.I(W27699), .ZN(O17051));
  INVX1 G36859 (.I(I574), .ZN(W2831));
  INVX1 G36860 (.I(I1506), .ZN(W2833));
  INVX1 G36861 (.I(W33961), .ZN(W48136));
  INVX1 G36862 (.I(W39396), .ZN(O17048));
  INVX1 G36863 (.I(W24004), .ZN(O17178));
  INVX1 G36864 (.I(W1827), .ZN(W2686));
  INVX1 G36865 (.I(W43003), .ZN(O17188));
  INVX1 G36866 (.I(W8481), .ZN(O17187));
  INVX1 G36867 (.I(W1122), .ZN(W2687));
  INVX1 G36868 (.I(W33389), .ZN(O17183));
  INVX1 G36869 (.I(W17610), .ZN(O17181));
  INVX1 G36870 (.I(I695), .ZN(W2696));
  INVX1 G36871 (.I(I1970), .ZN(W2697));
  INVX1 G36872 (.I(W2197), .ZN(W2698));
  INVX1 G36873 (.I(W7810), .ZN(O17190));
  INVX1 G36874 (.I(I1503), .ZN(W2699));
  INVX1 G36875 (.I(W2603), .ZN(W2700));
  INVX1 G36876 (.I(I238), .ZN(W2703));
  INVX1 G36877 (.I(W46826), .ZN(O17173));
  INVX1 G36878 (.I(W6136), .ZN(O17172));
  INVX1 G36879 (.I(I1468), .ZN(W2706));
  INVX1 G36880 (.I(W2975), .ZN(O17171));
  INVX1 G36881 (.I(W42288), .ZN(O17170));
  INVX1 G36882 (.I(W40), .ZN(W2672));
  INVX1 G36883 (.I(W12233), .ZN(O17216));
  INVX1 G36884 (.I(W41314), .ZN(O17215));
  INVX1 G36885 (.I(W6268), .ZN(O17213));
  INVX1 G36886 (.I(W1756), .ZN(W2664));
  INVX1 G36887 (.I(W34342), .ZN(O17210));
  INVX1 G36888 (.I(W2388), .ZN(W2667));
  INVX1 G36889 (.I(W17407), .ZN(O17206));
  INVX1 G36890 (.I(I1958), .ZN(W2669));
  INVX1 G36891 (.I(W46079), .ZN(O17204));
  INVX1 G36892 (.I(W1511), .ZN(W2708));
  INVX1 G36893 (.I(W15948), .ZN(O17201));
  INVX1 G36894 (.I(W11499), .ZN(O17200));
  INVX1 G36895 (.I(W5992), .ZN(O17199));
  INVX1 G36896 (.I(W1919), .ZN(W2673));
  INVX1 G36897 (.I(I161), .ZN(W2675));
  INVX1 G36898 (.I(W32212), .ZN(O17195));
  INVX1 G36899 (.I(W2541), .ZN(W2680));
  INVX1 G36900 (.I(W2570), .ZN(W2685));
  INVX1 G36901 (.I(W1907), .ZN(W48231));
  INVX1 G36902 (.I(I221), .ZN(O17148));
  INVX1 G36903 (.I(W7350), .ZN(O17147));
  INVX1 G36904 (.I(W45993), .ZN(O17146));
  INVX1 G36905 (.I(W29450), .ZN(O17145));
  INVX1 G36906 (.I(I428), .ZN(W2733));
  INVX1 G36907 (.I(W45788), .ZN(O17140));
  INVX1 G36908 (.I(W24388), .ZN(O17139));
  INVX1 G36909 (.I(W43380), .ZN(O17137));
  INVX1 G36910 (.I(W18731), .ZN(W48235));
  INVX1 G36911 (.I(W39129), .ZN(O17149));
  INVX1 G36912 (.I(W28125), .ZN(O17133));
  INVX1 G36913 (.I(W37307), .ZN(O17131));
  INVX1 G36914 (.I(I820), .ZN(W2744));
  INVX1 G36915 (.I(W1342), .ZN(W2748));
  INVX1 G36916 (.I(W1332), .ZN(W2755));
  INVX1 G36917 (.I(W960), .ZN(W2759));
  INVX1 G36918 (.I(W30116), .ZN(O17123));
  INVX1 G36919 (.I(I1350), .ZN(W2760));
  INVX1 G36920 (.I(W172), .ZN(W2725));
  INVX1 G36921 (.I(W406), .ZN(W2711));
  INVX1 G36922 (.I(I1069), .ZN(W2713));
  INVX1 G36923 (.I(W60), .ZN(W2716));
  INVX1 G36924 (.I(I1851), .ZN(W2722));
  INVX1 G36925 (.I(W2458), .ZN(W2723));
  INVX1 G36926 (.I(I1610), .ZN(O17160));
  INVX1 G36927 (.I(W26131), .ZN(O17159));
  INVX1 G36928 (.I(W28077), .ZN(O17158));
  INVX1 G36929 (.I(W1054), .ZN(W2865));
  INVX1 G36930 (.I(I1953), .ZN(W2726));
  INVX1 G36931 (.I(W34863), .ZN(O17155));
  INVX1 G36932 (.I(I229), .ZN(W2728));
  INVX1 G36933 (.I(I1225), .ZN(W2729));
  INVX1 G36934 (.I(W43221), .ZN(O17153));
  INVX1 G36935 (.I(W21376), .ZN(O17152));
  INVX1 G36936 (.I(W34959), .ZN(O17151));
  INVX1 G36937 (.I(I1671), .ZN(W2730));
  INVX1 G36938 (.I(W2161), .ZN(W3005));
  INVX1 G36939 (.I(W1516), .ZN(W2990));
  INVX1 G36940 (.I(W1459), .ZN(W2991));
  INVX1 G36941 (.I(I1108), .ZN(W2995));
  INVX1 G36942 (.I(I1571), .ZN(W2996));
  INVX1 G36943 (.I(I353), .ZN(W2998));
  INVX1 G36944 (.I(W38540), .ZN(O16891));
  INVX1 G36945 (.I(W35646), .ZN(W47968));
  INVX1 G36946 (.I(W1230), .ZN(W3001));
  INVX1 G36947 (.I(I1624), .ZN(W3002));
  INVX1 G36948 (.I(W1839), .ZN(W2989));
  INVX1 G36949 (.I(W38197), .ZN(O16887));
  INVX1 G36950 (.I(W4818), .ZN(O16884));
  INVX1 G36951 (.I(W2879), .ZN(O16883));
  INVX1 G36952 (.I(W32180), .ZN(O16880));
  INVX1 G36953 (.I(W2833), .ZN(W3019));
  INVX1 G36954 (.I(W1472), .ZN(W3021));
  INVX1 G36955 (.I(W46107), .ZN(O16875));
  INVX1 G36956 (.I(W12749), .ZN(O16874));
  INVX1 G36957 (.I(W46241), .ZN(O16915));
  INVX1 G36958 (.I(W10969), .ZN(O16928));
  INVX1 G36959 (.I(W650), .ZN(W2957));
  INVX1 G36960 (.I(W2636), .ZN(W2959));
  INVX1 G36961 (.I(I1277), .ZN(W2962));
  INVX1 G36962 (.I(W2162), .ZN(O16922));
  INVX1 G36963 (.I(I1619), .ZN(W2965));
  INVX1 G36964 (.I(W8061), .ZN(O16919));
  INVX1 G36965 (.I(W44403), .ZN(O16917));
  INVX1 G36966 (.I(W38360), .ZN(O16916));
  INVX1 G36967 (.I(W2674), .ZN(O16872));
  INVX1 G36968 (.I(W44753), .ZN(W47994));
  INVX1 G36969 (.I(W36139), .ZN(O16914));
  INVX1 G36970 (.I(I1011), .ZN(W2972));
  INVX1 G36971 (.I(W42653), .ZN(O16910));
  INVX1 G36972 (.I(W1744), .ZN(W2975));
  INVX1 G36973 (.I(I1578), .ZN(W2977));
  INVX1 G36974 (.I(W2127), .ZN(W2979));
  INVX1 G36975 (.I(W47510), .ZN(O16902));
  INVX1 G36976 (.I(W17477), .ZN(O16831));
  INVX1 G36977 (.I(I723), .ZN(W3061));
  INVX1 G36978 (.I(W639), .ZN(W3063));
  INVX1 G36979 (.I(I1150), .ZN(W3064));
  INVX1 G36980 (.I(W30635), .ZN(O16840));
  INVX1 G36981 (.I(W2090), .ZN(W3067));
  INVX1 G36982 (.I(W46587), .ZN(O16836));
  INVX1 G36983 (.I(W36245), .ZN(O16835));
  INVX1 G36984 (.I(W41072), .ZN(O16834));
  INVX1 G36985 (.I(I409), .ZN(W3070));
  INVX1 G36986 (.I(W38260), .ZN(O16845));
  INVX1 G36987 (.I(W1065), .ZN(O16829));
  INVX1 G36988 (.I(W2684), .ZN(W3082));
  INVX1 G36989 (.I(W9065), .ZN(O16824));
  INVX1 G36990 (.I(W34507), .ZN(O16823));
  INVX1 G36991 (.I(I764), .ZN(W3084));
  INVX1 G36992 (.I(I382), .ZN(W3085));
  INVX1 G36993 (.I(W3073), .ZN(W3087));
  INVX1 G36994 (.I(W893), .ZN(W3088));
  INVX1 G36995 (.I(W16), .ZN(W3045));
  INVX1 G36996 (.I(I992), .ZN(W3030));
  INVX1 G36997 (.I(W27549), .ZN(O16868));
  INVX1 G36998 (.I(W29976), .ZN(O16867));
  INVX1 G36999 (.I(W38675), .ZN(O16866));
  INVX1 G37000 (.I(W648), .ZN(W3033));
  INVX1 G37001 (.I(W47884), .ZN(O16864));
  INVX1 G37002 (.I(I1179), .ZN(W3037));
  INVX1 G37003 (.I(W2854), .ZN(W3038));
  INVX1 G37004 (.I(W45264), .ZN(O16929));
  INVX1 G37005 (.I(W43536), .ZN(O16858));
  INVX1 G37006 (.I(I1197), .ZN(W3046));
  INVX1 G37007 (.I(I259), .ZN(W3051));
  INVX1 G37008 (.I(W47385), .ZN(O16852));
  INVX1 G37009 (.I(W41784), .ZN(O16851));
  INVX1 G37010 (.I(W25045), .ZN(O16850));
  INVX1 G37011 (.I(W12686), .ZN(O16847));
  INVX1 G37012 (.I(W6886), .ZN(O16846));
  INVX1 G37013 (.I(W777), .ZN(W2897));
  INVX1 G37014 (.I(W979), .ZN(W2887));
  INVX1 G37015 (.I(W877), .ZN(W2890));
  INVX1 G37016 (.I(W33790), .ZN(O16993));
  INVX1 G37017 (.I(W1088), .ZN(W2891));
  INVX1 G37018 (.I(W2036), .ZN(W2892));
  INVX1 G37019 (.I(W960), .ZN(W2893));
  INVX1 G37020 (.I(W363), .ZN(W2895));
  INVX1 G37021 (.I(W5118), .ZN(O16990));
  INVX1 G37022 (.I(I1118), .ZN(W2896));
  INVX1 G37023 (.I(W39988), .ZN(O16997));
  INVX1 G37024 (.I(W27826), .ZN(O16987));
  INVX1 G37025 (.I(W1257), .ZN(W2899));
  INVX1 G37026 (.I(W36187), .ZN(O16984));
  INVX1 G37027 (.I(W24715), .ZN(O16983));
  INVX1 G37028 (.I(W1120), .ZN(W2902));
  INVX1 G37029 (.I(I1820), .ZN(W2904));
  INVX1 G37030 (.I(W3356), .ZN(O16981));
  INVX1 G37031 (.I(W847), .ZN(W2906));
  INVX1 G37032 (.I(I1172), .ZN(W2877));
  INVX1 G37033 (.I(W27519), .ZN(O17019));
  INVX1 G37034 (.I(W568), .ZN(W2869));
  INVX1 G37035 (.I(W4244), .ZN(O17017));
  INVX1 G37036 (.I(I1064), .ZN(W2871));
  INVX1 G37037 (.I(W43291), .ZN(O17015));
  INVX1 G37038 (.I(W1393), .ZN(O17014));
  INVX1 G37039 (.I(W35512), .ZN(O17012));
  INVX1 G37040 (.I(W11349), .ZN(O17011));
  INVX1 G37041 (.I(I1687), .ZN(W2875));
  INVX1 G37042 (.I(W12885), .ZN(O16978));
  INVX1 G37043 (.I(W18692), .ZN(O17007));
  INVX1 G37044 (.I(I633), .ZN(O17006));
  INVX1 G37045 (.I(W5612), .ZN(O17005));
  INVX1 G37046 (.I(I1461), .ZN(W2879));
  INVX1 G37047 (.I(W26693), .ZN(O17002));
  INVX1 G37048 (.I(W72), .ZN(W2883));
  INVX1 G37049 (.I(W836), .ZN(W2885));
  INVX1 G37050 (.I(W39748), .ZN(O16999));
  INVX1 G37051 (.I(I204), .ZN(W2946));
  INVX1 G37052 (.I(W16184), .ZN(O16953));
  INVX1 G37053 (.I(W2210), .ZN(W2929));
  INVX1 G37054 (.I(W134), .ZN(W2931));
  INVX1 G37055 (.I(I1853), .ZN(W2932));
  INVX1 G37056 (.I(W37695), .ZN(O16947));
  INVX1 G37057 (.I(I24), .ZN(W2936));
  INVX1 G37058 (.I(W2898), .ZN(W2937));
  INVX1 G37059 (.I(I700), .ZN(W2940));
  INVX1 G37060 (.I(W2160), .ZN(W2942));
  INVX1 G37061 (.I(W10626), .ZN(O16954));
  INVX1 G37062 (.I(W2226), .ZN(W2947));
  INVX1 G37063 (.I(W46814), .ZN(O16939));
  INVX1 G37064 (.I(W43658), .ZN(O16938));
  INVX1 G37065 (.I(W40871), .ZN(O16937));
  INVX1 G37066 (.I(I1956), .ZN(W2948));
  INVX1 G37067 (.I(W2635), .ZN(W2953));
  INVX1 G37068 (.I(W2245), .ZN(W2954));
  INVX1 G37069 (.I(W47933), .ZN(O16931));
  INVX1 G37070 (.I(W949), .ZN(W2918));
  INVX1 G37071 (.I(W1012), .ZN(W2909));
  INVX1 G37072 (.I(W21545), .ZN(O16976));
  INVX1 G37073 (.I(W31315), .ZN(O16975));
  INVX1 G37074 (.I(W23441), .ZN(O16974));
  INVX1 G37075 (.I(W39271), .ZN(O16970));
  INVX1 G37076 (.I(W1542), .ZN(W2916));
  INVX1 G37077 (.I(I983), .ZN(W2917));
  INVX1 G37078 (.I(W16062), .ZN(O16967));
  INVX1 G37079 (.I(I818), .ZN(W1771));
  INVX1 G37080 (.I(I987), .ZN(W2919));
  INVX1 G37081 (.I(W34857), .ZN(O16964));
  INVX1 G37082 (.I(W34784), .ZN(O16963));
  INVX1 G37083 (.I(W2475), .ZN(W2921));
  INVX1 G37084 (.I(W30845), .ZN(O16960));
  INVX1 G37085 (.I(W43361), .ZN(O16959));
  INVX1 G37086 (.I(W2374), .ZN(W2924));
  INVX1 G37087 (.I(W14036), .ZN(O16955));
  INVX1 G37088 (.I(I1236), .ZN(W618));
  INVX1 G37089 (.I(I1202), .ZN(W601));
  INVX1 G37090 (.I(I1204), .ZN(W602));
  INVX1 G37091 (.I(W33592), .ZN(O19174));
  INVX1 G37092 (.I(I1206), .ZN(W603));
  INVX1 G37093 (.I(W4303), .ZN(O19171));
  INVX1 G37094 (.I(W32734), .ZN(O19168));
  INVX1 G37095 (.I(I1222), .ZN(W611));
  INVX1 G37096 (.I(W46239), .ZN(O19165));
  INVX1 G37097 (.I(I1226), .ZN(W613));
  INVX1 G37098 (.I(W367), .ZN(W50410));
  INVX1 G37099 (.I(I1240), .ZN(W620));
  INVX1 G37100 (.I(I1248), .ZN(W624));
  INVX1 G37101 (.I(I1256), .ZN(W628));
  INVX1 G37102 (.I(W29475), .ZN(O19157));
  INVX1 G37103 (.I(W15286), .ZN(O19156));
  INVX1 G37104 (.I(W46811), .ZN(O19155));
  INVX1 G37105 (.I(W7350), .ZN(O19154));
  INVX1 G37106 (.I(W37029), .ZN(O19152));
  INVX1 G37107 (.I(I1182), .ZN(W591));
  INVX1 G37108 (.I(W18893), .ZN(O19209));
  INVX1 G37109 (.I(W30910), .ZN(O19205));
  INVX1 G37110 (.I(I1154), .ZN(W577));
  INVX1 G37111 (.I(W43967), .ZN(O19203));
  INVX1 G37112 (.I(W30779), .ZN(O19202));
  INVX1 G37113 (.I(I1168), .ZN(W584));
  INVX1 G37114 (.I(W47514), .ZN(O19195));
  INVX1 G37115 (.I(W25044), .ZN(O19193));
  INVX1 G37116 (.I(W47384), .ZN(O19192));
  INVX1 G37117 (.I(W23256), .ZN(O19151));
  INVX1 G37118 (.I(W28617), .ZN(O19190));
  INVX1 G37119 (.I(I1184), .ZN(W592));
  INVX1 G37120 (.I(W22048), .ZN(O19188));
  INVX1 G37121 (.I(W20698), .ZN(O19187));
  INVX1 G37122 (.I(W21799), .ZN(O19185));
  INVX1 G37123 (.I(W40630), .ZN(O19184));
  INVX1 G37124 (.I(W3033), .ZN(O19182));
  INVX1 G37125 (.I(I1190), .ZN(W595));
  INVX1 G37126 (.I(I1358), .ZN(W679));
  INVX1 G37127 (.I(W34974), .ZN(O19120));
  INVX1 G37128 (.I(W14733), .ZN(O19118));
  INVX1 G37129 (.I(I1326), .ZN(W663));
  INVX1 G37130 (.I(W17293), .ZN(O19115));
  INVX1 G37131 (.I(W14766), .ZN(O19112));
  INVX1 G37132 (.I(I1334), .ZN(W667));
  INVX1 G37133 (.I(I1348), .ZN(W674));
  INVX1 G37134 (.I(I1350), .ZN(W675));
  INVX1 G37135 (.I(W12013), .ZN(O19101));
  INVX1 G37136 (.I(I1314), .ZN(W657));
  INVX1 G37137 (.I(I1362), .ZN(W681));
  INVX1 G37138 (.I(W22038), .ZN(O19097));
  INVX1 G37139 (.I(I1368), .ZN(W684));
  INVX1 G37140 (.I(I1370), .ZN(W685));
  INVX1 G37141 (.I(W38782), .ZN(O19094));
  INVX1 G37142 (.I(W24952), .ZN(O19093));
  INVX1 G37143 (.I(W33234), .ZN(O19092));
  INVX1 G37144 (.I(W23648), .ZN(O19089));
  INVX1 G37145 (.I(W11834), .ZN(O19135));
  INVX1 G37146 (.I(W8913), .ZN(O19149));
  INVX1 G37147 (.I(I1268), .ZN(W634));
  INVX1 G37148 (.I(I1274), .ZN(W637));
  INVX1 G37149 (.I(I1278), .ZN(W639));
  INVX1 G37150 (.I(W38524), .ZN(O19142));
  INVX1 G37151 (.I(I1284), .ZN(W642));
  INVX1 G37152 (.I(W38067), .ZN(O19139));
  INVX1 G37153 (.I(W18513), .ZN(O19138));
  INVX1 G37154 (.I(I1290), .ZN(W645));
  INVX1 G37155 (.I(I1136), .ZN(W568));
  INVX1 G37156 (.I(I1294), .ZN(W647));
  INVX1 G37157 (.I(W34441), .ZN(O19133));
  INVX1 G37158 (.I(I1296), .ZN(W648));
  INVX1 G37159 (.I(W36344), .ZN(O19127));
  INVX1 G37160 (.I(I1308), .ZN(W654));
  INVX1 G37161 (.I(I1310), .ZN(W655));
  INVX1 G37162 (.I(W34622), .ZN(O19124));
  INVX1 G37163 (.I(I1312), .ZN(W656));
  INVX1 G37164 (.I(I970), .ZN(W485));
  INVX1 G37165 (.I(I954), .ZN(W477));
  INVX1 G37166 (.I(I958), .ZN(W479));
  INVX1 G37167 (.I(W46415), .ZN(O19296));
  INVX1 G37168 (.I(I960), .ZN(W480));
  INVX1 G37169 (.I(W5407), .ZN(O19294));
  INVX1 G37170 (.I(W48836), .ZN(O19292));
  INVX1 G37171 (.I(W25239), .ZN(O19291));
  INVX1 G37172 (.I(W7407), .ZN(O19290));
  INVX1 G37173 (.I(W15070), .ZN(O19289));
  INVX1 G37174 (.I(W49087), .ZN(O19300));
  INVX1 G37175 (.I(W45710), .ZN(O19284));
  INVX1 G37176 (.I(I978), .ZN(W489));
  INVX1 G37177 (.I(I984), .ZN(W492));
  INVX1 G37178 (.I(W36944), .ZN(O19276));
  INVX1 G37179 (.I(I996), .ZN(W498));
  INVX1 G37180 (.I(W10807), .ZN(O19273));
  INVX1 G37181 (.I(W30229), .ZN(O19271));
  INVX1 G37182 (.I(I1006), .ZN(W503));
  INVX1 G37183 (.I(I898), .ZN(W449));
  INVX1 G37184 (.I(I868), .ZN(W434));
  INVX1 G37185 (.I(W36344), .ZN(O19332));
  INVX1 G37186 (.I(W39045), .ZN(O19330));
  INVX1 G37187 (.I(W14048), .ZN(O19329));
  INVX1 G37188 (.I(W34573), .ZN(O19328));
  INVX1 G37189 (.I(W8967), .ZN(O19326));
  INVX1 G37190 (.I(I882), .ZN(W441));
  INVX1 G37191 (.I(I890), .ZN(W445));
  INVX1 G37192 (.I(I896), .ZN(W448));
  INVX1 G37193 (.I(I1008), .ZN(W504));
  INVX1 G37194 (.I(W28406), .ZN(O19315));
  INVX1 G37195 (.I(I930), .ZN(W465));
  INVX1 G37196 (.I(W2804), .ZN(O19310));
  INVX1 G37197 (.I(W43605), .ZN(O19309));
  INVX1 G37198 (.I(W44209), .ZN(O19308));
  INVX1 G37199 (.I(I934), .ZN(W467));
  INVX1 G37200 (.I(I948), .ZN(W474));
  INVX1 G37201 (.I(I950), .ZN(W475));
  INVX1 G37202 (.I(I1096), .ZN(W548));
  INVX1 G37203 (.I(W13633), .ZN(O19239));
  INVX1 G37204 (.I(I1070), .ZN(W535));
  INVX1 G37205 (.I(I1076), .ZN(W538));
  INVX1 G37206 (.I(I1080), .ZN(W540));
  INVX1 G37207 (.I(I1082), .ZN(W541));
  INVX1 G37208 (.I(I1084), .ZN(W542));
  INVX1 G37209 (.I(W4015), .ZN(O19231));
  INVX1 G37210 (.I(W8042), .ZN(O19229));
  INVX1 G37211 (.I(I1092), .ZN(W546));
  INVX1 G37212 (.I(I1062), .ZN(W531));
  INVX1 G37213 (.I(I1098), .ZN(W549));
  INVX1 G37214 (.I(I1100), .ZN(W550));
  INVX1 G37215 (.I(I1478), .ZN(O19223));
  INVX1 G37216 (.I(I1108), .ZN(W554));
  INVX1 G37217 (.I(W9833), .ZN(O19219));
  INVX1 G37218 (.I(I1684), .ZN(O19216));
  INVX1 G37219 (.I(I1124), .ZN(W562));
  INVX1 G37220 (.I(W50225), .ZN(O19211));
  INVX1 G37221 (.I(I1038), .ZN(W519));
  INVX1 G37222 (.I(I1016), .ZN(W508));
  INVX1 G37223 (.I(I1022), .ZN(W511));
  INVX1 G37224 (.I(W13689), .ZN(O19264));
  INVX1 G37225 (.I(I1034), .ZN(W517));
  INVX1 G37226 (.I(W48727), .ZN(O19261));
  INVX1 G37227 (.I(I1036), .ZN(W518));
  INVX1 G37228 (.I(W8038), .ZN(O19259));
  INVX1 G37229 (.I(W7704), .ZN(O19258));
  INVX1 G37230 (.I(I1378), .ZN(W689));
  INVX1 G37231 (.I(W20051), .ZN(O19254));
  INVX1 G37232 (.I(W16567), .ZN(O19253));
  INVX1 G37233 (.I(W5433), .ZN(O19251));
  INVX1 G37234 (.I(I1056), .ZN(W528));
  INVX1 G37235 (.I(W30885), .ZN(O19245));
  INVX1 G37236 (.I(W17988), .ZN(O19243));
  INVX1 G37237 (.I(I1060), .ZN(W530));
  INVX1 G37238 (.I(W35601), .ZN(O19241));
  INVX1 G37239 (.I(W8174), .ZN(O18938));
  INVX1 G37240 (.I(W45383), .ZN(O18952));
  INVX1 G37241 (.I(I1634), .ZN(W817));
  INVX1 G37242 (.I(I1640), .ZN(W820));
  INVX1 G37243 (.I(I1642), .ZN(W821));
  INVX1 G37244 (.I(I1644), .ZN(W822));
  INVX1 G37245 (.I(I1654), .ZN(W827));
  INVX1 G37246 (.I(W3678), .ZN(O18944));
  INVX1 G37247 (.I(I1660), .ZN(W830));
  INVX1 G37248 (.I(W34935), .ZN(O18942));
  INVX1 G37249 (.I(I1630), .ZN(W815));
  INVX1 G37250 (.I(W36556), .ZN(O18936));
  INVX1 G37251 (.I(I1672), .ZN(W836));
  INVX1 G37252 (.I(W3334), .ZN(O18933));
  INVX1 G37253 (.I(I1682), .ZN(W841));
  INVX1 G37254 (.I(W1584), .ZN(O18930));
  INVX1 G37255 (.I(I1690), .ZN(W845));
  INVX1 G37256 (.I(I1692), .ZN(W846));
  INVX1 G37257 (.I(W3314), .ZN(O18925));
  INVX1 G37258 (.I(I1600), .ZN(W800));
  INVX1 G37259 (.I(W3120), .ZN(O18978));
  INVX1 G37260 (.I(W13227), .ZN(O18977));
  INVX1 G37261 (.I(W29915), .ZN(O18976));
  INVX1 G37262 (.I(I1582), .ZN(W791));
  INVX1 G37263 (.I(I1586), .ZN(W793));
  INVX1 G37264 (.I(W15240), .ZN(O18971));
  INVX1 G37265 (.I(I1594), .ZN(W797));
  INVX1 G37266 (.I(W7774), .ZN(O18969));
  INVX1 G37267 (.I(W13256), .ZN(O18968));
  INVX1 G37268 (.I(I1698), .ZN(W849));
  INVX1 G37269 (.I(W5650), .ZN(O18966));
  INVX1 G37270 (.I(I1604), .ZN(W802));
  INVX1 G37271 (.I(I1606), .ZN(W803));
  INVX1 G37272 (.I(I1612), .ZN(W806));
  INVX1 G37273 (.I(I1614), .ZN(W807));
  INVX1 G37274 (.I(I1622), .ZN(W811));
  INVX1 G37275 (.I(I1624), .ZN(W812));
  INVX1 G37276 (.I(I1626), .ZN(W813));
  INVX1 G37277 (.I(I1790), .ZN(W895));
  INVX1 G37278 (.I(I1766), .ZN(W883));
  INVX1 G37279 (.I(I1770), .ZN(W885));
  INVX1 G37280 (.I(I1780), .ZN(W890));
  INVX1 G37281 (.I(I1784), .ZN(W892));
  INVX1 G37282 (.I(I1786), .ZN(W893));
  INVX1 G37283 (.I(W25705), .ZN(O18884));
  INVX1 G37284 (.I(W24137), .ZN(O18883));
  INVX1 G37285 (.I(W7588), .ZN(W50105));
  INVX1 G37286 (.I(I1788), .ZN(W894));
  INVX1 G37287 (.I(I1764), .ZN(W882));
  INVX1 G37288 (.I(I1796), .ZN(W898));
  INVX1 G37289 (.I(I1804), .ZN(W902));
  INVX1 G37290 (.I(W33182), .ZN(O18875));
  INVX1 G37291 (.I(W3917), .ZN(O18870));
  INVX1 G37292 (.I(W1596), .ZN(O18868));
  INVX1 G37293 (.I(W43291), .ZN(O18867));
  INVX1 G37294 (.I(I1816), .ZN(W908));
  INVX1 G37295 (.I(I1820), .ZN(W910));
  INVX1 G37296 (.I(W6887), .ZN(O18907));
  INVX1 G37297 (.I(I1704), .ZN(W852));
  INVX1 G37298 (.I(I1712), .ZN(W856));
  INVX1 G37299 (.I(W29489), .ZN(O18917));
  INVX1 G37300 (.I(W20245), .ZN(O18916));
  INVX1 G37301 (.I(I1720), .ZN(W860));
  INVX1 G37302 (.I(I1722), .ZN(W861));
  INVX1 G37303 (.I(W44942), .ZN(O18911));
  INVX1 G37304 (.I(I1734), .ZN(W867));
  INVX1 G37305 (.I(I1580), .ZN(W790));
  INVX1 G37306 (.I(W2575), .ZN(O18906));
  INVX1 G37307 (.I(I1740), .ZN(W870));
  INVX1 G37308 (.I(W10991), .ZN(O18903));
  INVX1 G37309 (.I(I1744), .ZN(W872));
  INVX1 G37310 (.I(W8781), .ZN(O18901));
  INVX1 G37311 (.I(W32404), .ZN(O18899));
  INVX1 G37312 (.I(I1756), .ZN(W878));
  INVX1 G37313 (.I(W29131), .ZN(O18895));
  INVX1 G37314 (.I(I1432), .ZN(W716));
  INVX1 G37315 (.I(W28630), .ZN(O19063));
  INVX1 G37316 (.I(I1416), .ZN(W708));
  INVX1 G37317 (.I(W24975), .ZN(O19061));
  INVX1 G37318 (.I(W44996), .ZN(O19060));
  INVX1 G37319 (.I(W41788), .ZN(O19059));
  INVX1 G37320 (.I(W4011), .ZN(O19058));
  INVX1 G37321 (.I(W28962), .ZN(O19056));
  INVX1 G37322 (.I(W2592), .ZN(O19054));
  INVX1 G37323 (.I(W19791), .ZN(O19053));
  INVX1 G37324 (.I(W8672), .ZN(O19064));
  INVX1 G37325 (.I(W41187), .ZN(O19049));
  INVX1 G37326 (.I(W28037), .ZN(O19047));
  INVX1 G37327 (.I(I1442), .ZN(W721));
  INVX1 G37328 (.I(W5368), .ZN(O19044));
  INVX1 G37329 (.I(W23781), .ZN(O19043));
  INVX1 G37330 (.I(W8809), .ZN(O19042));
  INVX1 G37331 (.I(I1450), .ZN(W725));
  INVX1 G37332 (.I(W27655), .ZN(O19037));
  INVX1 G37333 (.I(I624), .ZN(O19075));
  INVX1 G37334 (.I(W3788), .ZN(O19087));
  INVX1 G37335 (.I(W4966), .ZN(O19086));
  INVX1 G37336 (.I(I1382), .ZN(W691));
  INVX1 G37337 (.I(W39605), .ZN(O19084));
  INVX1 G37338 (.I(W3907), .ZN(O19083));
  INVX1 G37339 (.I(W8701), .ZN(O19082));
  INVX1 G37340 (.I(W24108), .ZN(O19080));
  INVX1 G37341 (.I(I1386), .ZN(W693));
  INVX1 G37342 (.I(W15936), .ZN(O19077));
  INVX1 G37343 (.I(I1468), .ZN(W734));
  INVX1 G37344 (.I(W47877), .ZN(O19074));
  INVX1 G37345 (.I(W46739), .ZN(O19073));
  INVX1 G37346 (.I(W36022), .ZN(O19072));
  INVX1 G37347 (.I(I1396), .ZN(W698));
  INVX1 G37348 (.I(I1404), .ZN(W702));
  INVX1 G37349 (.I(W9644), .ZN(O19069));
  INVX1 G37350 (.I(W46317), .ZN(O19066));
  INVX1 G37351 (.I(I1412), .ZN(W706));
  INVX1 G37352 (.I(I1542), .ZN(W771));
  INVX1 G37353 (.I(I1520), .ZN(W760));
  INVX1 G37354 (.I(I1524), .ZN(W762));
  INVX1 G37355 (.I(I1526), .ZN(W763));
  INVX1 G37356 (.I(W27911), .ZN(O19002));
  INVX1 G37357 (.I(W29275), .ZN(O19001));
  INVX1 G37358 (.I(I563), .ZN(O18999));
  INVX1 G37359 (.I(W42602), .ZN(O18997));
  INVX1 G37360 (.I(I1536), .ZN(W768));
  INVX1 G37361 (.I(I1538), .ZN(W769));
  INVX1 G37362 (.I(W2214), .ZN(O19007));
  INVX1 G37363 (.I(I1548), .ZN(W774));
  INVX1 G37364 (.I(W31417), .ZN(O18991));
  INVX1 G37365 (.I(I1550), .ZN(W775));
  INVX1 G37366 (.I(I1554), .ZN(W777));
  INVX1 G37367 (.I(W5380), .ZN(O18987));
  INVX1 G37368 (.I(I1558), .ZN(W779));
  INVX1 G37369 (.I(W29), .ZN(O18985));
  INVX1 G37370 (.I(I1566), .ZN(W783));
  INVX1 G37371 (.I(I1486), .ZN(W743));
  INVX1 G37372 (.I(I522), .ZN(O19034));
  INVX1 G37373 (.I(W28447), .ZN(O19031));
  INVX1 G37374 (.I(I1478), .ZN(W739));
  INVX1 G37375 (.I(I1480), .ZN(W740));
  INVX1 G37376 (.I(W44041), .ZN(O19027));
  INVX1 G37377 (.I(W14604), .ZN(O19026));
  INVX1 G37378 (.I(W43030), .ZN(O19025));
  INVX1 G37379 (.I(I1484), .ZN(W742));
  INVX1 G37380 (.I(W6185), .ZN(O19334));
  INVX1 G37381 (.I(I1498), .ZN(W749));
  INVX1 G37382 (.I(W33505), .ZN(O19017));
  INVX1 G37383 (.I(I1510), .ZN(W755));
  INVX1 G37384 (.I(W50198), .ZN(O19013));
  INVX1 G37385 (.I(I1514), .ZN(W757));
  INVX1 G37386 (.I(W46886), .ZN(O19011));
  INVX1 G37387 (.I(W33742), .ZN(O19010));
  INVX1 G37388 (.I(I1516), .ZN(W758));
  INVX1 G37389 (.I(I278), .ZN(W139));
  INVX1 G37390 (.I(W26289), .ZN(O19635));
  INVX1 G37391 (.I(I250), .ZN(W125));
  INVX1 G37392 (.I(I264), .ZN(W132));
  INVX1 G37393 (.I(W44034), .ZN(O19629));
  INVX1 G37394 (.I(W4762), .ZN(O19628));
  INVX1 G37395 (.I(W28200), .ZN(O19627));
  INVX1 G37396 (.I(W9663), .ZN(O19626));
  INVX1 G37397 (.I(I272), .ZN(W136));
  INVX1 G37398 (.I(I274), .ZN(W137));
  INVX1 G37399 (.I(W11885), .ZN(O19638));
  INVX1 G37400 (.I(W44263), .ZN(O19620));
  INVX1 G37401 (.I(W21320), .ZN(O19619));
  INVX1 G37402 (.I(I280), .ZN(W140));
  INVX1 G37403 (.I(I286), .ZN(W143));
  INVX1 G37404 (.I(W39036), .ZN(O19615));
  INVX1 G37405 (.I(W6304), .ZN(O19612));
  INVX1 G37406 (.I(I292), .ZN(O0));
  INVX1 G37407 (.I(W3716), .ZN(O19610));
  INVX1 G37408 (.I(I182), .ZN(W91));
  INVX1 G37409 (.I(I158), .ZN(W79));
  INVX1 G37410 (.I(W13138), .ZN(O19668));
  INVX1 G37411 (.I(I166), .ZN(W83));
  INVX1 G37412 (.I(W28183), .ZN(O19665));
  INVX1 G37413 (.I(I172), .ZN(W86));
  INVX1 G37414 (.I(W14019), .ZN(O19663));
  INVX1 G37415 (.I(W16624), .ZN(O19662));
  INVX1 G37416 (.I(I176), .ZN(W88));
  INVX1 G37417 (.I(W14614), .ZN(O19660));
  INVX1 G37418 (.I(I294), .ZN(W147));
  INVX1 G37419 (.I(I186), .ZN(W93));
  INVX1 G37420 (.I(I188), .ZN(W94));
  INVX1 G37421 (.I(W34567), .ZN(O19656));
  INVX1 G37422 (.I(I198), .ZN(W99));
  INVX1 G37423 (.I(I200), .ZN(W100));
  INVX1 G37424 (.I(I204), .ZN(W102));
  INVX1 G37425 (.I(I210), .ZN(W105));
  INVX1 G37426 (.I(W21252), .ZN(O19644));
  INVX1 G37427 (.I(W14502), .ZN(O19563));
  INVX1 G37428 (.I(I366), .ZN(O1));
  INVX1 G37429 (.I(W38869), .ZN(O19572));
  INVX1 G37430 (.I(W9511), .ZN(O19571));
  INVX1 G37431 (.I(I368), .ZN(W184));
  INVX1 G37432 (.I(I372), .ZN(W186));
  INVX1 G37433 (.I(W17832), .ZN(O19567));
  INVX1 G37434 (.I(I376), .ZN(W188));
  INVX1 G37435 (.I(I378), .ZN(W189));
  INVX1 G37436 (.I(I380), .ZN(W190));
  INVX1 G37437 (.I(W14432), .ZN(O19574));
  INVX1 G37438 (.I(I382), .ZN(W191));
  INVX1 G37439 (.I(W3485), .ZN(O19558));
  INVX1 G37440 (.I(W11341), .ZN(O19557));
  INVX1 G37441 (.I(I394), .ZN(W197));
  INVX1 G37442 (.I(I396), .ZN(W198));
  INVX1 G37443 (.I(I398), .ZN(W199));
  INVX1 G37444 (.I(I402), .ZN(W201));
  INVX1 G37445 (.I(W17483), .ZN(O19551));
  INVX1 G37446 (.I(W24167), .ZN(O19589));
  INVX1 G37447 (.I(I306), .ZN(W153));
  INVX1 G37448 (.I(W20999), .ZN(O19602));
  INVX1 G37449 (.I(I310), .ZN(W155));
  INVX1 G37450 (.I(W43394), .ZN(O19599));
  INVX1 G37451 (.I(I320), .ZN(W160));
  INVX1 G37452 (.I(I324), .ZN(W162));
  INVX1 G37453 (.I(I326), .ZN(W163));
  INVX1 G37454 (.I(I332), .ZN(W166));
  INVX1 G37455 (.I(W48558), .ZN(W50909));
  INVX1 G37456 (.I(I340), .ZN(W170));
  INVX1 G37457 (.I(I342), .ZN(W171));
  INVX1 G37458 (.I(I344), .ZN(W172));
  INVX1 G37459 (.I(W43710), .ZN(O19584));
  INVX1 G37460 (.I(W28049), .ZN(O19583));
  INVX1 G37461 (.I(W47531), .ZN(O19579));
  INVX1 G37462 (.I(I358), .ZN(W179));
  INVX1 G37463 (.I(I362), .ZN(W181));
  INVX1 G37464 (.I(I68), .ZN(W34));
  INVX1 G37465 (.I(W5563), .ZN(O19735));
  INVX1 G37466 (.I(I52), .ZN(W26));
  INVX1 G37467 (.I(W26252), .ZN(O19733));
  INVX1 G37468 (.I(I58), .ZN(W29));
  INVX1 G37469 (.I(W50437), .ZN(O19729));
  INVX1 G37470 (.I(W43986), .ZN(O19728));
  INVX1 G37471 (.I(I62), .ZN(W31));
  INVX1 G37472 (.I(I66), .ZN(W33));
  INVX1 G37473 (.I(W31250), .ZN(O19725));
  INVX1 G37474 (.I(W37110), .ZN(O19736));
  INVX1 G37475 (.I(W33348), .ZN(O19723));
  INVX1 G37476 (.I(I72), .ZN(W36));
  INVX1 G37477 (.I(I76), .ZN(W38));
  INVX1 G37478 (.I(W14651), .ZN(O19720));
  INVX1 G37479 (.I(I82), .ZN(W41));
  INVX1 G37480 (.I(W21781), .ZN(O19718));
  INVX1 G37481 (.I(I86), .ZN(W43));
  INVX1 G37482 (.I(W27368), .ZN(O19715));
  INVX1 G37483 (.I(W3856), .ZN(O19747));
  INVX1 G37484 (.I(W23040), .ZN(O19762));
  INVX1 G37485 (.I(W5), .ZN(O19761));
  INVX1 G37486 (.I(I0), .ZN(W0));
  INVX1 G37487 (.I(I14), .ZN(W7));
  INVX1 G37488 (.I(W46110), .ZN(O19756));
  INVX1 G37489 (.I(W4232), .ZN(O19755));
  INVX1 G37490 (.I(I24), .ZN(W12));
  INVX1 G37491 (.I(W17198), .ZN(O19750));
  INVX1 G37492 (.I(W15785), .ZN(O19749));
  INVX1 G37493 (.I(I88), .ZN(W44));
  INVX1 G37494 (.I(W7112), .ZN(O19746));
  INVX1 G37495 (.I(I32), .ZN(W16));
  INVX1 G37496 (.I(I34), .ZN(W17));
  INVX1 G37497 (.I(I36), .ZN(W18));
  INVX1 G37498 (.I(W27949), .ZN(O19742));
  INVX1 G37499 (.I(I40), .ZN(W20));
  INVX1 G37500 (.I(W35880), .ZN(O19738));
  INVX1 G37501 (.I(I46), .ZN(W23));
  INVX1 G37502 (.I(W8643), .ZN(O19680));
  INVX1 G37503 (.I(W2286), .ZN(O19691));
  INVX1 G37504 (.I(I124), .ZN(W62));
  INVX1 G37505 (.I(W9374), .ZN(O19689));
  INVX1 G37506 (.I(I126), .ZN(W63));
  INVX1 G37507 (.I(W41387), .ZN(O19687));
  INVX1 G37508 (.I(I128), .ZN(W64));
  INVX1 G37509 (.I(I130), .ZN(W65));
  INVX1 G37510 (.I(W991), .ZN(O19684));
  INVX1 G37511 (.I(I132), .ZN(W66));
  INVX1 G37512 (.I(W25355), .ZN(O19692));
  INVX1 G37513 (.I(W38006), .ZN(O19679));
  INVX1 G37514 (.I(W34598), .ZN(O19678));
  INVX1 G37515 (.I(I138), .ZN(W69));
  INVX1 G37516 (.I(I140), .ZN(W70));
  INVX1 G37517 (.I(I142), .ZN(W71));
  INVX1 G37518 (.I(I148), .ZN(W74));
  INVX1 G37519 (.I(I154), .ZN(W77));
  INVX1 G37520 (.I(W31911), .ZN(O19671));
  INVX1 G37521 (.I(I106), .ZN(W53));
  INVX1 G37522 (.I(I92), .ZN(W46));
  INVX1 G37523 (.I(I96), .ZN(W48));
  INVX1 G37524 (.I(I98), .ZN(W49));
  INVX1 G37525 (.I(I100), .ZN(W50));
  INVX1 G37526 (.I(W10074), .ZN(O19708));
  INVX1 G37527 (.I(W25119), .ZN(O19707));
  INVX1 G37528 (.I(W28674), .ZN(O19706));
  INVX1 G37529 (.I(I104), .ZN(W52));
  INVX1 G37530 (.I(I410), .ZN(W205));
  INVX1 G37531 (.I(W31608), .ZN(O19702));
  INVX1 G37532 (.I(W32653), .ZN(O19700));
  INVX1 G37533 (.I(W49362), .ZN(O19699));
  INVX1 G37534 (.I(I118), .ZN(W59));
  INVX1 G37535 (.I(W15209), .ZN(O19696));
  INVX1 G37536 (.I(W46037), .ZN(O19695));
  INVX1 G37537 (.I(W36774), .ZN(O19694));
  INVX1 G37538 (.I(W39466), .ZN(O19693));
  INVX1 G37539 (.I(I748), .ZN(W374));
  INVX1 G37540 (.I(W11830), .ZN(O19406));
  INVX1 G37541 (.I(I732), .ZN(W366));
  INVX1 G37542 (.I(I738), .ZN(W369));
  INVX1 G37543 (.I(W37465), .ZN(O19401));
  INVX1 G37544 (.I(W33042), .ZN(O19398));
  INVX1 G37545 (.I(W10820), .ZN(O19397));
  INVX1 G37546 (.I(W49893), .ZN(O19395));
  INVX1 G37547 (.I(W39065), .ZN(O19394));
  INVX1 G37548 (.I(W39454), .ZN(O19393));
  INVX1 G37549 (.I(I716), .ZN(W358));
  INVX1 G37550 (.I(W23296), .ZN(O19391));
  INVX1 G37551 (.I(W36239), .ZN(W50627));
  INVX1 G37552 (.I(I750), .ZN(W375));
  INVX1 G37553 (.I(I756), .ZN(W378));
  INVX1 G37554 (.I(W40307), .ZN(O19387));
  INVX1 G37555 (.I(W33762), .ZN(O19386));
  INVX1 G37556 (.I(W47952), .ZN(O19384));
  INVX1 G37557 (.I(I760), .ZN(W380));
  INVX1 G37558 (.I(W29104), .ZN(O19422));
  INVX1 G37559 (.I(W15195), .ZN(O19437));
  INVX1 G37560 (.I(I650), .ZN(W325));
  INVX1 G37561 (.I(I652), .ZN(W326));
  INVX1 G37562 (.I(W22327), .ZN(O19432));
  INVX1 G37563 (.I(W29547), .ZN(O19431));
  INVX1 G37564 (.I(I662), .ZN(W331));
  INVX1 G37565 (.I(W50), .ZN(O19427));
  INVX1 G37566 (.I(I666), .ZN(W333));
  INVX1 G37567 (.I(W40550), .ZN(O19425));
  INVX1 G37568 (.I(I762), .ZN(W381));
  INVX1 G37569 (.I(I688), .ZN(W344));
  INVX1 G37570 (.I(W6540), .ZN(O19417));
  INVX1 G37571 (.I(I698), .ZN(W349));
  INVX1 G37572 (.I(W29996), .ZN(O19415));
  INVX1 G37573 (.I(I702), .ZN(W351));
  INVX1 G37574 (.I(I708), .ZN(W354));
  INVX1 G37575 (.I(W50105), .ZN(O19410));
  INVX1 G37576 (.I(W34304), .ZN(O19409));
  INVX1 G37577 (.I(W40649), .ZN(O19344));
  INVX1 G37578 (.I(I804), .ZN(W402));
  INVX1 G37579 (.I(I806), .ZN(W403));
  INVX1 G37580 (.I(W36972), .ZN(O19355));
  INVX1 G37581 (.I(I822), .ZN(W411));
  INVX1 G37582 (.I(W46164), .ZN(O19352));
  INVX1 G37583 (.I(I834), .ZN(W417));
  INVX1 G37584 (.I(I836), .ZN(W418));
  INVX1 G37585 (.I(I840), .ZN(W420));
  INVX1 G37586 (.I(W47185), .ZN(O19345));
  INVX1 G37587 (.I(W24000), .ZN(O19360));
  INVX1 G37588 (.I(I844), .ZN(W422));
  INVX1 G37589 (.I(I846), .ZN(W423));
  INVX1 G37590 (.I(W14259), .ZN(O19340));
  INVX1 G37591 (.I(I850), .ZN(W425));
  INVX1 G37592 (.I(I854), .ZN(W427));
  INVX1 G37593 (.I(I864), .ZN(W432));
  INVX1 G37594 (.I(W14998), .ZN(O19336));
  INVX1 G37595 (.I(I866), .ZN(W433));
  INVX1 G37596 (.I(I794), .ZN(W397));
  INVX1 G37597 (.I(W11532), .ZN(O19381));
  INVX1 G37598 (.I(I768), .ZN(W384));
  INVX1 G37599 (.I(I774), .ZN(W387));
  INVX1 G37600 (.I(W32751), .ZN(O19376));
  INVX1 G37601 (.I(W47824), .ZN(O19375));
  INVX1 G37602 (.I(I782), .ZN(W391));
  INVX1 G37603 (.I(W517), .ZN(O19373));
  INVX1 G37604 (.I(I788), .ZN(W394));
  INVX1 G37605 (.I(I644), .ZN(W322));
  INVX1 G37606 (.I(W39376), .ZN(O19370));
  INVX1 G37607 (.I(W47195), .ZN(O19369));
  INVX1 G37608 (.I(W13712), .ZN(O19366));
  INVX1 G37609 (.I(I800), .ZN(W400));
  INVX1 G37610 (.I(W6225), .ZN(O19364));
  INVX1 G37611 (.I(I802), .ZN(W401));
  INVX1 G37612 (.I(W44457), .ZN(O19362));
  INVX1 G37613 (.I(W2934), .ZN(O19361));
  INVX1 G37614 (.I(I496), .ZN(W248));
  INVX1 G37615 (.I(I472), .ZN(W236));
  INVX1 G37616 (.I(W36884), .ZN(O19518));
  INVX1 G37617 (.I(W16076), .ZN(O19517));
  INVX1 G37618 (.I(W33929), .ZN(O19515));
  INVX1 G37619 (.I(W1010), .ZN(O19514));
  INVX1 G37620 (.I(W8529), .ZN(O19513));
  INVX1 G37621 (.I(W46754), .ZN(O19510));
  INVX1 G37622 (.I(I486), .ZN(W243));
  INVX1 G37623 (.I(W37149), .ZN(O19507));
  INVX1 G37624 (.I(I464), .ZN(W232));
  INVX1 G37625 (.I(W33846), .ZN(O19502));
  INVX1 G37626 (.I(W35150), .ZN(O19499));
  INVX1 G37627 (.I(W14740), .ZN(O19496));
  INVX1 G37628 (.I(I512), .ZN(W256));
  INVX1 G37629 (.I(I514), .ZN(W257));
  INVX1 G37630 (.I(W4385), .ZN(O19493));
  INVX1 G37631 (.I(I522), .ZN(W261));
  INVX1 G37632 (.I(W32306), .ZN(O19491));
  INVX1 G37633 (.I(I448), .ZN(W224));
  INVX1 G37634 (.I(I418), .ZN(W209));
  INVX1 G37635 (.I(I798), .ZN(O19546));
  INVX1 G37636 (.I(I424), .ZN(W212));
  INVX1 G37637 (.I(W44018), .ZN(O19543));
  INVX1 G37638 (.I(I426), .ZN(W213));
  INVX1 G37639 (.I(W30036), .ZN(O19541));
  INVX1 G37640 (.I(W6912), .ZN(O19539));
  INVX1 G37641 (.I(W14715), .ZN(O19536));
  INVX1 G37642 (.I(W45544), .ZN(O19534));
  INVX1 G37643 (.I(I528), .ZN(W264));
  INVX1 G37644 (.I(W11192), .ZN(O19531));
  INVX1 G37645 (.I(W20702), .ZN(O19530));
  INVX1 G37646 (.I(I452), .ZN(W226));
  INVX1 G37647 (.I(W13169), .ZN(O19528));
  INVX1 G37648 (.I(W18279), .ZN(O19527));
  INVX1 G37649 (.I(I460), .ZN(W230));
  INVX1 G37650 (.I(W19881), .ZN(O19524));
  INVX1 G37651 (.I(W41127), .ZN(O19523));
  INVX1 G37652 (.I(I610), .ZN(W305));
  INVX1 G37653 (.I(W49756), .ZN(O19463));
  INVX1 G37654 (.I(I404), .ZN(O19462));
  INVX1 G37655 (.I(W23359), .ZN(O19461));
  INVX1 G37656 (.I(W48708), .ZN(W50698));
  INVX1 G37657 (.I(W35114), .ZN(O19459));
  INVX1 G37658 (.I(I598), .ZN(W299));
  INVX1 G37659 (.I(W13512), .ZN(O19455));
  INVX1 G37660 (.I(W47004), .ZN(O19454));
  INVX1 G37661 (.I(W38267), .ZN(O19453));
  INVX1 G37662 (.I(W28035), .ZN(O19464));
  INVX1 G37663 (.I(W8821), .ZN(O19448));
  INVX1 G37664 (.I(W8849), .ZN(O19447));
  INVX1 G37665 (.I(I616), .ZN(W308));
  INVX1 G37666 (.I(W33634), .ZN(O19445));
  INVX1 G37667 (.I(I626), .ZN(W313));
  INVX1 G37668 (.I(I398), .ZN(O19442));
  INVX1 G37669 (.I(W21491), .ZN(O19441));
  INVX1 G37670 (.I(W41517), .ZN(O19440));
  INVX1 G37671 (.I(W29812), .ZN(O19475));
  INVX1 G37672 (.I(I544), .ZN(W272));
  INVX1 G37673 (.I(I552), .ZN(W276));
  INVX1 G37674 (.I(I560), .ZN(W280));
  INVX1 G37675 (.I(W7341), .ZN(O19482));
  INVX1 G37676 (.I(I568), .ZN(W284));
  INVX1 G37677 (.I(I570), .ZN(W285));
  INVX1 G37678 (.I(I572), .ZN(W286));
  INVX1 G37679 (.I(W32377), .ZN(O19476));
  INVX1 G37680 (.I(I1822), .ZN(W911));
  INVX1 G37681 (.I(W1685), .ZN(O19474));
  INVX1 G37682 (.I(I576), .ZN(W288));
  INVX1 G37683 (.I(I584), .ZN(W292));
  INVX1 G37684 (.I(I588), .ZN(W294));
  INVX1 G37685 (.I(I590), .ZN(W295));
  INVX1 G37686 (.I(W42864), .ZN(O19467));
  INVX1 G37687 (.I(W45625), .ZN(O19466));
  INVX1 G37688 (.I(I592), .ZN(W296));
  INVX1 G37689 (.I(I268), .ZN(O18306));
  INVX1 G37690 (.I(I1898), .ZN(W1490));
  INVX1 G37691 (.I(W13754), .ZN(O18318));
  INVX1 G37692 (.I(W6038), .ZN(O18317));
  INVX1 G37693 (.I(W39050), .ZN(O18316));
  INVX1 G37694 (.I(W30797), .ZN(O18315));
  INVX1 G37695 (.I(I1604), .ZN(W1491));
  INVX1 G37696 (.I(I262), .ZN(W1494));
  INVX1 G37697 (.I(W2033), .ZN(O18311));
  INVX1 G37698 (.I(W500), .ZN(O14));
  INVX1 G37699 (.I(W607), .ZN(W1489));
  INVX1 G37700 (.I(I1188), .ZN(W1505));
  INVX1 G37701 (.I(I1636), .ZN(W1506));
  INVX1 G37702 (.I(W36702), .ZN(O18302));
  INVX1 G37703 (.I(W16300), .ZN(O18300));
  INVX1 G37704 (.I(I1322), .ZN(W1509));
  INVX1 G37705 (.I(I120), .ZN(W1510));
  INVX1 G37706 (.I(W22624), .ZN(O18297));
  INVX1 G37707 (.I(W24302), .ZN(O18296));
  INVX1 G37708 (.I(W23179), .ZN(O18333));
  INVX1 G37709 (.I(W33699), .ZN(O18345));
  INVX1 G37710 (.I(W21530), .ZN(O18344));
  INVX1 G37711 (.I(W42254), .ZN(O18343));
  INVX1 G37712 (.I(I1029), .ZN(W1464));
  INVX1 G37713 (.I(I435), .ZN(W1467));
  INVX1 G37714 (.I(W22505), .ZN(O18337));
  INVX1 G37715 (.I(W1414), .ZN(W1471));
  INVX1 G37716 (.I(I1697), .ZN(W1473));
  INVX1 G37717 (.I(I1153), .ZN(W1475));
  INVX1 G37718 (.I(W577), .ZN(W1511));
  INVX1 G37719 (.I(W44904), .ZN(O18330));
  INVX1 G37720 (.I(W28750), .ZN(W49528));
  INVX1 G37721 (.I(I621), .ZN(W1479));
  INVX1 G37722 (.I(W39635), .ZN(O18329));
  INVX1 G37723 (.I(W31587), .ZN(O18328));
  INVX1 G37724 (.I(I644), .ZN(W1481));
  INVX1 G37725 (.I(I930), .ZN(W1482));
  INVX1 G37726 (.I(W6924), .ZN(O18322));
  INVX1 G37727 (.I(W41270), .ZN(O18256));
  INVX1 G37728 (.I(W1425), .ZN(W1533));
  INVX1 G37729 (.I(W25992), .ZN(O18267));
  INVX1 G37730 (.I(W13264), .ZN(O18266));
  INVX1 G37731 (.I(I1338), .ZN(W1538));
  INVX1 G37732 (.I(W27296), .ZN(O18264));
  INVX1 G37733 (.I(W26044), .ZN(O18261));
  INVX1 G37734 (.I(I740), .ZN(W1542));
  INVX1 G37735 (.I(W23687), .ZN(O18259));
  INVX1 G37736 (.I(W555), .ZN(W1544));
  INVX1 G37737 (.I(W654), .ZN(W1530));
  INVX1 G37738 (.I(I887), .ZN(W1545));
  INVX1 G37739 (.I(I185), .ZN(W1546));
  INVX1 G37740 (.I(W241), .ZN(W1550));
  INVX1 G37741 (.I(I1760), .ZN(O18252));
  INVX1 G37742 (.I(W4977), .ZN(O18251));
  INVX1 G37743 (.I(W664), .ZN(W1551));
  INVX1 G37744 (.I(W29264), .ZN(O18249));
  INVX1 G37745 (.I(W46415), .ZN(O18246));
  INVX1 G37746 (.I(W47649), .ZN(O18285));
  INVX1 G37747 (.I(W12328), .ZN(O18294));
  INVX1 G37748 (.I(I975), .ZN(W1512));
  INVX1 G37749 (.I(W1215), .ZN(W1513));
  INVX1 G37750 (.I(I315), .ZN(W1514));
  INVX1 G37751 (.I(W3321), .ZN(O18290));
  INVX1 G37752 (.I(W21113), .ZN(O18289));
  INVX1 G37753 (.I(I1066), .ZN(W1516));
  INVX1 G37754 (.I(I1889), .ZN(W1517));
  INVX1 G37755 (.I(W39322), .ZN(O18346));
  INVX1 G37756 (.I(I356), .ZN(W1521));
  INVX1 G37757 (.I(W14256), .ZN(O18280));
  INVX1 G37758 (.I(I459), .ZN(W1522));
  INVX1 G37759 (.I(I1214), .ZN(W1524));
  INVX1 G37760 (.I(W10360), .ZN(O18277));
  INVX1 G37761 (.I(I424), .ZN(W1526));
  INVX1 G37762 (.I(W20012), .ZN(O18274));
  INVX1 G37763 (.I(W1418), .ZN(W1528));
  INVX1 G37764 (.I(I1577), .ZN(W1401));
  INVX1 G37765 (.I(W4241), .ZN(O18419));
  INVX1 G37766 (.I(W940), .ZN(W1388));
  INVX1 G37767 (.I(W632), .ZN(W1390));
  INVX1 G37768 (.I(W102), .ZN(W1391));
  INVX1 G37769 (.I(W711), .ZN(W1392));
  INVX1 G37770 (.I(I970), .ZN(W1398));
  INVX1 G37771 (.I(W15968), .ZN(W49615));
  INVX1 G37772 (.I(W22254), .ZN(O18412));
  INVX1 G37773 (.I(W30910), .ZN(O18410));
  INVX1 G37774 (.I(W40904), .ZN(O18420));
  INVX1 G37775 (.I(W1493), .ZN(O18408));
  INVX1 G37776 (.I(W2904), .ZN(O18406));
  INVX1 G37777 (.I(W616), .ZN(W1403));
  INVX1 G37778 (.I(I1122), .ZN(W1405));
  INVX1 G37779 (.I(W48350), .ZN(O18401));
  INVX1 G37780 (.I(W44004), .ZN(O18400));
  INVX1 G37781 (.I(I1717), .ZN(W1411));
  INVX1 G37782 (.I(W32387), .ZN(O18397));
  INVX1 G37783 (.I(I1508), .ZN(W1384));
  INVX1 G37784 (.I(W723), .ZN(W1373));
  INVX1 G37785 (.I(W47458), .ZN(O18438));
  INVX1 G37786 (.I(W30975), .ZN(O18437));
  INVX1 G37787 (.I(W27829), .ZN(O18436));
  INVX1 G37788 (.I(I1544), .ZN(W1374));
  INVX1 G37789 (.I(I698), .ZN(W1376));
  INVX1 G37790 (.I(W20599), .ZN(O18432));
  INVX1 G37791 (.I(I1856), .ZN(W1379));
  INVX1 G37792 (.I(I1506), .ZN(W1383));
  INVX1 G37793 (.I(I1755), .ZN(O18396));
  INVX1 G37794 (.I(W838), .ZN(W1385));
  INVX1 G37795 (.I(W43482), .ZN(O18427));
  INVX1 G37796 (.I(I1103), .ZN(W1386));
  INVX1 G37797 (.I(W38323), .ZN(O18425));
  INVX1 G37798 (.I(W22470), .ZN(O18423));
  INVX1 G37799 (.I(W23959), .ZN(O18422));
  INVX1 G37800 (.I(W42769), .ZN(O18421));
  INVX1 G37801 (.I(W31913), .ZN(W49624));
  INVX1 G37802 (.I(I418), .ZN(W1451));
  INVX1 G37803 (.I(W1669), .ZN(O18368));
  INVX1 G37804 (.I(W176), .ZN(W1443));
  INVX1 G37805 (.I(I1088), .ZN(W1444));
  INVX1 G37806 (.I(W43232), .ZN(O18364));
  INVX1 G37807 (.I(W41193), .ZN(O18363));
  INVX1 G37808 (.I(I1597), .ZN(W1445));
  INVX1 G37809 (.I(W42354), .ZN(O18361));
  INVX1 G37810 (.I(W1129), .ZN(O13));
  INVX1 G37811 (.I(I444), .ZN(W1448));
  INVX1 G37812 (.I(W41582), .ZN(O18370));
  INVX1 G37813 (.I(I1976), .ZN(W1454));
  INVX1 G37814 (.I(W12925), .ZN(O18355));
  INVX1 G37815 (.I(W38512), .ZN(O18354));
  INVX1 G37816 (.I(I450), .ZN(W1459));
  INVX1 G37817 (.I(W46544), .ZN(O18350));
  INVX1 G37818 (.I(W18216), .ZN(W49549));
  INVX1 G37819 (.I(I405), .ZN(W1462));
  INVX1 G37820 (.I(W16704), .ZN(O18347));
  INVX1 G37821 (.I(W52), .ZN(W1423));
  INVX1 G37822 (.I(W33137), .ZN(O18395));
  INVX1 G37823 (.I(W21158), .ZN(O18393));
  INVX1 G37824 (.I(W447), .ZN(W1414));
  INVX1 G37825 (.I(I229), .ZN(W1419));
  INVX1 G37826 (.I(W1101), .ZN(W1420));
  INVX1 G37827 (.I(W3248), .ZN(O18387));
  INVX1 G37828 (.I(W46377), .ZN(O18386));
  INVX1 G37829 (.I(W57), .ZN(W1422));
  INVX1 G37830 (.I(W709), .ZN(O18243));
  INVX1 G37831 (.I(W17311), .ZN(O18383));
  INVX1 G37832 (.I(W29154), .ZN(O18382));
  INVX1 G37833 (.I(I1621), .ZN(W1424));
  INVX1 G37834 (.I(W47), .ZN(W1428));
  INVX1 G37835 (.I(I1168), .ZN(W1431));
  INVX1 G37836 (.I(W1158), .ZN(W1432));
  INVX1 G37837 (.I(W15047), .ZN(O18375));
  INVX1 G37838 (.I(W45641), .ZN(O18372));
  INVX1 G37839 (.I(W10064), .ZN(O18108));
  INVX1 G37840 (.I(W24807), .ZN(O18119));
  INVX1 G37841 (.I(I572), .ZN(W1696));
  INVX1 G37842 (.I(W4459), .ZN(O18117));
  INVX1 G37843 (.I(I1596), .ZN(W1697));
  INVX1 G37844 (.I(W531), .ZN(W1698));
  INVX1 G37845 (.I(W37533), .ZN(O18113));
  INVX1 G37846 (.I(W18435), .ZN(O18112));
  INVX1 G37847 (.I(W92), .ZN(W1704));
  INVX1 G37848 (.I(W26048), .ZN(O18109));
  INVX1 G37849 (.I(W662), .ZN(W1695));
  INVX1 G37850 (.I(W34075), .ZN(O18107));
  INVX1 G37851 (.I(W13941), .ZN(W49293));
  INVX1 G37852 (.I(W1224), .ZN(W1705));
  INVX1 G37853 (.I(I193), .ZN(W1707));
  INVX1 G37854 (.I(I1755), .ZN(W1709));
  INVX1 G37855 (.I(W1520), .ZN(W1710));
  INVX1 G37856 (.I(I331), .ZN(W1715));
  INVX1 G37857 (.I(W15667), .ZN(O18099));
  INVX1 G37858 (.I(W355), .ZN(W1676));
  INVX1 G37859 (.I(I1194), .ZN(W1660));
  INVX1 G37860 (.I(I524), .ZN(W1661));
  INVX1 G37861 (.I(W18922), .ZN(O18146));
  INVX1 G37862 (.I(W46), .ZN(W1670));
  INVX1 G37863 (.I(W27462), .ZN(O18139));
  INVX1 G37864 (.I(W1016), .ZN(W1672));
  INVX1 G37865 (.I(W27218), .ZN(O18137));
  INVX1 G37866 (.I(W9875), .ZN(O18136));
  INVX1 G37867 (.I(W15120), .ZN(O18135));
  INVX1 G37868 (.I(W16174), .ZN(O18098));
  INVX1 G37869 (.I(W14272), .ZN(O18133));
  INVX1 G37870 (.I(W302), .ZN(W1683));
  INVX1 G37871 (.I(W21313), .ZN(O18127));
  INVX1 G37872 (.I(I72), .ZN(W1686));
  INVX1 G37873 (.I(I1997), .ZN(W1687));
  INVX1 G37874 (.I(I1080), .ZN(W1689));
  INVX1 G37875 (.I(I236), .ZN(W1694));
  INVX1 G37876 (.I(W9314), .ZN(O18121));
  INVX1 G37877 (.I(W11721), .ZN(O18061));
  INVX1 G37878 (.I(W1338), .ZN(W1737));
  INVX1 G37879 (.I(I326), .ZN(W1739));
  INVX1 G37880 (.I(W43842), .ZN(O18070));
  INVX1 G37881 (.I(I1286), .ZN(W1747));
  INVX1 G37882 (.I(W42145), .ZN(O18068));
  INVX1 G37883 (.I(W17461), .ZN(O18067));
  INVX1 G37884 (.I(W2162), .ZN(O18066));
  INVX1 G37885 (.I(W46531), .ZN(O18064));
  INVX1 G37886 (.I(W15934), .ZN(O18063));
  INVX1 G37887 (.I(W268), .ZN(W1736));
  INVX1 G37888 (.I(W46361), .ZN(O18060));
  INVX1 G37889 (.I(W3422), .ZN(O18059));
  INVX1 G37890 (.I(W727), .ZN(W1750));
  INVX1 G37891 (.I(I1031), .ZN(W1755));
  INVX1 G37892 (.I(I1414), .ZN(W1756));
  INVX1 G37893 (.I(W1188), .ZN(W1764));
  INVX1 G37894 (.I(W25139), .ZN(O18050));
  INVX1 G37895 (.I(W1320), .ZN(W1766));
  INVX1 G37896 (.I(W790), .ZN(W1726));
  INVX1 G37897 (.I(I1126), .ZN(W1719));
  INVX1 G37898 (.I(I1147), .ZN(W1720));
  INVX1 G37899 (.I(W291), .ZN(W1721));
  INVX1 G37900 (.I(W17574), .ZN(O18093));
  INVX1 G37901 (.I(I1273), .ZN(W1722));
  INVX1 G37902 (.I(W1495), .ZN(O18091));
  INVX1 G37903 (.I(W1438), .ZN(W1723));
  INVX1 G37904 (.I(W10637), .ZN(O18089));
  INVX1 G37905 (.I(W5506), .ZN(O18149));
  INVX1 G37906 (.I(W37645), .ZN(O18087));
  INVX1 G37907 (.I(W45822), .ZN(O18086));
  INVX1 G37908 (.I(W2457), .ZN(O18085));
  INVX1 G37909 (.I(W1153), .ZN(W1728));
  INVX1 G37910 (.I(I43), .ZN(W1730));
  INVX1 G37911 (.I(W27229), .ZN(O18081));
  INVX1 G37912 (.I(W27542), .ZN(O18079));
  INVX1 G37913 (.I(I800), .ZN(W49262));
  INVX1 G37914 (.I(W21068), .ZN(O18209));
  INVX1 G37915 (.I(W1240), .ZN(W1583));
  INVX1 G37916 (.I(W1397), .ZN(W1584));
  INVX1 G37917 (.I(W2712), .ZN(O18218));
  INVX1 G37918 (.I(W37008), .ZN(O18217));
  INVX1 G37919 (.I(I1852), .ZN(W1587));
  INVX1 G37920 (.I(W1584), .ZN(W1588));
  INVX1 G37921 (.I(I1753), .ZN(W1590));
  INVX1 G37922 (.I(W14306), .ZN(O18211));
  INVX1 G37923 (.I(W1244), .ZN(W1592));
  INVX1 G37924 (.I(W792), .ZN(W1579));
  INVX1 G37925 (.I(W24433), .ZN(O18208));
  INVX1 G37926 (.I(W10737), .ZN(O18207));
  INVX1 G37927 (.I(W15126), .ZN(O18205));
  INVX1 G37928 (.I(W28521), .ZN(O18204));
  INVX1 G37929 (.I(I1696), .ZN(W1594));
  INVX1 G37930 (.I(W38843), .ZN(O18202));
  INVX1 G37931 (.I(I45), .ZN(W1595));
  INVX1 G37932 (.I(W7951), .ZN(O18200));
  INVX1 G37933 (.I(W36599), .ZN(O18233));
  INVX1 G37934 (.I(W1115), .ZN(W1558));
  INVX1 G37935 (.I(W10712), .ZN(O18242));
  INVX1 G37936 (.I(W1522), .ZN(W1561));
  INVX1 G37937 (.I(W1464), .ZN(W1563));
  INVX1 G37938 (.I(W42529), .ZN(O18239));
  INVX1 G37939 (.I(W2942), .ZN(O18237));
  INVX1 G37940 (.I(W36264), .ZN(O18236));
  INVX1 G37941 (.I(W40876), .ZN(O18234));
  INVX1 G37942 (.I(I654), .ZN(W1567));
  INVX1 G37943 (.I(I1118), .ZN(W1597));
  INVX1 G37944 (.I(I1611), .ZN(W1570));
  INVX1 G37945 (.I(I556), .ZN(W1572));
  INVX1 G37946 (.I(W519), .ZN(W1573));
  INVX1 G37947 (.I(W704), .ZN(W1574));
  INVX1 G37948 (.I(W814), .ZN(O18228));
  INVX1 G37949 (.I(I95), .ZN(W1575));
  INVX1 G37950 (.I(W14544), .ZN(O18226));
  INVX1 G37951 (.I(W1266), .ZN(W1576));
  INVX1 G37952 (.I(W6597), .ZN(O18162));
  INVX1 G37953 (.I(W34883), .ZN(W49362));
  INVX1 G37954 (.I(W954), .ZN(W1637));
  INVX1 G37955 (.I(W13569), .ZN(O18170));
  INVX1 G37956 (.I(I1506), .ZN(W1640));
  INVX1 G37957 (.I(W791), .ZN(W1644));
  INVX1 G37958 (.I(I20), .ZN(W1646));
  INVX1 G37959 (.I(W20872), .ZN(W49353));
  INVX1 G37960 (.I(W4371), .ZN(O18164));
  INVX1 G37961 (.I(W23850), .ZN(O18163));
  INVX1 G37962 (.I(W38267), .ZN(O18173));
  INVX1 G37963 (.I(W7328), .ZN(O18161));
  INVX1 G37964 (.I(W923), .ZN(W1647));
  INVX1 G37965 (.I(W1962), .ZN(O18158));
  INVX1 G37966 (.I(I1458), .ZN(W1653));
  INVX1 G37967 (.I(W1081), .ZN(W1654));
  INVX1 G37968 (.I(W118), .ZN(W1655));
  INVX1 G37969 (.I(W609), .ZN(W1656));
  INVX1 G37970 (.I(I1662), .ZN(W1657));
  INVX1 G37971 (.I(W3292), .ZN(O18184));
  INVX1 G37972 (.I(W28515), .ZN(O18196));
  INVX1 G37973 (.I(W113), .ZN(W1600));
  INVX1 G37974 (.I(I772), .ZN(W1604));
  INVX1 G37975 (.I(W28781), .ZN(O18192));
  INVX1 G37976 (.I(W814), .ZN(W1605));
  INVX1 G37977 (.I(W1230), .ZN(W1606));
  INVX1 G37978 (.I(I681), .ZN(W1611));
  INVX1 G37979 (.I(W11), .ZN(W1613));
  INVX1 G37980 (.I(I771), .ZN(W1371));
  INVX1 G37981 (.I(W33144), .ZN(O18183));
  INVX1 G37982 (.I(I1486), .ZN(W1616));
  INVX1 G37983 (.I(I289), .ZN(W1620));
  INVX1 G37984 (.I(W476), .ZN(W1625));
  INVX1 G37985 (.I(I1662), .ZN(W1626));
  INVX1 G37986 (.I(I1870), .ZN(W1627));
  INVX1 G37987 (.I(I637), .ZN(W1629));
  INVX1 G37988 (.I(W191), .ZN(W1631));
  INVX1 G37989 (.I(W18425), .ZN(O18718));
  INVX1 G37990 (.I(I247), .ZN(W1064));
  INVX1 G37991 (.I(I276), .ZN(O18728));
  INVX1 G37992 (.I(W20416), .ZN(O18725));
  INVX1 G37993 (.I(W12603), .ZN(W49942));
  INVX1 G37994 (.I(W602), .ZN(W1067));
  INVX1 G37995 (.I(W23205), .ZN(O18722));
  INVX1 G37996 (.I(I43), .ZN(W1069));
  INVX1 G37997 (.I(W39858), .ZN(O18720));
  INVX1 G37998 (.I(I619), .ZN(W1071));
  INVX1 G37999 (.I(W31015), .ZN(O18730));
  INVX1 G38000 (.I(W122), .ZN(W1072));
  INVX1 G38001 (.I(W11072), .ZN(O18715));
  INVX1 G38002 (.I(I1540), .ZN(W1076));
  INVX1 G38003 (.I(W686), .ZN(W1077));
  INVX1 G38004 (.I(W45811), .ZN(O18712));
  INVX1 G38005 (.I(I410), .ZN(W1078));
  INVX1 G38006 (.I(W19459), .ZN(O18710));
  INVX1 G38007 (.I(W34092), .ZN(O18709));
  INVX1 G38008 (.I(W21333), .ZN(O18742));
  INVX1 G38009 (.I(I1246), .ZN(W1040));
  INVX1 G38010 (.I(I1996), .ZN(W1042));
  INVX1 G38011 (.I(I1939), .ZN(W1043));
  INVX1 G38012 (.I(W12580), .ZN(O18753));
  INVX1 G38013 (.I(W421), .ZN(W1046));
  INVX1 G38014 (.I(W15575), .ZN(O18750));
  INVX1 G38015 (.I(W20493), .ZN(O18749));
  INVX1 G38016 (.I(W46621), .ZN(O18744));
  INVX1 G38017 (.I(I1476), .ZN(W1055));
  INVX1 G38018 (.I(W764), .ZN(W1080));
  INVX1 G38019 (.I(I1834), .ZN(W1057));
  INVX1 G38020 (.I(W29807), .ZN(O18739));
  INVX1 G38021 (.I(W27469), .ZN(O18738));
  INVX1 G38022 (.I(I1834), .ZN(W1058));
  INVX1 G38023 (.I(W40956), .ZN(O18736));
  INVX1 G38024 (.I(I1011), .ZN(W1062));
  INVX1 G38025 (.I(W49796), .ZN(O18733));
  INVX1 G38026 (.I(W46360), .ZN(O18732));
  INVX1 G38027 (.I(W42156), .ZN(O18669));
  INVX1 G38028 (.I(W35771), .ZN(O18684));
  INVX1 G38029 (.I(W41690), .ZN(O18682));
  INVX1 G38030 (.I(W17787), .ZN(O18680));
  INVX1 G38031 (.I(W717), .ZN(W1115));
  INVX1 G38032 (.I(W31181), .ZN(O18676));
  INVX1 G38033 (.I(I657), .ZN(W1122));
  INVX1 G38034 (.I(W928), .ZN(W1126));
  INVX1 G38035 (.I(I1969), .ZN(W1128));
  INVX1 G38036 (.I(W22812), .ZN(O18670));
  INVX1 G38037 (.I(W758), .ZN(W1106));
  INVX1 G38038 (.I(W11501), .ZN(O18665));
  INVX1 G38039 (.I(I1648), .ZN(W1134));
  INVX1 G38040 (.I(W28888), .ZN(O18663));
  INVX1 G38041 (.I(W159), .ZN(W1136));
  INVX1 G38042 (.I(I1666), .ZN(W1137));
  INVX1 G38043 (.I(W46686), .ZN(O18659));
  INVX1 G38044 (.I(I152), .ZN(W1141));
  INVX1 G38045 (.I(I704), .ZN(W1144));
  INVX1 G38046 (.I(I109), .ZN(W1092));
  INVX1 G38047 (.I(I1911), .ZN(W1081));
  INVX1 G38048 (.I(W153), .ZN(W1082));
  INVX1 G38049 (.I(I468), .ZN(W1084));
  INVX1 G38050 (.I(W44024), .ZN(O18703));
  INVX1 G38051 (.I(I1678), .ZN(W1086));
  INVX1 G38052 (.I(I1670), .ZN(W1087));
  INVX1 G38053 (.I(W21684), .ZN(O18699));
  INVX1 G38054 (.I(W9425), .ZN(O18698));
  INVX1 G38055 (.I(W7003), .ZN(O18758));
  INVX1 G38056 (.I(W43611), .ZN(O18696));
  INVX1 G38057 (.I(W3685), .ZN(O18695));
  INVX1 G38058 (.I(I933), .ZN(W1094));
  INVX1 G38059 (.I(W762), .ZN(W1095));
  INVX1 G38060 (.I(W16), .ZN(W1096));
  INVX1 G38061 (.I(W47968), .ZN(O18690));
  INVX1 G38062 (.I(I288), .ZN(W1100));
  INVX1 G38063 (.I(W27683), .ZN(O18687));
  INVX1 G38064 (.I(W29212), .ZN(O18826));
  INVX1 G38065 (.I(I1890), .ZN(W945));
  INVX1 G38066 (.I(I1896), .ZN(W948));
  INVX1 G38067 (.I(I1898), .ZN(W949));
  INVX1 G38068 (.I(I1904), .ZN(W952));
  INVX1 G38069 (.I(W17983), .ZN(O18832));
  INVX1 G38070 (.I(W34912), .ZN(O18831));
  INVX1 G38071 (.I(I1928), .ZN(W964));
  INVX1 G38072 (.I(W34562), .ZN(O18828));
  INVX1 G38073 (.I(W19763), .ZN(O18827));
  INVX1 G38074 (.I(I1884), .ZN(W942));
  INVX1 G38075 (.I(W16272), .ZN(O18825));
  INVX1 G38076 (.I(I1946), .ZN(W973));
  INVX1 G38077 (.I(W366), .ZN(O18819));
  INVX1 G38078 (.I(I1950), .ZN(W975));
  INVX1 G38079 (.I(I1960), .ZN(W980));
  INVX1 G38080 (.I(W10606), .ZN(O18813));
  INVX1 G38081 (.I(W13989), .ZN(O18811));
  INVX1 G38082 (.I(W47860), .ZN(O18810));
  INVX1 G38083 (.I(I1854), .ZN(W927));
  INVX1 G38084 (.I(I1826), .ZN(W913));
  INVX1 G38085 (.I(W14027), .ZN(O18860));
  INVX1 G38086 (.I(W3467), .ZN(O18859));
  INVX1 G38087 (.I(I1828), .ZN(W914));
  INVX1 G38088 (.I(W45089), .ZN(O18857));
  INVX1 G38089 (.I(W36910), .ZN(O18856));
  INVX1 G38090 (.I(I1832), .ZN(W916));
  INVX1 G38091 (.I(I1844), .ZN(W922));
  INVX1 G38092 (.I(I1848), .ZN(W924));
  INVX1 G38093 (.I(I1966), .ZN(W983));
  INVX1 G38094 (.I(I1856), .ZN(W928));
  INVX1 G38095 (.I(I1866), .ZN(W933));
  INVX1 G38096 (.I(I1868), .ZN(W934));
  INVX1 G38097 (.I(I1870), .ZN(W935));
  INVX1 G38098 (.I(W5784), .ZN(O18844));
  INVX1 G38099 (.I(W3135), .ZN(O18843));
  INVX1 G38100 (.I(I1878), .ZN(W939));
  INVX1 G38101 (.I(W43808), .ZN(O18841));
  INVX1 G38102 (.I(W33710), .ZN(O18770));
  INVX1 G38103 (.I(I1263), .ZN(W1017));
  INVX1 G38104 (.I(W23713), .ZN(O18779));
  INVX1 G38105 (.I(I1356), .ZN(W1018));
  INVX1 G38106 (.I(W299), .ZN(W1019));
  INVX1 G38107 (.I(W111), .ZN(W1022));
  INVX1 G38108 (.I(I234), .ZN(W1025));
  INVX1 G38109 (.I(I134), .ZN(W1026));
  INVX1 G38110 (.I(W4659), .ZN(O18773));
  INVX1 G38111 (.I(W16172), .ZN(O18771));
  INVX1 G38112 (.I(I238), .ZN(W1010));
  INVX1 G38113 (.I(W25), .ZN(W1028));
  INVX1 G38114 (.I(W28331), .ZN(W49987));
  INVX1 G38115 (.I(W7635), .ZN(O18767));
  INVX1 G38116 (.I(W848), .ZN(W1030));
  INVX1 G38117 (.I(W233), .ZN(W1032));
  INVX1 G38118 (.I(W11634), .ZN(O18762));
  INVX1 G38119 (.I(W14168), .ZN(O18761));
  INVX1 G38120 (.I(I1882), .ZN(W1036));
  INVX1 G38121 (.I(I1994), .ZN(W997));
  INVX1 G38122 (.I(I1970), .ZN(W985));
  INVX1 G38123 (.I(I1972), .ZN(W986));
  INVX1 G38124 (.I(W18791), .ZN(O18804));
  INVX1 G38125 (.I(W31202), .ZN(O18803));
  INVX1 G38126 (.I(W47122), .ZN(O18801));
  INVX1 G38127 (.I(I1988), .ZN(W994));
  INVX1 G38128 (.I(W29425), .ZN(O18798));
  INVX1 G38129 (.I(W46197), .ZN(O18797));
  INVX1 G38130 (.I(I1127), .ZN(W1147));
  INVX1 G38131 (.I(W18374), .ZN(O18795));
  INVX1 G38132 (.I(I1998), .ZN(W999));
  INVX1 G38133 (.I(W877), .ZN(W1001));
  INVX1 G38134 (.I(W9771), .ZN(O18790));
  INVX1 G38135 (.I(W38540), .ZN(O18788));
  INVX1 G38136 (.I(I566), .ZN(W1004));
  INVX1 G38137 (.I(W32057), .ZN(O18786));
  INVX1 G38138 (.I(W887), .ZN(W1008));
  INVX1 G38139 (.I(I1649), .ZN(W1292));
  INVX1 G38140 (.I(I1114), .ZN(W1277));
  INVX1 G38141 (.I(I1136), .ZN(W1286));
  INVX1 G38142 (.I(W36358), .ZN(O18510));
  INVX1 G38143 (.I(W12925), .ZN(O18509));
  INVX1 G38144 (.I(I1815), .ZN(W1289));
  INVX1 G38145 (.I(W13143), .ZN(O18507));
  INVX1 G38146 (.I(W40026), .ZN(O18506));
  INVX1 G38147 (.I(W609), .ZN(W1290));
  INVX1 G38148 (.I(I1065), .ZN(W1291));
  INVX1 G38149 (.I(W341), .ZN(W1276));
  INVX1 G38150 (.I(W882), .ZN(W1293));
  INVX1 G38151 (.I(W961), .ZN(O18502));
  INVX1 G38152 (.I(I116), .ZN(O18501));
  INVX1 G38153 (.I(W889), .ZN(W1296));
  INVX1 G38154 (.I(I1456), .ZN(W1298));
  INVX1 G38155 (.I(I626), .ZN(W1299));
  INVX1 G38156 (.I(W40513), .ZN(O18494));
  INVX1 G38157 (.I(I284), .ZN(W1300));
  INVX1 G38158 (.I(I1932), .ZN(W1251));
  INVX1 G38159 (.I(I885), .ZN(W1238));
  INVX1 G38160 (.I(I486), .ZN(W1239));
  INVX1 G38161 (.I(W691), .ZN(W1240));
  INVX1 G38162 (.I(W12), .ZN(W1243));
  INVX1 G38163 (.I(I1450), .ZN(W1245));
  INVX1 G38164 (.I(W417), .ZN(W1249));
  INVX1 G38165 (.I(W23361), .ZN(O18540));
  INVX1 G38166 (.I(W48600), .ZN(O18539));
  INVX1 G38167 (.I(I120), .ZN(W1250));
  INVX1 G38168 (.I(W48226), .ZN(O18492));
  INVX1 G38169 (.I(W46355), .ZN(O18533));
  INVX1 G38170 (.I(W33527), .ZN(O18532));
  INVX1 G38171 (.I(W137), .ZN(W1258));
  INVX1 G38172 (.I(W4503), .ZN(O18526));
  INVX1 G38173 (.I(I459), .ZN(W1270));
  INVX1 G38174 (.I(W41176), .ZN(O18522));
  INVX1 G38175 (.I(I23), .ZN(W1275));
  INVX1 G38176 (.I(W7166), .ZN(O18519));
  INVX1 G38177 (.I(I1552), .ZN(W1358));
  INVX1 G38178 (.I(I1594), .ZN(W1331));
  INVX1 G38179 (.I(W475), .ZN(W1334));
  INVX1 G38180 (.I(W31695), .ZN(O18465));
  INVX1 G38181 (.I(I850), .ZN(W1343));
  INVX1 G38182 (.I(I203), .ZN(W1346));
  INVX1 G38183 (.I(W44214), .ZN(O18460));
  INVX1 G38184 (.I(W15294), .ZN(O18459));
  INVX1 G38185 (.I(W763), .ZN(W1351));
  INVX1 G38186 (.I(W42311), .ZN(O18455));
  INVX1 G38187 (.I(W481), .ZN(W1328));
  INVX1 G38188 (.I(I729), .ZN(W1361));
  INVX1 G38189 (.I(W758), .ZN(W1362));
  INVX1 G38190 (.I(I1578), .ZN(W1363));
  INVX1 G38191 (.I(I759), .ZN(W1365));
  INVX1 G38192 (.I(W27227), .ZN(O18446));
  INVX1 G38193 (.I(I1166), .ZN(W1369));
  INVX1 G38194 (.I(W6984), .ZN(O18443));
  INVX1 G38195 (.I(W40826), .ZN(O18441));
  INVX1 G38196 (.I(W35), .ZN(W1309));
  INVX1 G38197 (.I(I878), .ZN(W1302));
  INVX1 G38198 (.I(W45679), .ZN(O18490));
  INVX1 G38199 (.I(W29211), .ZN(O18489));
  INVX1 G38200 (.I(W22732), .ZN(O18488));
  INVX1 G38201 (.I(W1138), .ZN(W1303));
  INVX1 G38202 (.I(W397), .ZN(O18486));
  INVX1 G38203 (.I(W42360), .ZN(O18483));
  INVX1 G38204 (.I(W21996), .ZN(O18482));
  INVX1 G38205 (.I(W17873), .ZN(O18549));
  INVX1 G38206 (.I(I1148), .ZN(W1312));
  INVX1 G38207 (.I(W47), .ZN(W1313));
  INVX1 G38208 (.I(I1165), .ZN(W1314));
  INVX1 G38209 (.I(W2172), .ZN(O18478));
  INVX1 G38210 (.I(I1322), .ZN(W1315));
  INVX1 G38211 (.I(W49293), .ZN(O18472));
  INVX1 G38212 (.I(I996), .ZN(W1324));
  INVX1 G38213 (.I(I989), .ZN(W1326));
  INVX1 G38214 (.I(I1858), .ZN(W1187));
  INVX1 G38215 (.I(W27736), .ZN(O18622));
  INVX1 G38216 (.I(I1278), .ZN(O18621));
  INVX1 G38217 (.I(W1221), .ZN(O18619));
  INVX1 G38218 (.I(W246), .ZN(W1176));
  INVX1 G38219 (.I(I619), .ZN(W1179));
  INVX1 G38220 (.I(I518), .ZN(W1180));
  INVX1 G38221 (.I(W6001), .ZN(O18612));
  INVX1 G38222 (.I(W69), .ZN(W1185));
  INVX1 G38223 (.I(W30497), .ZN(O18610));
  INVX1 G38224 (.I(W806), .ZN(O10));
  INVX1 G38225 (.I(W37158), .ZN(O18607));
  INVX1 G38226 (.I(W27638), .ZN(O18605));
  INVX1 G38227 (.I(I846), .ZN(W1193));
  INVX1 G38228 (.I(W660), .ZN(W1196));
  INVX1 G38229 (.I(W685), .ZN(W1197));
  INVX1 G38230 (.I(W28235), .ZN(O18598));
  INVX1 G38231 (.I(W975), .ZN(W1200));
  INVX1 G38232 (.I(W35139), .ZN(O18595));
  INVX1 G38233 (.I(W47074), .ZN(O18635));
  INVX1 G38234 (.I(W33375), .ZN(O18652));
  INVX1 G38235 (.I(I600), .ZN(W1151));
  INVX1 G38236 (.I(W22026), .ZN(O18646));
  INVX1 G38237 (.I(I246), .ZN(W1155));
  INVX1 G38238 (.I(W324), .ZN(W1157));
  INVX1 G38239 (.I(W14292), .ZN(O18642));
  INVX1 G38240 (.I(W30348), .ZN(O18641));
  INVX1 G38241 (.I(W33819), .ZN(O18639));
  INVX1 G38242 (.I(W19217), .ZN(O18638));
  INVX1 G38243 (.I(I1920), .ZN(W1203));
  INVX1 G38244 (.I(I605), .ZN(W1164));
  INVX1 G38245 (.I(W30556), .ZN(O18632));
  INVX1 G38246 (.I(I600), .ZN(W1167));
  INVX1 G38247 (.I(W2829), .ZN(O18629));
  INVX1 G38248 (.I(W31742), .ZN(O18627));
  INVX1 G38249 (.I(I62), .ZN(W1169));
  INVX1 G38250 (.I(W484), .ZN(O18625));
  INVX1 G38251 (.I(W83), .ZN(W1172));
  INVX1 G38252 (.I(I1152), .ZN(W1228));
  INVX1 G38253 (.I(I938), .ZN(W1216));
  INVX1 G38254 (.I(I1519), .ZN(W1218));
  INVX1 G38255 (.I(W2692), .ZN(O18572));
  INVX1 G38256 (.I(W4675), .ZN(O18571));
  INVX1 G38257 (.I(W32993), .ZN(O18570));
  INVX1 G38258 (.I(W42198), .ZN(O18569));
  INVX1 G38259 (.I(I1012), .ZN(W1220));
  INVX1 G38260 (.I(W38957), .ZN(O18566));
  INVX1 G38261 (.I(W101), .ZN(W1225));
  INVX1 G38262 (.I(W897), .ZN(W1215));
  INVX1 G38263 (.I(W16689), .ZN(O18562));
  INVX1 G38264 (.I(W37961), .ZN(O18561));
  INVX1 G38265 (.I(W5264), .ZN(O18560));
  INVX1 G38266 (.I(W44864), .ZN(O18556));
  INVX1 G38267 (.I(I503), .ZN(W1233));
  INVX1 G38268 (.I(W22269), .ZN(O18554));
  INVX1 G38269 (.I(W687), .ZN(W1234));
  INVX1 G38270 (.I(W32455), .ZN(O18552));
  INVX1 G38271 (.I(W12998), .ZN(O18584));
  INVX1 G38272 (.I(W655), .ZN(W1205));
  INVX1 G38273 (.I(W17197), .ZN(O18592));
  INVX1 G38274 (.I(W29421), .ZN(O18591));
  INVX1 G38275 (.I(W12767), .ZN(O18590));
  INVX1 G38276 (.I(W583), .ZN(W1207));
  INVX1 G38277 (.I(I1509), .ZN(W1208));
  INVX1 G38278 (.I(W26836), .ZN(O18587));
  INVX1 G38279 (.I(W49086), .ZN(O18585));
  INVX1 G38280 (.I(W2544), .ZN(W3523));
  INVX1 G38281 (.I(I579), .ZN(W1210));
  INVX1 G38282 (.I(W27594), .ZN(O18583));
  INVX1 G38283 (.I(W1053), .ZN(W1212));
  INVX1 G38284 (.I(W544), .ZN(W1213));
  INVX1 G38285 (.I(W36274), .ZN(O18579));
  INVX1 G38286 (.I(W37476), .ZN(O18578));
  INVX1 G38287 (.I(I1939), .ZN(W1214));
  INVX1 G38288 (.I(W15657), .ZN(O18576));
  INVX1 G38289 (.I(W5563), .ZN(W5787));
  INVX1 G38290 (.I(W1999), .ZN(O14485));
  INVX1 G38291 (.I(W3940), .ZN(W5772));
  INVX1 G38292 (.I(W889), .ZN(W5774));
  INVX1 G38293 (.I(I528), .ZN(W5775));
  INVX1 G38294 (.I(I499), .ZN(W5776));
  INVX1 G38295 (.I(W12223), .ZN(O14479));
  INVX1 G38296 (.I(W4428), .ZN(W5779));
  INVX1 G38297 (.I(I334), .ZN(W5780));
  INVX1 G38298 (.I(W3862), .ZN(W5783));
  INVX1 G38299 (.I(W271), .ZN(W5764));
  INVX1 G38300 (.I(W1332), .ZN(W5790));
  INVX1 G38301 (.I(W6265), .ZN(O14471));
  INVX1 G38302 (.I(W44789), .ZN(O14470));
  INVX1 G38303 (.I(W5219), .ZN(W5795));
  INVX1 G38304 (.I(W17285), .ZN(O14465));
  INVX1 G38305 (.I(W872), .ZN(W5799));
  INVX1 G38306 (.I(W2795), .ZN(W5809));
  INVX1 G38307 (.I(W25157), .ZN(O14459));
  INVX1 G38308 (.I(W23144), .ZN(O14498));
  INVX1 G38309 (.I(W40654), .ZN(O14511));
  INVX1 G38310 (.I(W17806), .ZN(O14509));
  INVX1 G38311 (.I(W20279), .ZN(O14508));
  INVX1 G38312 (.I(W40327), .ZN(O14507));
  INVX1 G38313 (.I(W35072), .ZN(W45179));
  INVX1 G38314 (.I(I467), .ZN(W5736));
  INVX1 G38315 (.I(W44183), .ZN(O14504));
  INVX1 G38316 (.I(W2670), .ZN(W5738));
  INVX1 G38317 (.I(W115), .ZN(W5751));
  INVX1 G38318 (.I(I1524), .ZN(W5810));
  INVX1 G38319 (.I(W535), .ZN(W5753));
  INVX1 G38320 (.I(W4771), .ZN(W5754));
  INVX1 G38321 (.I(W5428), .ZN(W45165));
  INVX1 G38322 (.I(W14973), .ZN(O14494));
  INVX1 G38323 (.I(I480), .ZN(W5755));
  INVX1 G38324 (.I(W467), .ZN(W5756));
  INVX1 G38325 (.I(W36861), .ZN(O14490));
  INVX1 G38326 (.I(I957), .ZN(W5759));
  INVX1 G38327 (.I(W265), .ZN(W5860));
  INVX1 G38328 (.I(W4977), .ZN(W5848));
  INVX1 G38329 (.I(I1220), .ZN(W5849));
  INVX1 G38330 (.I(W4384), .ZN(W5850));
  INVX1 G38331 (.I(W41456), .ZN(O14431));
  INVX1 G38332 (.I(W3873), .ZN(W5853));
  INVX1 G38333 (.I(W20074), .ZN(O14428));
  INVX1 G38334 (.I(W960), .ZN(W5855));
  INVX1 G38335 (.I(W1002), .ZN(W5857));
  INVX1 G38336 (.I(W40521), .ZN(O14425));
  INVX1 G38337 (.I(W5309), .ZN(W5842));
  INVX1 G38338 (.I(W1883), .ZN(O14423));
  INVX1 G38339 (.I(W36235), .ZN(O14422));
  INVX1 G38340 (.I(W17556), .ZN(W45075));
  INVX1 G38341 (.I(W23056), .ZN(O14421));
  INVX1 G38342 (.I(W12097), .ZN(O14420));
  INVX1 G38343 (.I(W5607), .ZN(W5865));
  INVX1 G38344 (.I(W2863), .ZN(W45068));
  INVX1 G38345 (.I(W42754), .ZN(O14414));
  INVX1 G38346 (.I(W2159), .ZN(W5822));
  INVX1 G38347 (.I(I1403), .ZN(O103));
  INVX1 G38348 (.I(W3633), .ZN(W5814));
  INVX1 G38349 (.I(W703), .ZN(O14456));
  INVX1 G38350 (.I(W20095), .ZN(O14454));
  INVX1 G38351 (.I(W38490), .ZN(O14453));
  INVX1 G38352 (.I(W1751), .ZN(W5817));
  INVX1 G38353 (.I(W20666), .ZN(O14451));
  INVX1 G38354 (.I(W18634), .ZN(W45111));
  INVX1 G38355 (.I(W5251), .ZN(O104));
  INVX1 G38356 (.I(W18990), .ZN(O14512));
  INVX1 G38357 (.I(W15166), .ZN(O14446));
  INVX1 G38358 (.I(W2748), .ZN(W5830));
  INVX1 G38359 (.I(W1198), .ZN(W5832));
  INVX1 G38360 (.I(W17252), .ZN(O14442));
  INVX1 G38361 (.I(W31873), .ZN(O14441));
  INVX1 G38362 (.I(W44844), .ZN(O14440));
  INVX1 G38363 (.I(W2193), .ZN(O14438));
  INVX1 G38364 (.I(W5633), .ZN(W5838));
  INVX1 G38365 (.I(W3808), .ZN(O96));
  INVX1 G38366 (.I(W1567), .ZN(W5650));
  INVX1 G38367 (.I(W38892), .ZN(W45269));
  INVX1 G38368 (.I(W9378), .ZN(W45267));
  INVX1 G38369 (.I(W30747), .ZN(O14576));
  INVX1 G38370 (.I(I1477), .ZN(W45264));
  INVX1 G38371 (.I(W531), .ZN(W5654));
  INVX1 G38372 (.I(W35440), .ZN(O14573));
  INVX1 G38373 (.I(W338), .ZN(W5658));
  INVX1 G38374 (.I(W2363), .ZN(W5659));
  INVX1 G38375 (.I(W5254), .ZN(W5649));
  INVX1 G38376 (.I(W27770), .ZN(W45255));
  INVX1 G38377 (.I(W3859), .ZN(W5667));
  INVX1 G38378 (.I(W5198), .ZN(W45251));
  INVX1 G38379 (.I(I538), .ZN(W5669));
  INVX1 G38380 (.I(W18165), .ZN(O14563));
  INVX1 G38381 (.I(W12083), .ZN(O14559));
  INVX1 G38382 (.I(W22522), .ZN(O14558));
  INVX1 G38383 (.I(W39233), .ZN(W45237));
  INVX1 G38384 (.I(W17442), .ZN(O14590));
  INVX1 G38385 (.I(W3085), .ZN(W5622));
  INVX1 G38386 (.I(W27075), .ZN(O14598));
  INVX1 G38387 (.I(W30138), .ZN(O14596));
  INVX1 G38388 (.I(W140), .ZN(O14595));
  INVX1 G38389 (.I(I1809), .ZN(W5624));
  INVX1 G38390 (.I(W25034), .ZN(O14593));
  INVX1 G38391 (.I(W2953), .ZN(W5625));
  INVX1 G38392 (.I(W5520), .ZN(W5627));
  INVX1 G38393 (.I(W3065), .ZN(W5629));
  INVX1 G38394 (.I(W366), .ZN(W5683));
  INVX1 G38395 (.I(I55), .ZN(W5631));
  INVX1 G38396 (.I(I358), .ZN(W5633));
  INVX1 G38397 (.I(I102), .ZN(W5634));
  INVX1 G38398 (.I(W1953), .ZN(W5640));
  INVX1 G38399 (.I(W2917), .ZN(W5644));
  INVX1 G38400 (.I(W20059), .ZN(O14583));
  INVX1 G38401 (.I(W563), .ZN(W5645));
  INVX1 G38402 (.I(I1799), .ZN(W5648));
  INVX1 G38403 (.I(W4005), .ZN(W5719));
  INVX1 G38404 (.I(W35454), .ZN(O14532));
  INVX1 G38405 (.I(W111), .ZN(W5712));
  INVX1 G38406 (.I(W30665), .ZN(W45205));
  INVX1 G38407 (.I(W4157), .ZN(W5713));
  INVX1 G38408 (.I(W30086), .ZN(O14530));
  INVX1 G38409 (.I(W6004), .ZN(O14529));
  INVX1 G38410 (.I(W2195), .ZN(O98));
  INVX1 G38411 (.I(W7565), .ZN(O14525));
  INVX1 G38412 (.I(W4019), .ZN(W5718));
  INVX1 G38413 (.I(W19638), .ZN(W45209));
  INVX1 G38414 (.I(W5271), .ZN(W5721));
  INVX1 G38415 (.I(W1386), .ZN(W5723));
  INVX1 G38416 (.I(I172), .ZN(W5725));
  INVX1 G38417 (.I(W4412), .ZN(W5726));
  INVX1 G38418 (.I(W1030), .ZN(W5727));
  INVX1 G38419 (.I(W747), .ZN(W5728));
  INVX1 G38420 (.I(I1025), .ZN(W5729));
  INVX1 G38421 (.I(W31061), .ZN(O14514));
  INVX1 G38422 (.I(W31566), .ZN(O14547));
  INVX1 G38423 (.I(W5147), .ZN(W5685));
  INVX1 G38424 (.I(W24307), .ZN(O14554));
  INVX1 G38425 (.I(I1875), .ZN(W5686));
  INVX1 G38426 (.I(W19092), .ZN(O14553));
  INVX1 G38427 (.I(W663), .ZN(W5687));
  INVX1 G38428 (.I(W39819), .ZN(O14551));
  INVX1 G38429 (.I(W2754), .ZN(O14549));
  INVX1 G38430 (.I(I1069), .ZN(W45225));
  INVX1 G38431 (.I(W13190), .ZN(O14412));
  INVX1 G38432 (.I(W1349), .ZN(O14546));
  INVX1 G38433 (.I(W4215), .ZN(W5694));
  INVX1 G38434 (.I(W5167), .ZN(W5695));
  INVX1 G38435 (.I(W2226), .ZN(W5699));
  INVX1 G38436 (.I(W2032), .ZN(W5700));
  INVX1 G38437 (.I(W43319), .ZN(O14540));
  INVX1 G38438 (.I(W4677), .ZN(O14538));
  INVX1 G38439 (.I(W42180), .ZN(W45211));
  INVX1 G38440 (.I(W502), .ZN(W6031));
  INVX1 G38441 (.I(W3994), .ZN(W6014));
  INVX1 G38442 (.I(W22530), .ZN(O14289));
  INVX1 G38443 (.I(W3331), .ZN(W6016));
  INVX1 G38444 (.I(W28307), .ZN(O14287));
  INVX1 G38445 (.I(W8669), .ZN(O14286));
  INVX1 G38446 (.I(I1347), .ZN(W6017));
  INVX1 G38447 (.I(W3712), .ZN(W6020));
  INVX1 G38448 (.I(W34400), .ZN(O14280));
  INVX1 G38449 (.I(W3929), .ZN(W6024));
  INVX1 G38450 (.I(W43377), .ZN(O14293));
  INVX1 G38451 (.I(W4741), .ZN(W6032));
  INVX1 G38452 (.I(W4859), .ZN(W6033));
  INVX1 G38453 (.I(W39812), .ZN(W44901));
  INVX1 G38454 (.I(W32455), .ZN(O14275));
  INVX1 G38455 (.I(I235), .ZN(W6037));
  INVX1 G38456 (.I(W826), .ZN(W6038));
  INVX1 G38457 (.I(W3171), .ZN(W6042));
  INVX1 G38458 (.I(I233), .ZN(W6043));
  INVX1 G38459 (.I(W2550), .ZN(W5978));
  INVX1 G38460 (.I(W827), .ZN(W5968));
  INVX1 G38461 (.I(W40854), .ZN(O14315));
  INVX1 G38462 (.I(W7246), .ZN(O14314));
  INVX1 G38463 (.I(I768), .ZN(W44950));
  INVX1 G38464 (.I(W5540), .ZN(W5971));
  INVX1 G38465 (.I(W4259), .ZN(W5972));
  INVX1 G38466 (.I(I431), .ZN(W5974));
  INVX1 G38467 (.I(W2176), .ZN(W5977));
  INVX1 G38468 (.I(W4276), .ZN(O14309));
  INVX1 G38469 (.I(W212), .ZN(W6044));
  INVX1 G38470 (.I(W2739), .ZN(O113));
  INVX1 G38471 (.I(W4081), .ZN(O114));
  INVX1 G38472 (.I(W14933), .ZN(O14303));
  INVX1 G38473 (.I(W2006), .ZN(W5999));
  INVX1 G38474 (.I(W1545), .ZN(W6002));
  INVX1 G38475 (.I(I1256), .ZN(W6003));
  INVX1 G38476 (.I(W5887), .ZN(W6004));
  INVX1 G38477 (.I(W3626), .ZN(W6007));
  INVX1 G38478 (.I(W31356), .ZN(O14238));
  INVX1 G38479 (.I(W100), .ZN(W6065));
  INVX1 G38480 (.I(W4737), .ZN(W44862));
  INVX1 G38481 (.I(W21551), .ZN(W44861));
  INVX1 G38482 (.I(W2833), .ZN(W6066));
  INVX1 G38483 (.I(W2340), .ZN(W6069));
  INVX1 G38484 (.I(I1742), .ZN(W6070));
  INVX1 G38485 (.I(I1243), .ZN(W6071));
  INVX1 G38486 (.I(I44), .ZN(W6072));
  INVX1 G38487 (.I(W301), .ZN(W6074));
  INVX1 G38488 (.I(W34449), .ZN(W44864));
  INVX1 G38489 (.I(W4428), .ZN(W6075));
  INVX1 G38490 (.I(W5109), .ZN(W6076));
  INVX1 G38491 (.I(W17017), .ZN(O14234));
  INVX1 G38492 (.I(W4563), .ZN(W6081));
  INVX1 G38493 (.I(W30160), .ZN(O14231));
  INVX1 G38494 (.I(I557), .ZN(W6088));
  INVX1 G38495 (.I(W4055), .ZN(W6093));
  INVX1 G38496 (.I(W10667), .ZN(W44836));
  INVX1 G38497 (.I(W21731), .ZN(O14258));
  INVX1 G38498 (.I(W26165), .ZN(O14267));
  INVX1 G38499 (.I(W36342), .ZN(O14265));
  INVX1 G38500 (.I(W18926), .ZN(O14264));
  INVX1 G38501 (.I(W41643), .ZN(O14263));
  INVX1 G38502 (.I(W33079), .ZN(O14262));
  INVX1 G38503 (.I(W20807), .ZN(O14261));
  INVX1 G38504 (.I(W317), .ZN(W6051));
  INVX1 G38505 (.I(W41235), .ZN(O14259));
  INVX1 G38506 (.I(I954), .ZN(W5965));
  INVX1 G38507 (.I(W19461), .ZN(O14257));
  INVX1 G38508 (.I(W27889), .ZN(O14254));
  INVX1 G38509 (.I(W523), .ZN(W6058));
  INVX1 G38510 (.I(W16685), .ZN(O14250));
  INVX1 G38511 (.I(W36825), .ZN(O14249));
  INVX1 G38512 (.I(W32049), .ZN(W44868));
  INVX1 G38513 (.I(I624), .ZN(W6063));
  INVX1 G38514 (.I(W13569), .ZN(O14247));
  INVX1 G38515 (.I(I1238), .ZN(W5903));
  INVX1 G38516 (.I(W40049), .ZN(O14385));
  INVX1 G38517 (.I(W35690), .ZN(O14383));
  INVX1 G38518 (.I(I1317), .ZN(W5896));
  INVX1 G38519 (.I(W24946), .ZN(O14382));
  INVX1 G38520 (.I(W7245), .ZN(O14381));
  INVX1 G38521 (.I(W846), .ZN(W5898));
  INVX1 G38522 (.I(W3256), .ZN(O14379));
  INVX1 G38523 (.I(W5077), .ZN(W5899));
  INVX1 G38524 (.I(W39315), .ZN(O14377));
  INVX1 G38525 (.I(W2329), .ZN(W5892));
  INVX1 G38526 (.I(W42305), .ZN(O14375));
  INVX1 G38527 (.I(W3897), .ZN(W5907));
  INVX1 G38528 (.I(W27140), .ZN(O14372));
  INVX1 G38529 (.I(I1348), .ZN(W5909));
  INVX1 G38530 (.I(W16990), .ZN(W45018));
  INVX1 G38531 (.I(I1980), .ZN(W5911));
  INVX1 G38532 (.I(W33218), .ZN(O14367));
  INVX1 G38533 (.I(W5123), .ZN(W5912));
  INVX1 G38534 (.I(W5229), .ZN(W5877));
  INVX1 G38535 (.I(W30029), .ZN(O14411));
  INVX1 G38536 (.I(W21964), .ZN(O14410));
  INVX1 G38537 (.I(W4071), .ZN(O14409));
  INVX1 G38538 (.I(W10851), .ZN(O14408));
  INVX1 G38539 (.I(W5856), .ZN(W5871));
  INVX1 G38540 (.I(W9632), .ZN(O14406));
  INVX1 G38541 (.I(W39479), .ZN(O14405));
  INVX1 G38542 (.I(W11800), .ZN(O14404));
  INVX1 G38543 (.I(W2812), .ZN(W5874));
  INVX1 G38544 (.I(W19739), .ZN(O14365));
  INVX1 G38545 (.I(I1819), .ZN(W5878));
  INVX1 G38546 (.I(W19570), .ZN(O14399));
  INVX1 G38547 (.I(W23515), .ZN(O14398));
  INVX1 G38548 (.I(W27026), .ZN(O14397));
  INVX1 G38549 (.I(I1000), .ZN(W5887));
  INVX1 G38550 (.I(W3240), .ZN(W5888));
  INVX1 G38551 (.I(W5660), .ZN(W5889));
  INVX1 G38552 (.I(W6297), .ZN(O14388));
  INVX1 G38553 (.I(W4641), .ZN(W5959));
  INVX1 G38554 (.I(W30557), .ZN(O14342));
  INVX1 G38555 (.I(W44660), .ZN(O14339));
  INVX1 G38556 (.I(W44794), .ZN(O14338));
  INVX1 G38557 (.I(W5816), .ZN(W5950));
  INVX1 G38558 (.I(W3741), .ZN(O108));
  INVX1 G38559 (.I(W42542), .ZN(W44974));
  INVX1 G38560 (.I(W5198), .ZN(O14336));
  INVX1 G38561 (.I(W2311), .ZN(W5953));
  INVX1 G38562 (.I(W11430), .ZN(O14331));
  INVX1 G38563 (.I(W850), .ZN(W5945));
  INVX1 G38564 (.I(W30095), .ZN(O14328));
  INVX1 G38565 (.I(W3424), .ZN(W5960));
  INVX1 G38566 (.I(W104), .ZN(O14326));
  INVX1 G38567 (.I(W40783), .ZN(O14325));
  INVX1 G38568 (.I(W17464), .ZN(O14323));
  INVX1 G38569 (.I(W5749), .ZN(W5962));
  INVX1 G38570 (.I(W36950), .ZN(O14321));
  INVX1 G38571 (.I(W14615), .ZN(O14320));
  INVX1 G38572 (.I(W2779), .ZN(W5932));
  INVX1 G38573 (.I(W4565), .ZN(W5916));
  INVX1 G38574 (.I(I1404), .ZN(W5918));
  INVX1 G38575 (.I(W3307), .ZN(W5920));
  INVX1 G38576 (.I(W39725), .ZN(O14358));
  INVX1 G38577 (.I(I1556), .ZN(O14355));
  INVX1 G38578 (.I(W5), .ZN(W5925));
  INVX1 G38579 (.I(W44908), .ZN(O14353));
  INVX1 G38580 (.I(W44035), .ZN(W44999));
  INVX1 G38581 (.I(W30817), .ZN(O14601));
  INVX1 G38582 (.I(W4175), .ZN(W5934));
  INVX1 G38583 (.I(W2741), .ZN(W5936));
  INVX1 G38584 (.I(I234), .ZN(W5938));
  INVX1 G38585 (.I(W5331), .ZN(W5940));
  INVX1 G38586 (.I(W5378), .ZN(W5941));
  INVX1 G38587 (.I(W44441), .ZN(O14347));
  INVX1 G38588 (.I(W11987), .ZN(O14346));
  INVX1 G38589 (.I(W3475), .ZN(W5942));
  INVX1 G38590 (.I(W5104), .ZN(W5348));
  INVX1 G38591 (.I(I1217), .ZN(W5336));
  INVX1 G38592 (.I(I1563), .ZN(W5337));
  INVX1 G38593 (.I(W30505), .ZN(O14844));
  INVX1 G38594 (.I(W32411), .ZN(W45595));
  INVX1 G38595 (.I(I223), .ZN(W5340));
  INVX1 G38596 (.I(W17982), .ZN(O14842));
  INVX1 G38597 (.I(W10249), .ZN(O14841));
  INVX1 G38598 (.I(I457), .ZN(W5344));
  INVX1 G38599 (.I(W44226), .ZN(O14839));
  INVX1 G38600 (.I(W12418), .ZN(O14847));
  INVX1 G38601 (.I(W27648), .ZN(O14837));
  INVX1 G38602 (.I(W4897), .ZN(W5350));
  INVX1 G38603 (.I(I92), .ZN(W5354));
  INVX1 G38604 (.I(W16402), .ZN(O14834));
  INVX1 G38605 (.I(W4974), .ZN(W5355));
  INVX1 G38606 (.I(W41256), .ZN(O14831));
  INVX1 G38607 (.I(I1064), .ZN(W5361));
  INVX1 G38608 (.I(W29310), .ZN(O14829));
  INVX1 G38609 (.I(W1239), .ZN(W5322));
  INVX1 G38610 (.I(W3894), .ZN(W5309));
  INVX1 G38611 (.I(W31594), .ZN(O14870));
  INVX1 G38612 (.I(W2586), .ZN(W5310));
  INVX1 G38613 (.I(W4642), .ZN(W5311));
  INVX1 G38614 (.I(W1249), .ZN(W5312));
  INVX1 G38615 (.I(W13899), .ZN(O14866));
  INVX1 G38616 (.I(W10587), .ZN(O14863));
  INVX1 G38617 (.I(W40184), .ZN(O14862));
  INVX1 G38618 (.I(W832), .ZN(W5315));
  INVX1 G38619 (.I(W30017), .ZN(O14828));
  INVX1 G38620 (.I(W3287), .ZN(O14854));
  INVX1 G38621 (.I(W2082), .ZN(W5331));
  INVX1 G38622 (.I(W5356), .ZN(W45606));
  INVX1 G38623 (.I(W2339), .ZN(W5333));
  INVX1 G38624 (.I(W20507), .ZN(O14851));
  INVX1 G38625 (.I(I879), .ZN(O14850));
  INVX1 G38626 (.I(W2590), .ZN(W5335));
  INVX1 G38627 (.I(W25979), .ZN(O14848));
  INVX1 G38628 (.I(W44988), .ZN(O14795));
  INVX1 G38629 (.I(W15771), .ZN(O14805));
  INVX1 G38630 (.I(W40643), .ZN(O14804));
  INVX1 G38631 (.I(I1298), .ZN(W5396));
  INVX1 G38632 (.I(W26305), .ZN(O14801));
  INVX1 G38633 (.I(W4109), .ZN(O14800));
  INVX1 G38634 (.I(W4809), .ZN(W5398));
  INVX1 G38635 (.I(W45018), .ZN(O14797));
  INVX1 G38636 (.I(W32983), .ZN(W45533));
  INVX1 G38637 (.I(W8951), .ZN(O14796));
  INVX1 G38638 (.I(W4272), .ZN(O84));
  INVX1 G38639 (.I(W2982), .ZN(W5404));
  INVX1 G38640 (.I(I932), .ZN(W5407));
  INVX1 G38641 (.I(W13824), .ZN(W45525));
  INVX1 G38642 (.I(W3782), .ZN(W5408));
  INVX1 G38643 (.I(I324), .ZN(W5410));
  INVX1 G38644 (.I(I1550), .ZN(W5411));
  INVX1 G38645 (.I(W30770), .ZN(O14788));
  INVX1 G38646 (.I(W3224), .ZN(O14787));
  INVX1 G38647 (.I(W10202), .ZN(W45559));
  INVX1 G38648 (.I(W40781), .ZN(W45574));
  INVX1 G38649 (.I(W44352), .ZN(O14826));
  INVX1 G38650 (.I(I784), .ZN(W5363));
  INVX1 G38651 (.I(W40296), .ZN(O14825));
  INVX1 G38652 (.I(W238), .ZN(W5368));
  INVX1 G38653 (.I(W30661), .ZN(W45564));
  INVX1 G38654 (.I(W20800), .ZN(O14821));
  INVX1 G38655 (.I(W39050), .ZN(O14820));
  INVX1 G38656 (.I(W13139), .ZN(O14871));
  INVX1 G38657 (.I(W27885), .ZN(W45558));
  INVX1 G38658 (.I(W28824), .ZN(O14817));
  INVX1 G38659 (.I(W4516), .ZN(W5378));
  INVX1 G38660 (.I(W4093), .ZN(W5379));
  INVX1 G38661 (.I(W10260), .ZN(O14813));
  INVX1 G38662 (.I(W1747), .ZN(W5383));
  INVX1 G38663 (.I(W4209), .ZN(W5387));
  INVX1 G38664 (.I(W43055), .ZN(O14808));
  INVX1 G38665 (.I(W3074), .ZN(W5238));
  INVX1 G38666 (.I(W1272), .ZN(W5230));
  INVX1 G38667 (.I(W32132), .ZN(O14943));
  INVX1 G38668 (.I(W41994), .ZN(O14942));
  INVX1 G38669 (.I(W14156), .ZN(O14941));
  INVX1 G38670 (.I(W1077), .ZN(W5233));
  INVX1 G38671 (.I(W137), .ZN(O78));
  INVX1 G38672 (.I(W5033), .ZN(O14937));
  INVX1 G38673 (.I(W2068), .ZN(W5237));
  INVX1 G38674 (.I(W30579), .ZN(O14935));
  INVX1 G38675 (.I(W22922), .ZN(W45710));
  INVX1 G38676 (.I(W22387), .ZN(O14933));
  INVX1 G38677 (.I(W1816), .ZN(W5239));
  INVX1 G38678 (.I(W19), .ZN(O14931));
  INVX1 G38679 (.I(W907), .ZN(W45693));
  INVX1 G38680 (.I(W25387), .ZN(W45692));
  INVX1 G38681 (.I(W1703), .ZN(W5241));
  INVX1 G38682 (.I(W26248), .ZN(O14928));
  INVX1 G38683 (.I(W2356), .ZN(W5243));
  INVX1 G38684 (.I(W4378), .ZN(W5219));
  INVX1 G38685 (.I(W29616), .ZN(O14960));
  INVX1 G38686 (.I(W43380), .ZN(W45732));
  INVX1 G38687 (.I(W1225), .ZN(W5215));
  INVX1 G38688 (.I(W39193), .ZN(O14958));
  INVX1 G38689 (.I(W23076), .ZN(O14957));
  INVX1 G38690 (.I(I1944), .ZN(W45728));
  INVX1 G38691 (.I(W37597), .ZN(W45726));
  INVX1 G38692 (.I(W41911), .ZN(O14955));
  INVX1 G38693 (.I(I1225), .ZN(W5218));
  INVX1 G38694 (.I(W42536), .ZN(O14926));
  INVX1 G38695 (.I(W27380), .ZN(O14951));
  INVX1 G38696 (.I(W40174), .ZN(O14950));
  INVX1 G38697 (.I(W3522), .ZN(W5222));
  INVX1 G38698 (.I(I1950), .ZN(W5223));
  INVX1 G38699 (.I(I116), .ZN(W5224));
  INVX1 G38700 (.I(W3047), .ZN(W5225));
  INVX1 G38701 (.I(W2830), .ZN(W45714));
  INVX1 G38702 (.I(W3857), .ZN(W5227));
  INVX1 G38703 (.I(W598), .ZN(W5299));
  INVX1 G38704 (.I(W30273), .ZN(O14897));
  INVX1 G38705 (.I(W6367), .ZN(O14896));
  INVX1 G38706 (.I(W10164), .ZN(O14895));
  INVX1 G38707 (.I(W19003), .ZN(O14894));
  INVX1 G38708 (.I(W2140), .ZN(W5286));
  INVX1 G38709 (.I(W25803), .ZN(O14890));
  INVX1 G38710 (.I(W28684), .ZN(O14885));
  INVX1 G38711 (.I(W1439), .ZN(W5297));
  INVX1 G38712 (.I(W2014), .ZN(W5298));
  INVX1 G38713 (.I(W19426), .ZN(O14899));
  INVX1 G38714 (.I(W3005), .ZN(W5300));
  INVX1 G38715 (.I(W45205), .ZN(O14880));
  INVX1 G38716 (.I(W21461), .ZN(O14879));
  INVX1 G38717 (.I(W1012), .ZN(W5304));
  INVX1 G38718 (.I(W21270), .ZN(O14876));
  INVX1 G38719 (.I(W28002), .ZN(O14875));
  INVX1 G38720 (.I(W32618), .ZN(O14874));
  INVX1 G38721 (.I(W3812), .ZN(W5305));
  INVX1 G38722 (.I(W963), .ZN(W5259));
  INVX1 G38723 (.I(W4518), .ZN(W5244));
  INVX1 G38724 (.I(I685), .ZN(W5248));
  INVX1 G38725 (.I(W3720), .ZN(W5250));
  INVX1 G38726 (.I(W594), .ZN(W5251));
  INVX1 G38727 (.I(W355), .ZN(W5252));
  INVX1 G38728 (.I(W8180), .ZN(W45679));
  INVX1 G38729 (.I(W30679), .ZN(W45678));
  INVX1 G38730 (.I(W37190), .ZN(O14917));
  INVX1 G38731 (.I(W1381), .ZN(W5412));
  INVX1 G38732 (.I(W38917), .ZN(O14915));
  INVX1 G38733 (.I(W5073), .ZN(O14914));
  INVX1 G38734 (.I(W961), .ZN(W5263));
  INVX1 G38735 (.I(I1760), .ZN(W5266));
  INVX1 G38736 (.I(W1505), .ZN(W5270));
  INVX1 G38737 (.I(W434), .ZN(W5272));
  INVX1 G38738 (.I(W678), .ZN(W5276));
  INVX1 G38739 (.I(W18), .ZN(W5277));
  INVX1 G38740 (.I(I121), .ZN(W5554));
  INVX1 G38741 (.I(I44), .ZN(O91));
  INVX1 G38742 (.I(W22544), .ZN(W45373));
  INVX1 G38743 (.I(W1223), .ZN(W5539));
  INVX1 G38744 (.I(W4570), .ZN(O92));
  INVX1 G38745 (.I(I1432), .ZN(W5545));
  INVX1 G38746 (.I(W43709), .ZN(O14660));
  INVX1 G38747 (.I(W2118), .ZN(O93));
  INVX1 G38748 (.I(W4835), .ZN(W5551));
  INVX1 G38749 (.I(W3162), .ZN(W5552));
  INVX1 G38750 (.I(W9375), .ZN(O14666));
  INVX1 G38751 (.I(W27346), .ZN(O14658));
  INVX1 G38752 (.I(W22759), .ZN(O14657));
  INVX1 G38753 (.I(W1645), .ZN(W5555));
  INVX1 G38754 (.I(W3477), .ZN(W5556));
  INVX1 G38755 (.I(W44861), .ZN(O14654));
  INVX1 G38756 (.I(W32280), .ZN(O14653));
  INVX1 G38757 (.I(W6419), .ZN(O14652));
  INVX1 G38758 (.I(I1760), .ZN(W5557));
  INVX1 G38759 (.I(I1758), .ZN(O14679));
  INVX1 G38760 (.I(I132), .ZN(O14696));
  INVX1 G38761 (.I(W3005), .ZN(W5506));
  INVX1 G38762 (.I(W3007), .ZN(O14694));
  INVX1 G38763 (.I(W710), .ZN(W5508));
  INVX1 G38764 (.I(W3166), .ZN(W5510));
  INVX1 G38765 (.I(W32451), .ZN(O14686));
  INVX1 G38766 (.I(W3297), .ZN(O88));
  INVX1 G38767 (.I(W1481), .ZN(W5517));
  INVX1 G38768 (.I(W41245), .ZN(O14681));
  INVX1 G38769 (.I(W1942), .ZN(W5560));
  INVX1 G38770 (.I(W2), .ZN(O14678));
  INVX1 G38771 (.I(W30708), .ZN(O14676));
  INVX1 G38772 (.I(W2756), .ZN(W5523));
  INVX1 G38773 (.I(I294), .ZN(W5524));
  INVX1 G38774 (.I(W2568), .ZN(W5528));
  INVX1 G38775 (.I(W2062), .ZN(W5531));
  INVX1 G38776 (.I(W1187), .ZN(W5533));
  INVX1 G38777 (.I(W7170), .ZN(O14667));
  INVX1 G38778 (.I(W785), .ZN(W5600));
  INVX1 G38779 (.I(I1928), .ZN(W5581));
  INVX1 G38780 (.I(W2282), .ZN(W5583));
  INVX1 G38781 (.I(I1506), .ZN(W5588));
  INVX1 G38782 (.I(W13484), .ZN(O14624));
  INVX1 G38783 (.I(W27193), .ZN(O14623));
  INVX1 G38784 (.I(W1574), .ZN(W5594));
  INVX1 G38785 (.I(W2373), .ZN(W5597));
  INVX1 G38786 (.I(W3981), .ZN(O14618));
  INVX1 G38787 (.I(W25677), .ZN(O14615));
  INVX1 G38788 (.I(W3750), .ZN(W5579));
  INVX1 G38789 (.I(W36780), .ZN(O14612));
  INVX1 G38790 (.I(W1401), .ZN(W5604));
  INVX1 G38791 (.I(W2913), .ZN(W5605));
  INVX1 G38792 (.I(W50), .ZN(W5610));
  INVX1 G38793 (.I(W103), .ZN(W5611));
  INVX1 G38794 (.I(W29000), .ZN(O14604));
  INVX1 G38795 (.I(I784), .ZN(W5614));
  INVX1 G38796 (.I(W4675), .ZN(W5616));
  INVX1 G38797 (.I(I715), .ZN(W5567));
  INVX1 G38798 (.I(W3185), .ZN(W5563));
  INVX1 G38799 (.I(W43685), .ZN(O14645));
  INVX1 G38800 (.I(W15452), .ZN(W45349));
  INVX1 G38801 (.I(I962), .ZN(O94));
  INVX1 G38802 (.I(W15314), .ZN(O14643));
  INVX1 G38803 (.I(W1430), .ZN(W5565));
  INVX1 G38804 (.I(W5442), .ZN(O14641));
  INVX1 G38805 (.I(W38161), .ZN(O14640));
  INVX1 G38806 (.I(W4363), .ZN(W5502));
  INVX1 G38807 (.I(I820), .ZN(W5572));
  INVX1 G38808 (.I(W2162), .ZN(W5573));
  INVX1 G38809 (.I(I1118), .ZN(W45337));
  INVX1 G38810 (.I(I1523), .ZN(W5576));
  INVX1 G38811 (.I(W33110), .ZN(O14633));
  INVX1 G38812 (.I(W20514), .ZN(O14632));
  INVX1 G38813 (.I(W4178), .ZN(W5577));
  INVX1 G38814 (.I(W17378), .ZN(O14629));
  INVX1 G38815 (.I(W3206), .ZN(O14752));
  INVX1 G38816 (.I(W15647), .ZN(O14762));
  INVX1 G38817 (.I(W42111), .ZN(O14761));
  INVX1 G38818 (.I(W20546), .ZN(O14760));
  INVX1 G38819 (.I(W3708), .ZN(W5439));
  INVX1 G38820 (.I(W2704), .ZN(W5440));
  INVX1 G38821 (.I(W8035), .ZN(O14757));
  INVX1 G38822 (.I(W4715), .ZN(W5444));
  INVX1 G38823 (.I(W294), .ZN(W5447));
  INVX1 G38824 (.I(W484), .ZN(W5448));
  INVX1 G38825 (.I(W1660), .ZN(W5433));
  INVX1 G38826 (.I(W1968), .ZN(W5450));
  INVX1 G38827 (.I(W6433), .ZN(O14750));
  INVX1 G38828 (.I(I1129), .ZN(O14749));
  INVX1 G38829 (.I(W3939), .ZN(W5451));
  INVX1 G38830 (.I(W10611), .ZN(O14747));
  INVX1 G38831 (.I(I1540), .ZN(W5453));
  INVX1 G38832 (.I(W1990), .ZN(W5457));
  INVX1 G38833 (.I(W251), .ZN(W5458));
  INVX1 G38834 (.I(I1477), .ZN(W5419));
  INVX1 G38835 (.I(W7175), .ZN(O14785));
  INVX1 G38836 (.I(W22316), .ZN(W45517));
  INVX1 G38837 (.I(I1743), .ZN(W5416));
  INVX1 G38838 (.I(W38446), .ZN(O14782));
  INVX1 G38839 (.I(W2742), .ZN(W5417));
  INVX1 G38840 (.I(I1058), .ZN(W5418));
  INVX1 G38841 (.I(W15439), .ZN(O14779));
  INVX1 G38842 (.I(W19290), .ZN(O14778));
  INVX1 G38843 (.I(W44071), .ZN(O14777));
  INVX1 G38844 (.I(W1082), .ZN(W5460));
  INVX1 G38845 (.I(W2122), .ZN(W5420));
  INVX1 G38846 (.I(W818), .ZN(W5425));
  INVX1 G38847 (.I(I192), .ZN(W5426));
  INVX1 G38848 (.I(W37019), .ZN(O14770));
  INVX1 G38849 (.I(I1798), .ZN(O14769));
  INVX1 G38850 (.I(W4266), .ZN(W5429));
  INVX1 G38851 (.I(W3925), .ZN(W5431));
  INVX1 G38852 (.I(W17122), .ZN(O14765));
  INVX1 G38853 (.I(W247), .ZN(W5494));
  INVX1 G38854 (.I(W39778), .ZN(O14717));
  INVX1 G38855 (.I(W399), .ZN(W5488));
  INVX1 G38856 (.I(W18763), .ZN(O14713));
  INVX1 G38857 (.I(I147), .ZN(W5492));
  INVX1 G38858 (.I(W40477), .ZN(W45429));
  INVX1 G38859 (.I(W14884), .ZN(O14711));
  INVX1 G38860 (.I(W22934), .ZN(O14710));
  INVX1 G38861 (.I(W20637), .ZN(W45426));
  INVX1 G38862 (.I(W13490), .ZN(O14708));
  INVX1 G38863 (.I(W391), .ZN(W5486));
  INVX1 G38864 (.I(W12397), .ZN(O14705));
  INVX1 G38865 (.I(W1225), .ZN(W5497));
  INVX1 G38866 (.I(W7603), .ZN(O14703));
  INVX1 G38867 (.I(W12822), .ZN(O14702));
  INVX1 G38868 (.I(W13085), .ZN(O14701));
  INVX1 G38869 (.I(I1545), .ZN(W5498));
  INVX1 G38870 (.I(I873), .ZN(W5500));
  INVX1 G38871 (.I(W14076), .ZN(W45413));
  INVX1 G38872 (.I(W3283), .ZN(W5468));
  INVX1 G38873 (.I(W26165), .ZN(O14742));
  INVX1 G38874 (.I(W32624), .ZN(O14741));
  INVX1 G38875 (.I(W41833), .ZN(O14740));
  INVX1 G38876 (.I(W45383), .ZN(W45463));
  INVX1 G38877 (.I(I1076), .ZN(W5461));
  INVX1 G38878 (.I(I1401), .ZN(W5465));
  INVX1 G38879 (.I(W3887), .ZN(W5466));
  INVX1 G38880 (.I(I809), .ZN(O14734));
  INVX1 G38881 (.I(W4176), .ZN(W6096));
  INVX1 G38882 (.I(W29134), .ZN(O14728));
  INVX1 G38883 (.I(W13896), .ZN(O14727));
  INVX1 G38884 (.I(W2070), .ZN(W5477));
  INVX1 G38885 (.I(W3264), .ZN(W5479));
  INVX1 G38886 (.I(W31425), .ZN(O14724));
  INVX1 G38887 (.I(W1393), .ZN(W5481));
  INVX1 G38888 (.I(W861), .ZN(W5482));
  INVX1 G38889 (.I(W38203), .ZN(O14721));
  INVX1 G38890 (.I(W40), .ZN(W6692));
  INVX1 G38891 (.I(W605), .ZN(W6682));
  INVX1 G38892 (.I(I1468), .ZN(O13732));
  INVX1 G38893 (.I(W4854), .ZN(W6684));
  INVX1 G38894 (.I(W37737), .ZN(W44226));
  INVX1 G38895 (.I(W5227), .ZN(W6686));
  INVX1 G38896 (.I(W3907), .ZN(O13728));
  INVX1 G38897 (.I(W1482), .ZN(W6688));
  INVX1 G38898 (.I(W4581), .ZN(W6690));
  INVX1 G38899 (.I(W5859), .ZN(W6691));
  INVX1 G38900 (.I(W5088), .ZN(W6681));
  INVX1 G38901 (.I(W897), .ZN(O13723));
  INVX1 G38902 (.I(W12993), .ZN(O13722));
  INVX1 G38903 (.I(W22746), .ZN(O13721));
  INVX1 G38904 (.I(W6207), .ZN(W6698));
  INVX1 G38905 (.I(I1856), .ZN(W6700));
  INVX1 G38906 (.I(W24446), .ZN(O13716));
  INVX1 G38907 (.I(W22336), .ZN(W44209));
  INVX1 G38908 (.I(I819), .ZN(W6702));
  INVX1 G38909 (.I(W104), .ZN(W6675));
  INVX1 G38910 (.I(W16886), .ZN(O13749));
  INVX1 G38911 (.I(W6639), .ZN(O13748));
  INVX1 G38912 (.I(W1429), .ZN(O13747));
  INVX1 G38913 (.I(W30009), .ZN(O13746));
  INVX1 G38914 (.I(W32003), .ZN(W44249));
  INVX1 G38915 (.I(W1936), .ZN(W6671));
  INVX1 G38916 (.I(W23029), .ZN(W44246));
  INVX1 G38917 (.I(W6261), .ZN(W6673));
  INVX1 G38918 (.I(W2685), .ZN(W6674));
  INVX1 G38919 (.I(W13606), .ZN(O13712));
  INVX1 G38920 (.I(W37603), .ZN(O13741));
  INVX1 G38921 (.I(W356), .ZN(W44241));
  INVX1 G38922 (.I(W3219), .ZN(W44239));
  INVX1 G38923 (.I(W5497), .ZN(O13738));
  INVX1 G38924 (.I(W27821), .ZN(O13737));
  INVX1 G38925 (.I(W5246), .ZN(O13736));
  INVX1 G38926 (.I(W5253), .ZN(W6680));
  INVX1 G38927 (.I(W3076), .ZN(O13734));
  INVX1 G38928 (.I(I108), .ZN(W6743));
  INVX1 G38929 (.I(W18138), .ZN(O13688));
  INVX1 G38930 (.I(W17187), .ZN(O13687));
  INVX1 G38931 (.I(W25667), .ZN(O13685));
  INVX1 G38932 (.I(W4118), .ZN(O13683));
  INVX1 G38933 (.I(W580), .ZN(W6740));
  INVX1 G38934 (.I(W15482), .ZN(W44167));
  INVX1 G38935 (.I(W1894), .ZN(W6741));
  INVX1 G38936 (.I(I1421), .ZN(O13680));
  INVX1 G38937 (.I(W41287), .ZN(O13679));
  INVX1 G38938 (.I(W32183), .ZN(O13689));
  INVX1 G38939 (.I(W2671), .ZN(W6744));
  INVX1 G38940 (.I(I908), .ZN(W44159));
  INVX1 G38941 (.I(W236), .ZN(O13677));
  INVX1 G38942 (.I(W427), .ZN(W6751));
  INVX1 G38943 (.I(W29662), .ZN(W44154));
  INVX1 G38944 (.I(W28573), .ZN(W44153));
  INVX1 G38945 (.I(W39286), .ZN(O13674));
  INVX1 G38946 (.I(I676), .ZN(W6754));
  INVX1 G38947 (.I(W3944), .ZN(W6720));
  INVX1 G38948 (.I(W6641), .ZN(W6706));
  INVX1 G38949 (.I(I1985), .ZN(O143));
  INVX1 G38950 (.I(W40683), .ZN(O13706));
  INVX1 G38951 (.I(W5916), .ZN(W6712));
  INVX1 G38952 (.I(W33066), .ZN(O13702));
  INVX1 G38953 (.I(W6801), .ZN(O13701));
  INVX1 G38954 (.I(I856), .ZN(W6715));
  INVX1 G38955 (.I(W5531), .ZN(W6716));
  INVX1 G38956 (.I(W3275), .ZN(O13750));
  INVX1 G38957 (.I(W40986), .ZN(W44190));
  INVX1 G38958 (.I(W8208), .ZN(O13697));
  INVX1 G38959 (.I(I54), .ZN(O13696));
  INVX1 G38960 (.I(W2486), .ZN(W6721));
  INVX1 G38961 (.I(I605), .ZN(O147));
  INVX1 G38962 (.I(W21144), .ZN(W44183));
  INVX1 G38963 (.I(I1853), .ZN(W6726));
  INVX1 G38964 (.I(W40169), .ZN(O13690));
  INVX1 G38965 (.I(W24665), .ZN(O13802));
  INVX1 G38966 (.I(I1080), .ZN(O13811));
  INVX1 G38967 (.I(W6450), .ZN(O13810));
  INVX1 G38968 (.I(W9660), .ZN(O13809));
  INVX1 G38969 (.I(W14505), .ZN(O13808));
  INVX1 G38970 (.I(W380), .ZN(W6607));
  INVX1 G38971 (.I(I537), .ZN(W6609));
  INVX1 G38972 (.I(W857), .ZN(W6610));
  INVX1 G38973 (.I(W26377), .ZN(O13804));
  INVX1 G38974 (.I(W38772), .ZN(O13803));
  INVX1 G38975 (.I(W5785), .ZN(O138));
  INVX1 G38976 (.I(W4242), .ZN(W6611));
  INVX1 G38977 (.I(I836), .ZN(W6612));
  INVX1 G38978 (.I(I1684), .ZN(W6613));
  INVX1 G38979 (.I(W89), .ZN(W6620));
  INVX1 G38980 (.I(W35374), .ZN(O13796));
  INVX1 G38981 (.I(W30100), .ZN(O13794));
  INVX1 G38982 (.I(W6803), .ZN(O13792));
  INVX1 G38983 (.I(W13259), .ZN(O13791));
  INVX1 G38984 (.I(W4458), .ZN(W6587));
  INVX1 G38985 (.I(W19014), .ZN(O13833));
  INVX1 G38986 (.I(W5069), .ZN(W6579));
  INVX1 G38987 (.I(W24990), .ZN(W44348));
  INVX1 G38988 (.I(W40276), .ZN(O13830));
  INVX1 G38989 (.I(W32597), .ZN(O13829));
  INVX1 G38990 (.I(W5692), .ZN(W6581));
  INVX1 G38991 (.I(W3254), .ZN(W6583));
  INVX1 G38992 (.I(I554), .ZN(W6584));
  INVX1 G38993 (.I(W979), .ZN(W6585));
  INVX1 G38994 (.I(W30729), .ZN(O13790));
  INVX1 G38995 (.I(W1261), .ZN(W6588));
  INVX1 G38996 (.I(I208), .ZN(W6591));
  INVX1 G38997 (.I(I541), .ZN(W6593));
  INVX1 G38998 (.I(W16698), .ZN(O13819));
  INVX1 G38999 (.I(W1638), .ZN(W6596));
  INVX1 G39000 (.I(W16611), .ZN(O13816));
  INVX1 G39001 (.I(W6352), .ZN(W6598));
  INVX1 G39002 (.I(W431), .ZN(W6599));
  INVX1 G39003 (.I(W2623), .ZN(W6663));
  INVX1 G39004 (.I(W373), .ZN(W6658));
  INVX1 G39005 (.I(W15362), .ZN(O13767));
  INVX1 G39006 (.I(W41242), .ZN(O13766));
  INVX1 G39007 (.I(W22), .ZN(O13765));
  INVX1 G39008 (.I(W20116), .ZN(O13763));
  INVX1 G39009 (.I(W20735), .ZN(O13761));
  INVX1 G39010 (.I(I1156), .ZN(W6662));
  INVX1 G39011 (.I(W11354), .ZN(O13759));
  INVX1 G39012 (.I(W8078), .ZN(O13758));
  INVX1 G39013 (.I(I278), .ZN(W6656));
  INVX1 G39014 (.I(W4811), .ZN(W6664));
  INVX1 G39015 (.I(W4143), .ZN(W6665));
  INVX1 G39016 (.I(W26402), .ZN(W44261));
  INVX1 G39017 (.I(W4319), .ZN(W6667));
  INVX1 G39018 (.I(W7931), .ZN(O13754));
  INVX1 G39019 (.I(W37930), .ZN(O13752));
  INVX1 G39020 (.I(W7632), .ZN(O13751));
  INVX1 G39021 (.I(W214), .ZN(W6670));
  INVX1 G39022 (.I(W42006), .ZN(O13781));
  INVX1 G39023 (.I(W8454), .ZN(O13789));
  INVX1 G39024 (.I(I1589), .ZN(W6631));
  INVX1 G39025 (.I(W1575), .ZN(W6639));
  INVX1 G39026 (.I(W15849), .ZN(W44296));
  INVX1 G39027 (.I(W7195), .ZN(O13784));
  INVX1 G39028 (.I(W42901), .ZN(W44293));
  INVX1 G39029 (.I(W14551), .ZN(W44292));
  INVX1 G39030 (.I(W38899), .ZN(O13782));
  INVX1 G39031 (.I(I669), .ZN(W6755));
  INVX1 G39032 (.I(I1538), .ZN(W6645));
  INVX1 G39033 (.I(W5642), .ZN(W6648));
  INVX1 G39034 (.I(W3076), .ZN(O13778));
  INVX1 G39035 (.I(I697), .ZN(W6650));
  INVX1 G39036 (.I(W25169), .ZN(O13776));
  INVX1 G39037 (.I(W13227), .ZN(O13774));
  INVX1 G39038 (.I(W42419), .ZN(O13773));
  INVX1 G39039 (.I(I1563), .ZN(W6655));
  INVX1 G39040 (.I(W256), .ZN(W6922));
  INVX1 G39041 (.I(W1259), .ZN(W6909));
  INVX1 G39042 (.I(W31500), .ZN(O13551));
  INVX1 G39043 (.I(W520), .ZN(W6913));
  INVX1 G39044 (.I(I1952), .ZN(O13548));
  INVX1 G39045 (.I(W2515), .ZN(W6916));
  INVX1 G39046 (.I(I938), .ZN(W43992));
  INVX1 G39047 (.I(W19957), .ZN(O13544));
  INVX1 G39048 (.I(I294), .ZN(O13543));
  INVX1 G39049 (.I(W3887), .ZN(W6921));
  INVX1 G39050 (.I(W34685), .ZN(O13554));
  INVX1 G39051 (.I(W6415), .ZN(W6925));
  INVX1 G39052 (.I(W14049), .ZN(O13540));
  INVX1 G39053 (.I(W2717), .ZN(W6926));
  INVX1 G39054 (.I(W1762), .ZN(W6928));
  INVX1 G39055 (.I(W442), .ZN(W6929));
  INVX1 G39056 (.I(W2307), .ZN(W6931));
  INVX1 G39057 (.I(W1486), .ZN(W6932));
  INVX1 G39058 (.I(W39880), .ZN(O13534));
  INVX1 G39059 (.I(W30328), .ZN(O13566));
  INVX1 G39060 (.I(I1090), .ZN(W6872));
  INVX1 G39061 (.I(W1343), .ZN(W6876));
  INVX1 G39062 (.I(W795), .ZN(O155));
  INVX1 G39063 (.I(W2702), .ZN(W6885));
  INVX1 G39064 (.I(W31727), .ZN(W44024));
  INVX1 G39065 (.I(W18180), .ZN(W44023));
  INVX1 G39066 (.I(W12014), .ZN(O13570));
  INVX1 G39067 (.I(W34799), .ZN(O13568));
  INVX1 G39068 (.I(W8031), .ZN(O13567));
  INVX1 G39069 (.I(W38539), .ZN(W43976));
  INVX1 G39070 (.I(W8539), .ZN(O13564));
  INVX1 G39071 (.I(W6708), .ZN(W6896));
  INVX1 G39072 (.I(W5507), .ZN(W6898));
  INVX1 G39073 (.I(W904), .ZN(W6900));
  INVX1 G39074 (.I(W291), .ZN(W6902));
  INVX1 G39075 (.I(W513), .ZN(W6906));
  INVX1 G39076 (.I(W27376), .ZN(W44004));
  INVX1 G39077 (.I(W21479), .ZN(O13555));
  INVX1 G39078 (.I(W3263), .ZN(W6967));
  INVX1 G39079 (.I(W23108), .ZN(W43947));
  INVX1 G39080 (.I(W31700), .ZN(O13509));
  INVX1 G39081 (.I(W29237), .ZN(O13507));
  INVX1 G39082 (.I(W6638), .ZN(W6960));
  INVX1 G39083 (.I(I1442), .ZN(O158));
  INVX1 G39084 (.I(W38695), .ZN(O13503));
  INVX1 G39085 (.I(W24651), .ZN(O13502));
  INVX1 G39086 (.I(W1360), .ZN(W6966));
  INVX1 G39087 (.I(W8450), .ZN(O13500));
  INVX1 G39088 (.I(W18199), .ZN(O13510));
  INVX1 G39089 (.I(W3111), .ZN(W6968));
  INVX1 G39090 (.I(W1134), .ZN(W6972));
  INVX1 G39091 (.I(I1758), .ZN(W6976));
  INVX1 G39092 (.I(W2142), .ZN(W6977));
  INVX1 G39093 (.I(W38939), .ZN(O13494));
  INVX1 G39094 (.I(W14636), .ZN(O13493));
  INVX1 G39095 (.I(W42364), .ZN(O13491));
  INVX1 G39096 (.I(W27055), .ZN(O13490));
  INVX1 G39097 (.I(W33014), .ZN(O13520));
  INVX1 G39098 (.I(W2434), .ZN(W6933));
  INVX1 G39099 (.I(W25351), .ZN(O13532));
  INVX1 G39100 (.I(I1658), .ZN(W6937));
  INVX1 G39101 (.I(I488), .ZN(W6942));
  INVX1 G39102 (.I(W4947), .ZN(W6943));
  INVX1 G39103 (.I(I635), .ZN(W6944));
  INVX1 G39104 (.I(W13524), .ZN(O13522));
  INVX1 G39105 (.I(I315), .ZN(W6950));
  INVX1 G39106 (.I(W135), .ZN(W6871));
  INVX1 G39107 (.I(W27652), .ZN(O13519));
  INVX1 G39108 (.I(W5441), .ZN(W6951));
  INVX1 G39109 (.I(W3732), .ZN(W43958));
  INVX1 G39110 (.I(W6295), .ZN(W6955));
  INVX1 G39111 (.I(W40996), .ZN(O13514));
  INVX1 G39112 (.I(W17776), .ZN(O13513));
  INVX1 G39113 (.I(W1708), .ZN(W6956));
  INVX1 G39114 (.I(W32160), .ZN(W43950));
  INVX1 G39115 (.I(W35269), .ZN(O13639));
  INVX1 G39116 (.I(W33715), .ZN(O13650));
  INVX1 G39117 (.I(W3098), .ZN(W44120));
  INVX1 G39118 (.I(I443), .ZN(W6790));
  INVX1 G39119 (.I(W3551), .ZN(W6793));
  INVX1 G39120 (.I(W29200), .ZN(O13646));
  INVX1 G39121 (.I(W5390), .ZN(O13645));
  INVX1 G39122 (.I(W33276), .ZN(O13643));
  INVX1 G39123 (.I(W28468), .ZN(O13641));
  INVX1 G39124 (.I(W7190), .ZN(O13640));
  INVX1 G39125 (.I(W3807), .ZN(W6787));
  INVX1 G39126 (.I(W6413), .ZN(W6799));
  INVX1 G39127 (.I(W21477), .ZN(O13636));
  INVX1 G39128 (.I(W34032), .ZN(O13635));
  INVX1 G39129 (.I(W1261), .ZN(W6807));
  INVX1 G39130 (.I(W30705), .ZN(O13631));
  INVX1 G39131 (.I(I797), .ZN(W6808));
  INVX1 G39132 (.I(W2674), .ZN(W6810));
  INVX1 G39133 (.I(W4025), .ZN(W6811));
  INVX1 G39134 (.I(W1672), .ZN(W6770));
  INVX1 G39135 (.I(W630), .ZN(O13672));
  INVX1 G39136 (.I(I839), .ZN(O13671));
  INVX1 G39137 (.I(W5075), .ZN(W6758));
  INVX1 G39138 (.I(W121), .ZN(W6759));
  INVX1 G39139 (.I(W3567), .ZN(O13667));
  INVX1 G39140 (.I(W1830), .ZN(W6761));
  INVX1 G39141 (.I(W358), .ZN(W6762));
  INVX1 G39142 (.I(W21175), .ZN(W44139));
  INVX1 G39143 (.I(W11966), .ZN(O13663));
  INVX1 G39144 (.I(W233), .ZN(W6812));
  INVX1 G39145 (.I(W4884), .ZN(W6771));
  INVX1 G39146 (.I(W5743), .ZN(W6774));
  INVX1 G39147 (.I(W5739), .ZN(W44132));
  INVX1 G39148 (.I(I1523), .ZN(W6776));
  INVX1 G39149 (.I(W3168), .ZN(W6777));
  INVX1 G39150 (.I(I904), .ZN(W6778));
  INVX1 G39151 (.I(W16185), .ZN(O13655));
  INVX1 G39152 (.I(W5742), .ZN(W6786));
  INVX1 G39153 (.I(W134), .ZN(W6846));
  INVX1 G39154 (.I(W4413), .ZN(W6835));
  INVX1 G39155 (.I(W31844), .ZN(O13605));
  INVX1 G39156 (.I(W2530), .ZN(W6837));
  INVX1 G39157 (.I(W18030), .ZN(W44064));
  INVX1 G39158 (.I(W4538), .ZN(W6839));
  INVX1 G39159 (.I(W36350), .ZN(O13601));
  INVX1 G39160 (.I(W21351), .ZN(O13599));
  INVX1 G39161 (.I(W42334), .ZN(O13598));
  INVX1 G39162 (.I(W11173), .ZN(O13596));
  INVX1 G39163 (.I(W5879), .ZN(W6833));
  INVX1 G39164 (.I(W4129), .ZN(W6849));
  INVX1 G39165 (.I(W631), .ZN(O13591));
  INVX1 G39166 (.I(W1531), .ZN(W6858));
  INVX1 G39167 (.I(W28236), .ZN(O13588));
  INVX1 G39168 (.I(W6236), .ZN(W6860));
  INVX1 G39169 (.I(W5901), .ZN(O13586));
  INVX1 G39170 (.I(W28345), .ZN(O13583));
  INVX1 G39171 (.I(W10832), .ZN(O13581));
  INVX1 G39172 (.I(I1430), .ZN(W6828));
  INVX1 G39173 (.I(W262), .ZN(W6815));
  INVX1 G39174 (.I(W5146), .ZN(W6819));
  INVX1 G39175 (.I(I1621), .ZN(W6820));
  INVX1 G39176 (.I(W3097), .ZN(W6822));
  INVX1 G39177 (.I(I1794), .ZN(W6823));
  INVX1 G39178 (.I(W10665), .ZN(O13620));
  INVX1 G39179 (.I(W1493), .ZN(W6826));
  INVX1 G39180 (.I(W4239), .ZN(W6827));
  INVX1 G39181 (.I(W39294), .ZN(O13835));
  INVX1 G39182 (.I(W40889), .ZN(O13616));
  INVX1 G39183 (.I(W24537), .ZN(W44077));
  INVX1 G39184 (.I(W22442), .ZN(W44075));
  INVX1 G39185 (.I(W21536), .ZN(O13612));
  INVX1 G39186 (.I(W28199), .ZN(O13611));
  INVX1 G39187 (.I(W38704), .ZN(O13610));
  INVX1 G39188 (.I(W1290), .ZN(W6832));
  INVX1 G39189 (.I(W8934), .ZN(O13609));
  INVX1 G39190 (.I(W4649), .ZN(W6251));
  INVX1 G39191 (.I(W13880), .ZN(W44682));
  INVX1 G39192 (.I(W1874), .ZN(W6244));
  INVX1 G39193 (.I(W24862), .ZN(W44680));
  INVX1 G39194 (.I(W16770), .ZN(O14103));
  INVX1 G39195 (.I(W3662), .ZN(W6248));
  INVX1 G39196 (.I(W3254), .ZN(O14099));
  INVX1 G39197 (.I(W5355), .ZN(O14098));
  INVX1 G39198 (.I(W3060), .ZN(W6250));
  INVX1 G39199 (.I(W14727), .ZN(O14095));
  INVX1 G39200 (.I(W4416), .ZN(W6242));
  INVX1 G39201 (.I(I319), .ZN(W6252));
  INVX1 G39202 (.I(W20528), .ZN(W44668));
  INVX1 G39203 (.I(W5228), .ZN(O14092));
  INVX1 G39204 (.I(W36435), .ZN(O14091));
  INVX1 G39205 (.I(W4583), .ZN(W6258));
  INVX1 G39206 (.I(W39771), .ZN(O14089));
  INVX1 G39207 (.I(W20237), .ZN(O14088));
  INVX1 G39208 (.I(W40664), .ZN(O14087));
  INVX1 G39209 (.I(W3902), .ZN(W6227));
  INVX1 G39210 (.I(W15833), .ZN(O14131));
  INVX1 G39211 (.I(W5076), .ZN(W6203));
  INVX1 G39212 (.I(W5849), .ZN(W6210));
  INVX1 G39213 (.I(W16187), .ZN(O14125));
  INVX1 G39214 (.I(I1355), .ZN(O123));
  INVX1 G39215 (.I(W1780), .ZN(W6216));
  INVX1 G39216 (.I(W1652), .ZN(W6220));
  INVX1 G39217 (.I(W22542), .ZN(O14119));
  INVX1 G39218 (.I(W11338), .ZN(O14117));
  INVX1 G39219 (.I(W4788), .ZN(W6259));
  INVX1 G39220 (.I(W21661), .ZN(W44698));
  INVX1 G39221 (.I(W5760), .ZN(W6228));
  INVX1 G39222 (.I(W17621), .ZN(O14114));
  INVX1 G39223 (.I(W4837), .ZN(W44694));
  INVX1 G39224 (.I(I744), .ZN(W6233));
  INVX1 G39225 (.I(W12776), .ZN(O14108));
  INVX1 G39226 (.I(W3000), .ZN(W6238));
  INVX1 G39227 (.I(I817), .ZN(W6240));
  INVX1 G39228 (.I(W26715), .ZN(O14047));
  INVX1 G39229 (.I(W291), .ZN(W6279));
  INVX1 G39230 (.I(W21508), .ZN(O14062));
  INVX1 G39231 (.I(W1696), .ZN(W6285));
  INVX1 G39232 (.I(W37859), .ZN(O14057));
  INVX1 G39233 (.I(W3165), .ZN(W6287));
  INVX1 G39234 (.I(W3530), .ZN(W6294));
  INVX1 G39235 (.I(W1229), .ZN(W6296));
  INVX1 G39236 (.I(W33839), .ZN(O14049));
  INVX1 G39237 (.I(W3797), .ZN(W6298));
  INVX1 G39238 (.I(I1164), .ZN(W6278));
  INVX1 G39239 (.I(W4274), .ZN(O127));
  INVX1 G39240 (.I(W3136), .ZN(W6301));
  INVX1 G39241 (.I(W2496), .ZN(W6302));
  INVX1 G39242 (.I(W31), .ZN(W6304));
  INVX1 G39243 (.I(W2119), .ZN(W6305));
  INVX1 G39244 (.I(W11316), .ZN(W44603));
  INVX1 G39245 (.I(W2028), .ZN(W6311));
  INVX1 G39246 (.I(I842), .ZN(W6312));
  INVX1 G39247 (.I(W4690), .ZN(W6268));
  INVX1 G39248 (.I(W37094), .ZN(W44655));
  INVX1 G39249 (.I(W5793), .ZN(W6260));
  INVX1 G39250 (.I(W26407), .ZN(O14085));
  INVX1 G39251 (.I(W39010), .ZN(O14082));
  INVX1 G39252 (.I(I444), .ZN(W6266));
  INVX1 G39253 (.I(W3482), .ZN(W44647));
  INVX1 G39254 (.I(W39680), .ZN(W44646));
  INVX1 G39255 (.I(W36654), .ZN(W44645));
  INVX1 G39256 (.I(W27840), .ZN(O14132));
  INVX1 G39257 (.I(W3438), .ZN(W6270));
  INVX1 G39258 (.I(I1301), .ZN(W6272));
  INVX1 G39259 (.I(W3745), .ZN(W6273));
  INVX1 G39260 (.I(W21277), .ZN(O14073));
  INVX1 G39261 (.I(W14738), .ZN(O14072));
  INVX1 G39262 (.I(W1707), .ZN(O14071));
  INVX1 G39263 (.I(W15363), .ZN(O14070));
  INVX1 G39264 (.I(W2926), .ZN(O14066));
  INVX1 G39265 (.I(W3490), .ZN(W6133));
  INVX1 G39266 (.I(W2383), .ZN(W6120));
  INVX1 G39267 (.I(I50), .ZN(O14201));
  INVX1 G39268 (.I(W11442), .ZN(O14200));
  INVX1 G39269 (.I(W11755), .ZN(O14197));
  INVX1 G39270 (.I(W2407), .ZN(W6126));
  INVX1 G39271 (.I(W1106), .ZN(W6131));
  INVX1 G39272 (.I(W39263), .ZN(O14193));
  INVX1 G39273 (.I(W27674), .ZN(O14192));
  INVX1 G39274 (.I(W39864), .ZN(O14190));
  INVX1 G39275 (.I(W3206), .ZN(W6116));
  INVX1 G39276 (.I(W4280), .ZN(W6134));
  INVX1 G39277 (.I(W44702), .ZN(O14187));
  INVX1 G39278 (.I(W1983), .ZN(W6137));
  INVX1 G39279 (.I(W32086), .ZN(O14186));
  INVX1 G39280 (.I(W852), .ZN(W6142));
  INVX1 G39281 (.I(W1627), .ZN(W6151));
  INVX1 G39282 (.I(I1116), .ZN(W6154));
  INVX1 G39283 (.I(W3723), .ZN(W6156));
  INVX1 G39284 (.I(W2967), .ZN(W6109));
  INVX1 G39285 (.I(I1588), .ZN(W6100));
  INVX1 G39286 (.I(W8517), .ZN(O14220));
  INVX1 G39287 (.I(W1322), .ZN(W6101));
  INVX1 G39288 (.I(W2749), .ZN(W6103));
  INVX1 G39289 (.I(W25291), .ZN(O14217));
  INVX1 G39290 (.I(W34537), .ZN(O14215));
  INVX1 G39291 (.I(W15240), .ZN(O14214));
  INVX1 G39292 (.I(W42239), .ZN(W44824));
  INVX1 G39293 (.I(W5159), .ZN(W6106));
  INVX1 G39294 (.I(I1807), .ZN(W6159));
  INVX1 G39295 (.I(W43646), .ZN(O14211));
  INVX1 G39296 (.I(W23648), .ZN(O14210));
  INVX1 G39297 (.I(W2074), .ZN(W6110));
  INVX1 G39298 (.I(W7182), .ZN(W44816));
  INVX1 G39299 (.I(W1809), .ZN(W6111));
  INVX1 G39300 (.I(I285), .ZN(W6113));
  INVX1 G39301 (.I(W6862), .ZN(O14207));
  INVX1 G39302 (.I(W6198), .ZN(W44812));
  INVX1 G39303 (.I(W8256), .ZN(O14145));
  INVX1 G39304 (.I(W11885), .ZN(O14156));
  INVX1 G39305 (.I(W23912), .ZN(O14155));
  INVX1 G39306 (.I(W2213), .ZN(O122));
  INVX1 G39307 (.I(W32782), .ZN(O14150));
  INVX1 G39308 (.I(W2057), .ZN(W6195));
  INVX1 G39309 (.I(W3095), .ZN(O14148));
  INVX1 G39310 (.I(W40488), .ZN(O14147));
  INVX1 G39311 (.I(W10136), .ZN(O14146));
  INVX1 G39312 (.I(W8380), .ZN(W44735));
  INVX1 G39313 (.I(W37522), .ZN(O14157));
  INVX1 G39314 (.I(W7695), .ZN(O14144));
  INVX1 G39315 (.I(W43276), .ZN(O14141));
  INVX1 G39316 (.I(W13852), .ZN(O14140));
  INVX1 G39317 (.I(W40179), .ZN(O14139));
  INVX1 G39318 (.I(I1892), .ZN(O14136));
  INVX1 G39319 (.I(W3862), .ZN(W6201));
  INVX1 G39320 (.I(W2359), .ZN(W6202));
  INVX1 G39321 (.I(W24007), .ZN(O14133));
  INVX1 G39322 (.I(W23506), .ZN(W44763));
  INVX1 G39323 (.I(W18616), .ZN(O14175));
  INVX1 G39324 (.I(W572), .ZN(W6164));
  INVX1 G39325 (.I(W2434), .ZN(W6167));
  INVX1 G39326 (.I(W33494), .ZN(O14173));
  INVX1 G39327 (.I(W3347), .ZN(W6170));
  INVX1 G39328 (.I(W5988), .ZN(O14170));
  INVX1 G39329 (.I(I1870), .ZN(W6172));
  INVX1 G39330 (.I(W41462), .ZN(O14167));
  INVX1 G39331 (.I(I163), .ZN(W6313));
  INVX1 G39332 (.I(W29893), .ZN(W44762));
  INVX1 G39333 (.I(W3100), .ZN(W6177));
  INVX1 G39334 (.I(W10748), .ZN(O14164));
  INVX1 G39335 (.I(I583), .ZN(O14163));
  INVX1 G39336 (.I(W6293), .ZN(O14161));
  INVX1 G39337 (.I(W2085), .ZN(W6182));
  INVX1 G39338 (.I(W14516), .ZN(O14159));
  INVX1 G39339 (.I(W1642), .ZN(W6187));
  INVX1 G39340 (.I(W5011), .ZN(O13896));
  INVX1 G39341 (.I(W20537), .ZN(O13908));
  INVX1 G39342 (.I(I1547), .ZN(W6481));
  INVX1 G39343 (.I(W2107), .ZN(W44441));
  INVX1 G39344 (.I(W4125), .ZN(W6484));
  INVX1 G39345 (.I(W13724), .ZN(O13904));
  INVX1 G39346 (.I(W5100), .ZN(O13903));
  INVX1 G39347 (.I(W27), .ZN(W6488));
  INVX1 G39348 (.I(W11798), .ZN(O13899));
  INVX1 G39349 (.I(W4686), .ZN(W6490));
  INVX1 G39350 (.I(W5809), .ZN(W6480));
  INVX1 G39351 (.I(I1465), .ZN(W6491));
  INVX1 G39352 (.I(W33070), .ZN(O13893));
  INVX1 G39353 (.I(W4843), .ZN(W6497));
  INVX1 G39354 (.I(W16393), .ZN(O13889));
  INVX1 G39355 (.I(W13915), .ZN(O13888));
  INVX1 G39356 (.I(W33473), .ZN(O13887));
  INVX1 G39357 (.I(W687), .ZN(O13886));
  INVX1 G39358 (.I(W4641), .ZN(W6499));
  INVX1 G39359 (.I(I896), .ZN(W6458));
  INVX1 G39360 (.I(W4306), .ZN(W6442));
  INVX1 G39361 (.I(W11138), .ZN(W44474));
  INVX1 G39362 (.I(W4444), .ZN(W6445));
  INVX1 G39363 (.I(W1228), .ZN(W6446));
  INVX1 G39364 (.I(I316), .ZN(W6448));
  INVX1 G39365 (.I(W3332), .ZN(W6451));
  INVX1 G39366 (.I(W18), .ZN(W6452));
  INVX1 G39367 (.I(W31398), .ZN(O13929));
  INVX1 G39368 (.I(W3106), .ZN(W6454));
  INVX1 G39369 (.I(W15396), .ZN(O13883));
  INVX1 G39370 (.I(W31098), .ZN(O13925));
  INVX1 G39371 (.I(I380), .ZN(O13920));
  INVX1 G39372 (.I(W26050), .ZN(O13919));
  INVX1 G39373 (.I(W20969), .ZN(O13918));
  INVX1 G39374 (.I(W6315), .ZN(W6467));
  INVX1 G39375 (.I(W6839), .ZN(O13916));
  INVX1 G39376 (.I(W43002), .ZN(O13915));
  INVX1 G39377 (.I(I554), .ZN(W6476));
  INVX1 G39378 (.I(W9685), .ZN(O13849));
  INVX1 G39379 (.I(W2113), .ZN(W6526));
  INVX1 G39380 (.I(I909), .ZN(W6527));
  INVX1 G39381 (.I(I1320), .ZN(W44384));
  INVX1 G39382 (.I(W2910), .ZN(O13859));
  INVX1 G39383 (.I(W7629), .ZN(O13858));
  INVX1 G39384 (.I(W6164), .ZN(W6536));
  INVX1 G39385 (.I(W4875), .ZN(W6540));
  INVX1 G39386 (.I(I1197), .ZN(W6552));
  INVX1 G39387 (.I(W5208), .ZN(W6555));
  INVX1 G39388 (.I(W2942), .ZN(W6524));
  INVX1 G39389 (.I(W1582), .ZN(O13845));
  INVX1 G39390 (.I(W28258), .ZN(O13844));
  INVX1 G39391 (.I(W6002), .ZN(W6566));
  INVX1 G39392 (.I(I1818), .ZN(W6567));
  INVX1 G39393 (.I(W31184), .ZN(O13840));
  INVX1 G39394 (.I(W5597), .ZN(W44359));
  INVX1 G39395 (.I(W476), .ZN(W6570));
  INVX1 G39396 (.I(W5082), .ZN(O13836));
  INVX1 G39397 (.I(W10483), .ZN(O13873));
  INVX1 G39398 (.I(W5577), .ZN(O13882));
  INVX1 G39399 (.I(W6014), .ZN(W6501));
  INVX1 G39400 (.I(W11535), .ZN(O13881));
  INVX1 G39401 (.I(W41763), .ZN(O13880));
  INVX1 G39402 (.I(W32213), .ZN(O13879));
  INVX1 G39403 (.I(W31998), .ZN(O13878));
  INVX1 G39404 (.I(W1539), .ZN(O13876));
  INVX1 G39405 (.I(W1264), .ZN(W6509));
  INVX1 G39406 (.I(W15135), .ZN(O13937));
  INVX1 G39407 (.I(W3918), .ZN(O13871));
  INVX1 G39408 (.I(W5560), .ZN(O13870));
  INVX1 G39409 (.I(W1303), .ZN(W6515));
  INVX1 G39410 (.I(W31350), .ZN(O13868));
  INVX1 G39411 (.I(W5482), .ZN(W6517));
  INVX1 G39412 (.I(W3166), .ZN(W6519));
  INVX1 G39413 (.I(W3689), .ZN(W6520));
  INVX1 G39414 (.I(W40945), .ZN(O13863));
  INVX1 G39415 (.I(I235), .ZN(W6365));
  INVX1 G39416 (.I(I1816), .ZN(W6351));
  INVX1 G39417 (.I(W33657), .ZN(W44561));
  INVX1 G39418 (.I(W5187), .ZN(W6352));
  INVX1 G39419 (.I(W25891), .ZN(O14005));
  INVX1 G39420 (.I(W4667), .ZN(W6356));
  INVX1 G39421 (.I(W4483), .ZN(W6358));
  INVX1 G39422 (.I(W18208), .ZN(O14000));
  INVX1 G39423 (.I(W2411), .ZN(W6364));
  INVX1 G39424 (.I(W20310), .ZN(O13998));
  INVX1 G39425 (.I(W23484), .ZN(O14008));
  INVX1 G39426 (.I(W1496), .ZN(O13996));
  INVX1 G39427 (.I(I1366), .ZN(W6367));
  INVX1 G39428 (.I(W30932), .ZN(O13994));
  INVX1 G39429 (.I(W594), .ZN(W6369));
  INVX1 G39430 (.I(W10121), .ZN(W44545));
  INVX1 G39431 (.I(I676), .ZN(O13992));
  INVX1 G39432 (.I(W23815), .ZN(O13991));
  INVX1 G39433 (.I(W324), .ZN(W6371));
  INVX1 G39434 (.I(I1665), .ZN(W6334));
  INVX1 G39435 (.I(W39431), .ZN(O14035));
  INVX1 G39436 (.I(W2667), .ZN(O14034));
  INVX1 G39437 (.I(W12144), .ZN(O14030));
  INVX1 G39438 (.I(W43889), .ZN(W44590));
  INVX1 G39439 (.I(W917), .ZN(W6326));
  INVX1 G39440 (.I(W3293), .ZN(O14026));
  INVX1 G39441 (.I(I18), .ZN(W6330));
  INVX1 G39442 (.I(W40529), .ZN(W44581));
  INVX1 G39443 (.I(I1983), .ZN(W6333));
  INVX1 G39444 (.I(W5729), .ZN(W6372));
  INVX1 G39445 (.I(W3486), .ZN(W6336));
  INVX1 G39446 (.I(I370), .ZN(O14018));
  INVX1 G39447 (.I(W3142), .ZN(W6339));
  INVX1 G39448 (.I(W5077), .ZN(W6341));
  INVX1 G39449 (.I(I858), .ZN(W6343));
  INVX1 G39450 (.I(W4971), .ZN(W6344));
  INVX1 G39451 (.I(W8645), .ZN(O14012));
  INVX1 G39452 (.I(W15610), .ZN(O14011));
  INVX1 G39453 (.I(W3039), .ZN(W6414));
  INVX1 G39454 (.I(W31166), .ZN(O13967));
  INVX1 G39455 (.I(W15778), .ZN(O13966));
  INVX1 G39456 (.I(W1246), .ZN(W6405));
  INVX1 G39457 (.I(W4421), .ZN(O13963));
  INVX1 G39458 (.I(W2213), .ZN(W6407));
  INVX1 G39459 (.I(W693), .ZN(W6409));
  INVX1 G39460 (.I(W13745), .ZN(O13960));
  INVX1 G39461 (.I(W15281), .ZN(W44504));
  INVX1 G39462 (.I(W15562), .ZN(O13956));
  INVX1 G39463 (.I(W4733), .ZN(W6401));
  INVX1 G39464 (.I(W33153), .ZN(O13954));
  INVX1 G39465 (.I(W7830), .ZN(O13951));
  INVX1 G39466 (.I(I1322), .ZN(W6422));
  INVX1 G39467 (.I(I1718), .ZN(W6430));
  INVX1 G39468 (.I(W32881), .ZN(W44486));
  INVX1 G39469 (.I(W1279), .ZN(W6433));
  INVX1 G39470 (.I(W5618), .ZN(O13941));
  INVX1 G39471 (.I(W9456), .ZN(O13939));
  INVX1 G39472 (.I(W3341), .ZN(W6388));
  INVX1 G39473 (.I(W5867), .ZN(W6373));
  INVX1 G39474 (.I(W4775), .ZN(W6374));
  INVX1 G39475 (.I(W10843), .ZN(O13986));
  INVX1 G39476 (.I(W24941), .ZN(O13985));
  INVX1 G39477 (.I(W30468), .ZN(O13983));
  INVX1 G39478 (.I(I164), .ZN(W6381));
  INVX1 G39479 (.I(W16185), .ZN(W44531));
  INVX1 G39480 (.I(W26160), .ZN(O13980));
  INVX1 G39481 (.I(W233), .ZN(W5211));
  INVX1 G39482 (.I(W3105), .ZN(O13978));
  INVX1 G39483 (.I(I1278), .ZN(W6389));
  INVX1 G39484 (.I(I778), .ZN(O129));
  INVX1 G39485 (.I(W40421), .ZN(O13975));
  INVX1 G39486 (.I(W701), .ZN(W6397));
  INVX1 G39487 (.I(W31740), .ZN(O13971));
  INVX1 G39488 (.I(W1262), .ZN(O13970));
  INVX1 G39489 (.I(I1726), .ZN(W6399));
  INVX1 G39490 (.I(W36372), .ZN(O15909));
  INVX1 G39491 (.I(W2691), .ZN(W4083));
  INVX1 G39492 (.I(W2548), .ZN(W4086));
  INVX1 G39493 (.I(I1913), .ZN(W4087));
  INVX1 G39494 (.I(W3108), .ZN(W4088));
  INVX1 G39495 (.I(I410), .ZN(W4092));
  INVX1 G39496 (.I(W44703), .ZN(O15918));
  INVX1 G39497 (.I(W1812), .ZN(W4096));
  INVX1 G39498 (.I(W81), .ZN(W4097));
  INVX1 G39499 (.I(I1054), .ZN(W4102));
  INVX1 G39500 (.I(W14339), .ZN(O15924));
  INVX1 G39501 (.I(W2615), .ZN(W4106));
  INVX1 G39502 (.I(W13733), .ZN(O15907));
  INVX1 G39503 (.I(W2345), .ZN(W4109));
  INVX1 G39504 (.I(W14069), .ZN(W46867));
  INVX1 G39505 (.I(W1866), .ZN(W4112));
  INVX1 G39506 (.I(W2994), .ZN(W4114));
  INVX1 G39507 (.I(W17903), .ZN(O15902));
  INVX1 G39508 (.I(W3558), .ZN(W4115));
  INVX1 G39509 (.I(W5465), .ZN(O15934));
  INVX1 G39510 (.I(W1289), .ZN(W4053));
  INVX1 G39511 (.I(W46473), .ZN(O15947));
  INVX1 G39512 (.I(W16193), .ZN(W46914));
  INVX1 G39513 (.I(W33757), .ZN(O15946));
  INVX1 G39514 (.I(W7890), .ZN(O15945));
  INVX1 G39515 (.I(W163), .ZN(W4060));
  INVX1 G39516 (.I(W3479), .ZN(W4061));
  INVX1 G39517 (.I(W3409), .ZN(W4064));
  INVX1 G39518 (.I(W2641), .ZN(W4071));
  INVX1 G39519 (.I(W3145), .ZN(W4116));
  INVX1 G39520 (.I(W3216), .ZN(W4075));
  INVX1 G39521 (.I(W11877), .ZN(O15931));
  INVX1 G39522 (.I(W2565), .ZN(O15929));
  INVX1 G39523 (.I(I1466), .ZN(W4079));
  INVX1 G39524 (.I(W755), .ZN(W4080));
  INVX1 G39525 (.I(W16393), .ZN(O15927));
  INVX1 G39526 (.I(W8803), .ZN(O15926));
  INVX1 G39527 (.I(W2391), .ZN(W4082));
  INVX1 G39528 (.I(W18618), .ZN(O15866));
  INVX1 G39529 (.I(W46203), .ZN(O15879));
  INVX1 G39530 (.I(W740), .ZN(W4144));
  INVX1 G39531 (.I(I626), .ZN(W4147));
  INVX1 G39532 (.I(W2217), .ZN(W4148));
  INVX1 G39533 (.I(W2765), .ZN(W4150));
  INVX1 G39534 (.I(W2538), .ZN(W4154));
  INVX1 G39535 (.I(W1438), .ZN(O15872));
  INVX1 G39536 (.I(W2132), .ZN(W4158));
  INVX1 G39537 (.I(W9090), .ZN(O15867));
  INVX1 G39538 (.I(W129), .ZN(W4142));
  INVX1 G39539 (.I(I1801), .ZN(W4166));
  INVX1 G39540 (.I(W8431), .ZN(W46814));
  INVX1 G39541 (.I(W1943), .ZN(W4169));
  INVX1 G39542 (.I(W3597), .ZN(W4170));
  INVX1 G39543 (.I(W3199), .ZN(W4171));
  INVX1 G39544 (.I(W1294), .ZN(W4172));
  INVX1 G39545 (.I(W35839), .ZN(O15861));
  INVX1 G39546 (.I(W45925), .ZN(O15859));
  INVX1 G39547 (.I(W790), .ZN(W4125));
  INVX1 G39548 (.I(W2029), .ZN(W46860));
  INVX1 G39549 (.I(W27626), .ZN(O15899));
  INVX1 G39550 (.I(W10219), .ZN(W46858));
  INVX1 G39551 (.I(W41744), .ZN(O15898));
  INVX1 G39552 (.I(W37785), .ZN(O15897));
  INVX1 G39553 (.I(W1754), .ZN(W4117));
  INVX1 G39554 (.I(W2605), .ZN(W4118));
  INVX1 G39555 (.I(W9410), .ZN(W46852));
  INVX1 G39556 (.I(W9443), .ZN(O15892));
  INVX1 G39557 (.I(W1795), .ZN(W4052));
  INVX1 G39558 (.I(W4), .ZN(W4126));
  INVX1 G39559 (.I(I635), .ZN(W4132));
  INVX1 G39560 (.I(W42302), .ZN(O15887));
  INVX1 G39561 (.I(W25583), .ZN(O15885));
  INVX1 G39562 (.I(W35027), .ZN(W46841));
  INVX1 G39563 (.I(W2204), .ZN(W4136));
  INVX1 G39564 (.I(W28715), .ZN(W46836));
  INVX1 G39565 (.I(I1578), .ZN(W4139));
  INVX1 G39566 (.I(W1748), .ZN(W3987));
  INVX1 G39567 (.I(W591), .ZN(W3980));
  INVX1 G39568 (.I(W2525), .ZN(W3982));
  INVX1 G39569 (.I(W19911), .ZN(O16011));
  INVX1 G39570 (.I(W40052), .ZN(O16010));
  INVX1 G39571 (.I(I404), .ZN(W3983));
  INVX1 G39572 (.I(I1440), .ZN(W3985));
  INVX1 G39573 (.I(I870), .ZN(W3986));
  INVX1 G39574 (.I(W43638), .ZN(O16007));
  INVX1 G39575 (.I(W32622), .ZN(O16006));
  INVX1 G39576 (.I(W438), .ZN(O16016));
  INVX1 G39577 (.I(W1815), .ZN(W3988));
  INVX1 G39578 (.I(W102), .ZN(W3991));
  INVX1 G39579 (.I(W103), .ZN(W3993));
  INVX1 G39580 (.I(I1883), .ZN(W3996));
  INVX1 G39581 (.I(I1158), .ZN(W3998));
  INVX1 G39582 (.I(I1678), .ZN(O15998));
  INVX1 G39583 (.I(W2225), .ZN(W4000));
  INVX1 G39584 (.I(W7076), .ZN(O15997));
  INVX1 G39585 (.I(W12051), .ZN(W47010));
  INVX1 G39586 (.I(W43832), .ZN(O16035));
  INVX1 G39587 (.I(W10723), .ZN(O16034));
  INVX1 G39588 (.I(I1095), .ZN(W3958));
  INVX1 G39589 (.I(W41452), .ZN(O16032));
  INVX1 G39590 (.I(W2626), .ZN(W3959));
  INVX1 G39591 (.I(W3760), .ZN(O16030));
  INVX1 G39592 (.I(I467), .ZN(O50));
  INVX1 G39593 (.I(W9278), .ZN(O16028));
  INVX1 G39594 (.I(W42580), .ZN(O16027));
  INVX1 G39595 (.I(W3702), .ZN(W4001));
  INVX1 G39596 (.I(W28769), .ZN(W47008));
  INVX1 G39597 (.I(I1488), .ZN(W3963));
  INVX1 G39598 (.I(I1793), .ZN(W3966));
  INVX1 G39599 (.I(W3226), .ZN(W3967));
  INVX1 G39600 (.I(W1406), .ZN(W3970));
  INVX1 G39601 (.I(W1847), .ZN(W3971));
  INVX1 G39602 (.I(W1664), .ZN(W3973));
  INVX1 G39603 (.I(I741), .ZN(O16017));
  INVX1 G39604 (.I(W626), .ZN(W4030));
  INVX1 G39605 (.I(W789), .ZN(W4017));
  INVX1 G39606 (.I(W1211), .ZN(W4019));
  INVX1 G39607 (.I(W3306), .ZN(W4020));
  INVX1 G39608 (.I(I673), .ZN(W4022));
  INVX1 G39609 (.I(W16318), .ZN(O15974));
  INVX1 G39610 (.I(W3315), .ZN(W4024));
  INVX1 G39611 (.I(W15643), .ZN(O15971));
  INVX1 G39612 (.I(W29600), .ZN(O15970));
  INVX1 G39613 (.I(W10255), .ZN(O15966));
  INVX1 G39614 (.I(W240), .ZN(W4015));
  INVX1 G39615 (.I(W20494), .ZN(O15961));
  INVX1 G39616 (.I(W2194), .ZN(W4039));
  INVX1 G39617 (.I(W1556), .ZN(W4040));
  INVX1 G39618 (.I(I525), .ZN(W4041));
  INVX1 G39619 (.I(I1561), .ZN(W4043));
  INVX1 G39620 (.I(W1932), .ZN(W4045));
  INVX1 G39621 (.I(W781), .ZN(W4049));
  INVX1 G39622 (.I(W1787), .ZN(W4051));
  INVX1 G39623 (.I(W44926), .ZN(O15990));
  INVX1 G39624 (.I(W2762), .ZN(W4002));
  INVX1 G39625 (.I(W41003), .ZN(O15994));
  INVX1 G39626 (.I(I1957), .ZN(W4004));
  INVX1 G39627 (.I(W42824), .ZN(W46968));
  INVX1 G39628 (.I(W44868), .ZN(O15993));
  INVX1 G39629 (.I(W1346), .ZN(W4005));
  INVX1 G39630 (.I(I526), .ZN(O15992));
  INVX1 G39631 (.I(I1194), .ZN(W4006));
  INVX1 G39632 (.I(W1072), .ZN(O52));
  INVX1 G39633 (.I(W18348), .ZN(O15989));
  INVX1 G39634 (.I(W13710), .ZN(O15988));
  INVX1 G39635 (.I(I966), .ZN(W4009));
  INVX1 G39636 (.I(W45988), .ZN(O15985));
  INVX1 G39637 (.I(W2687), .ZN(W4010));
  INVX1 G39638 (.I(W3545), .ZN(W4011));
  INVX1 G39639 (.I(W14330), .ZN(O15982));
  INVX1 G39640 (.I(W18652), .ZN(O15979));
  INVX1 G39641 (.I(W1070), .ZN(W4340));
  INVX1 G39642 (.I(W13845), .ZN(O15741));
  INVX1 G39643 (.I(W13374), .ZN(O15740));
  INVX1 G39644 (.I(W46176), .ZN(O15738));
  INVX1 G39645 (.I(W391), .ZN(W4330));
  INVX1 G39646 (.I(W11967), .ZN(O15736));
  INVX1 G39647 (.I(W1329), .ZN(W4336));
  INVX1 G39648 (.I(W35265), .ZN(W46660));
  INVX1 G39649 (.I(W4874), .ZN(O15734));
  INVX1 G39650 (.I(W18481), .ZN(O15732));
  INVX1 G39651 (.I(W988), .ZN(W4325));
  INVX1 G39652 (.I(W28365), .ZN(O15729));
  INVX1 G39653 (.I(W18740), .ZN(O15725));
  INVX1 G39654 (.I(W44456), .ZN(O15724));
  INVX1 G39655 (.I(I1303), .ZN(W4351));
  INVX1 G39656 (.I(W3315), .ZN(W4352));
  INVX1 G39657 (.I(W2670), .ZN(W4355));
  INVX1 G39658 (.I(I1950), .ZN(O15719));
  INVX1 G39659 (.I(W35670), .ZN(O15718));
  INVX1 G39660 (.I(W45964), .ZN(O15756));
  INVX1 G39661 (.I(W14725), .ZN(O15765));
  INVX1 G39662 (.I(W3177), .ZN(W4297));
  INVX1 G39663 (.I(W1905), .ZN(W4300));
  INVX1 G39664 (.I(W36132), .ZN(O15762));
  INVX1 G39665 (.I(W15538), .ZN(O15761));
  INVX1 G39666 (.I(W4196), .ZN(W4306));
  INVX1 G39667 (.I(W36037), .ZN(O15759));
  INVX1 G39668 (.I(W1654), .ZN(W4310));
  INVX1 G39669 (.I(W41392), .ZN(W46686));
  INVX1 G39670 (.I(W276), .ZN(W4357));
  INVX1 G39671 (.I(W3762), .ZN(W4311));
  INVX1 G39672 (.I(I1445), .ZN(W4312));
  INVX1 G39673 (.I(W27972), .ZN(W46681));
  INVX1 G39674 (.I(W3921), .ZN(W4317));
  INVX1 G39675 (.I(W2511), .ZN(O55));
  INVX1 G39676 (.I(W2932), .ZN(W4320));
  INVX1 G39677 (.I(W19869), .ZN(O15747));
  INVX1 G39678 (.I(I207), .ZN(W4322));
  INVX1 G39679 (.I(I371), .ZN(O57));
  INVX1 G39680 (.I(W2056), .ZN(W4405));
  INVX1 G39681 (.I(W3796), .ZN(W4406));
  INVX1 G39682 (.I(W5937), .ZN(O15688));
  INVX1 G39683 (.I(I1193), .ZN(W4407));
  INVX1 G39684 (.I(W4299), .ZN(W4411));
  INVX1 G39685 (.I(W14928), .ZN(O15684));
  INVX1 G39686 (.I(W24160), .ZN(O15683));
  INVX1 G39687 (.I(W27994), .ZN(O15682));
  INVX1 G39688 (.I(W21083), .ZN(O15681));
  INVX1 G39689 (.I(W2412), .ZN(W4401));
  INVX1 G39690 (.I(W12242), .ZN(O15680));
  INVX1 G39691 (.I(I912), .ZN(W4416));
  INVX1 G39692 (.I(I58), .ZN(W4417));
  INVX1 G39693 (.I(W4076), .ZN(W4418));
  INVX1 G39694 (.I(I1940), .ZN(W4419));
  INVX1 G39695 (.I(W12799), .ZN(O15673));
  INVX1 G39696 (.I(I1402), .ZN(W4425));
  INVX1 G39697 (.I(W1758), .ZN(W4426));
  INVX1 G39698 (.I(W1486), .ZN(W4378));
  INVX1 G39699 (.I(W475), .ZN(W4358));
  INVX1 G39700 (.I(W41714), .ZN(O15716));
  INVX1 G39701 (.I(I1016), .ZN(W4360));
  INVX1 G39702 (.I(W1833), .ZN(W4362));
  INVX1 G39703 (.I(W1657), .ZN(W4365));
  INVX1 G39704 (.I(W1245), .ZN(W4368));
  INVX1 G39705 (.I(W2154), .ZN(W4373));
  INVX1 G39706 (.I(W425), .ZN(W4375));
  INVX1 G39707 (.I(W3667), .ZN(W4296));
  INVX1 G39708 (.I(W22264), .ZN(O15701));
  INVX1 G39709 (.I(W1481), .ZN(W4389));
  INVX1 G39710 (.I(I772), .ZN(W46617));
  INVX1 G39711 (.I(W2249), .ZN(O15698));
  INVX1 G39712 (.I(W1218), .ZN(W4396));
  INVX1 G39713 (.I(W44901), .ZN(O15696));
  INVX1 G39714 (.I(W2662), .ZN(W4398));
  INVX1 G39715 (.I(W4254), .ZN(W4399));
  INVX1 G39716 (.I(W14340), .ZN(O15822));
  INVX1 G39717 (.I(I252), .ZN(W4210));
  INVX1 G39718 (.I(W1824), .ZN(W4211));
  INVX1 G39719 (.I(W30924), .ZN(W46776));
  INVX1 G39720 (.I(W2048), .ZN(W4213));
  INVX1 G39721 (.I(I276), .ZN(W4215));
  INVX1 G39722 (.I(I879), .ZN(W4216));
  INVX1 G39723 (.I(W19023), .ZN(W46769));
  INVX1 G39724 (.I(W3202), .ZN(W4221));
  INVX1 G39725 (.I(W1225), .ZN(W4224));
  INVX1 G39726 (.I(W34623), .ZN(O15834));
  INVX1 G39727 (.I(I804), .ZN(W4229));
  INVX1 G39728 (.I(W460), .ZN(W4231));
  INVX1 G39729 (.I(I1273), .ZN(W4235));
  INVX1 G39730 (.I(W1124), .ZN(W4237));
  INVX1 G39731 (.I(W3884), .ZN(W4238));
  INVX1 G39732 (.I(W12900), .ZN(O15817));
  INVX1 G39733 (.I(I1306), .ZN(O15816));
  INVX1 G39734 (.I(W3517), .ZN(W4239));
  INVX1 G39735 (.I(W3759), .ZN(W4204));
  INVX1 G39736 (.I(W23903), .ZN(O15856));
  INVX1 G39737 (.I(W1859), .ZN(W4184));
  INVX1 G39738 (.I(W32168), .ZN(O15853));
  INVX1 G39739 (.I(W185), .ZN(W4185));
  INVX1 G39740 (.I(W3841), .ZN(W4186));
  INVX1 G39741 (.I(W3654), .ZN(W4187));
  INVX1 G39742 (.I(W212), .ZN(W4190));
  INVX1 G39743 (.I(W3855), .ZN(W4198));
  INVX1 G39744 (.I(W2909), .ZN(W4199));
  INVX1 G39745 (.I(W38253), .ZN(O15814));
  INVX1 G39746 (.I(W5330), .ZN(O15845));
  INVX1 G39747 (.I(I853), .ZN(O15843));
  INVX1 G39748 (.I(I684), .ZN(O15842));
  INVX1 G39749 (.I(W27637), .ZN(O15840));
  INVX1 G39750 (.I(W5775), .ZN(O15839));
  INVX1 G39751 (.I(W30372), .ZN(O15838));
  INVX1 G39752 (.I(W33942), .ZN(O15836));
  INVX1 G39753 (.I(W27595), .ZN(O15835));
  INVX1 G39754 (.I(W546), .ZN(W4274));
  INVX1 G39755 (.I(W1448), .ZN(W4262));
  INVX1 G39756 (.I(W1197), .ZN(W4263));
  INVX1 G39757 (.I(W34079), .ZN(O15789));
  INVX1 G39758 (.I(W3433), .ZN(W4266));
  INVX1 G39759 (.I(W2051), .ZN(W4267));
  INVX1 G39760 (.I(I239), .ZN(W4271));
  INVX1 G39761 (.I(W9724), .ZN(O15782));
  INVX1 G39762 (.I(W4222), .ZN(W4272));
  INVX1 G39763 (.I(W1374), .ZN(W4273));
  INVX1 G39764 (.I(W33354), .ZN(O15796));
  INVX1 G39765 (.I(W15927), .ZN(O15779));
  INVX1 G39766 (.I(W34487), .ZN(W46709));
  INVX1 G39767 (.I(W19290), .ZN(W46708));
  INVX1 G39768 (.I(W1580), .ZN(W4279));
  INVX1 G39769 (.I(W497), .ZN(W4291));
  INVX1 G39770 (.I(W137), .ZN(W4295));
  INVX1 G39771 (.I(I1418), .ZN(O15768));
  INVX1 G39772 (.I(W14059), .ZN(O15767));
  INVX1 G39773 (.I(W462), .ZN(O15805));
  INVX1 G39774 (.I(W6063), .ZN(O15813));
  INVX1 G39775 (.I(W37354), .ZN(W46754));
  INVX1 G39776 (.I(W1073), .ZN(W4240));
  INVX1 G39777 (.I(W3271), .ZN(W4241));
  INVX1 G39778 (.I(W32948), .ZN(O15811));
  INVX1 G39779 (.I(W3743), .ZN(W4243));
  INVX1 G39780 (.I(W25574), .ZN(O15808));
  INVX1 G39781 (.I(W17976), .ZN(O15807));
  INVX1 G39782 (.I(W9838), .ZN(O16040));
  INVX1 G39783 (.I(W14301), .ZN(O15804));
  INVX1 G39784 (.I(W35065), .ZN(O15803));
  INVX1 G39785 (.I(W2024), .ZN(W4249));
  INVX1 G39786 (.I(W15509), .ZN(O15800));
  INVX1 G39787 (.I(W16393), .ZN(O15799));
  INVX1 G39788 (.I(W3853), .ZN(W4250));
  INVX1 G39789 (.I(W1715), .ZN(W4254));
  INVX1 G39790 (.I(W3153), .ZN(W4255));
  INVX1 G39791 (.I(I773), .ZN(W3675));
  INVX1 G39792 (.I(I521), .ZN(W3665));
  INVX1 G39793 (.I(W15282), .ZN(O16298));
  INVX1 G39794 (.I(I1620), .ZN(W3668));
  INVX1 G39795 (.I(W19160), .ZN(O16294));
  INVX1 G39796 (.I(W2656), .ZN(W3669));
  INVX1 G39797 (.I(W729), .ZN(W47309));
  INVX1 G39798 (.I(W46815), .ZN(W47308));
  INVX1 G39799 (.I(I1380), .ZN(W3670));
  INVX1 G39800 (.I(I614), .ZN(W3672));
  INVX1 G39801 (.I(W1515), .ZN(W3657));
  INVX1 G39802 (.I(I1018), .ZN(O16287));
  INVX1 G39803 (.I(W29955), .ZN(O16286));
  INVX1 G39804 (.I(W1193), .ZN(O16285));
  INVX1 G39805 (.I(I924), .ZN(W3676));
  INVX1 G39806 (.I(W3368), .ZN(O16283));
  INVX1 G39807 (.I(W40681), .ZN(W47296));
  INVX1 G39808 (.I(W9598), .ZN(O16282));
  INVX1 G39809 (.I(W369), .ZN(W3678));
  INVX1 G39810 (.I(W20338), .ZN(O16312));
  INVX1 G39811 (.I(W22667), .ZN(O16322));
  INVX1 G39812 (.I(I551), .ZN(O16321));
  INVX1 G39813 (.I(W556), .ZN(O16320));
  INVX1 G39814 (.I(W3331), .ZN(W3637));
  INVX1 G39815 (.I(W46215), .ZN(O16319));
  INVX1 G39816 (.I(W368), .ZN(W3641));
  INVX1 G39817 (.I(W219), .ZN(W3648));
  INVX1 G39818 (.I(W2646), .ZN(O16314));
  INVX1 G39819 (.I(W29032), .ZN(O16313));
  INVX1 G39820 (.I(W615), .ZN(W3679));
  INVX1 G39821 (.I(W894), .ZN(W3649));
  INVX1 G39822 (.I(W33132), .ZN(O16310));
  INVX1 G39823 (.I(W1255), .ZN(O16309));
  INVX1 G39824 (.I(I445), .ZN(W3650));
  INVX1 G39825 (.I(W29896), .ZN(O16307));
  INVX1 G39826 (.I(W8790), .ZN(O16306));
  INVX1 G39827 (.I(W39127), .ZN(O16305));
  INVX1 G39828 (.I(W3089), .ZN(W3656));
  INVX1 G39829 (.I(W329), .ZN(W3719));
  INVX1 G39830 (.I(W23358), .ZN(O16258));
  INVX1 G39831 (.I(W2586), .ZN(W3705));
  INVX1 G39832 (.I(W30715), .ZN(O16257));
  INVX1 G39833 (.I(W231), .ZN(W3706));
  INVX1 G39834 (.I(W5378), .ZN(O16255));
  INVX1 G39835 (.I(W25504), .ZN(O16253));
  INVX1 G39836 (.I(W2045), .ZN(W3713));
  INVX1 G39837 (.I(W23678), .ZN(O16252));
  INVX1 G39838 (.I(W30802), .ZN(O16250));
  INVX1 G39839 (.I(W17662), .ZN(O16260));
  INVX1 G39840 (.I(I512), .ZN(W3720));
  INVX1 G39841 (.I(W45249), .ZN(O16244));
  INVX1 G39842 (.I(W24549), .ZN(O16243));
  INVX1 G39843 (.I(W2068), .ZN(W3726));
  INVX1 G39844 (.I(I1513), .ZN(O16241));
  INVX1 G39845 (.I(W15243), .ZN(O16240));
  INVX1 G39846 (.I(W40317), .ZN(O16239));
  INVX1 G39847 (.I(I455), .ZN(W3729));
  INVX1 G39848 (.I(W1530), .ZN(O16273));
  INVX1 G39849 (.I(I191), .ZN(W3680));
  INVX1 G39850 (.I(I16), .ZN(W3681));
  INVX1 G39851 (.I(W1868), .ZN(W3682));
  INVX1 G39852 (.I(W3171), .ZN(W3683));
  INVX1 G39853 (.I(I263), .ZN(W3685));
  INVX1 G39854 (.I(W29506), .ZN(W47287));
  INVX1 G39855 (.I(W2607), .ZN(W3687));
  INVX1 G39856 (.I(I1809), .ZN(W3689));
  INVX1 G39857 (.I(I720), .ZN(W3631));
  INVX1 G39858 (.I(W1356), .ZN(W3690));
  INVX1 G39859 (.I(W27955), .ZN(O16271));
  INVX1 G39860 (.I(W2453), .ZN(W3691));
  INVX1 G39861 (.I(W2757), .ZN(W3692));
  INVX1 G39862 (.I(W17133), .ZN(O16265));
  INVX1 G39863 (.I(W2264), .ZN(W3698));
  INVX1 G39864 (.I(W14229), .ZN(O16262));
  INVX1 G39865 (.I(W1072), .ZN(W3702));
  INVX1 G39866 (.I(I1629), .ZN(W3573));
  INVX1 G39867 (.I(W1616), .ZN(W3563));
  INVX1 G39868 (.I(W3377), .ZN(O16386));
  INVX1 G39869 (.I(W2154), .ZN(W3564));
  INVX1 G39870 (.I(W5009), .ZN(O16385));
  INVX1 G39871 (.I(W2963), .ZN(W3570));
  INVX1 G39872 (.I(W2860), .ZN(O16380));
  INVX1 G39873 (.I(W424), .ZN(W3572));
  INVX1 G39874 (.I(I1737), .ZN(O16378));
  INVX1 G39875 (.I(W31540), .ZN(O16377));
  INVX1 G39876 (.I(W100), .ZN(W3562));
  INVX1 G39877 (.I(W12589), .ZN(O16376));
  INVX1 G39878 (.I(W45678), .ZN(O16375));
  INVX1 G39879 (.I(W3888), .ZN(O16374));
  INVX1 G39880 (.I(I743), .ZN(W3579));
  INVX1 G39881 (.I(W46748), .ZN(O16371));
  INVX1 G39882 (.I(W1035), .ZN(W3580));
  INVX1 G39883 (.I(W5006), .ZN(O16369));
  INVX1 G39884 (.I(W3088), .ZN(W3586));
  INVX1 G39885 (.I(W1797), .ZN(W3545));
  INVX1 G39886 (.I(I784), .ZN(W3526));
  INVX1 G39887 (.I(W1659), .ZN(O38));
  INVX1 G39888 (.I(W13601), .ZN(O16413));
  INVX1 G39889 (.I(W2166), .ZN(W3533));
  INVX1 G39890 (.I(I1619), .ZN(W3534));
  INVX1 G39891 (.I(I75), .ZN(W3540));
  INVX1 G39892 (.I(W51), .ZN(W3542));
  INVX1 G39893 (.I(W9138), .ZN(O16403));
  INVX1 G39894 (.I(W1786), .ZN(W3543));
  INVX1 G39895 (.I(W7544), .ZN(O16365));
  INVX1 G39896 (.I(W2669), .ZN(W3548));
  INVX1 G39897 (.I(I1810), .ZN(W3551));
  INVX1 G39898 (.I(W3504), .ZN(W3554));
  INVX1 G39899 (.I(I1416), .ZN(W3557));
  INVX1 G39900 (.I(W35877), .ZN(O16392));
  INVX1 G39901 (.I(W17310), .ZN(O16391));
  INVX1 G39902 (.I(W25813), .ZN(O16390));
  INVX1 G39903 (.I(W627), .ZN(W3561));
  INVX1 G39904 (.I(W62), .ZN(W3620));
  INVX1 G39905 (.I(W4290), .ZN(O16347));
  INVX1 G39906 (.I(I1396), .ZN(W3609));
  INVX1 G39907 (.I(W14961), .ZN(O16345));
  INVX1 G39908 (.I(I518), .ZN(W3611));
  INVX1 G39909 (.I(I1333), .ZN(W3612));
  INVX1 G39910 (.I(W6357), .ZN(O16342));
  INVX1 G39911 (.I(W44364), .ZN(O16340));
  INVX1 G39912 (.I(W10148), .ZN(O16338));
  INVX1 G39913 (.I(W2907), .ZN(W3618));
  INVX1 G39914 (.I(W22415), .ZN(O16348));
  INVX1 G39915 (.I(W15905), .ZN(O16333));
  INVX1 G39916 (.I(W24004), .ZN(O16332));
  INVX1 G39917 (.I(W1617), .ZN(W3624));
  INVX1 G39918 (.I(W1572), .ZN(W3626));
  INVX1 G39919 (.I(W26183), .ZN(O16329));
  INVX1 G39920 (.I(W1235), .ZN(W3627));
  INVX1 G39921 (.I(W24844), .ZN(O16327));
  INVX1 G39922 (.I(W1544), .ZN(W3628));
  INVX1 G39923 (.I(W43692), .ZN(W47381));
  INVX1 G39924 (.I(W17835), .ZN(O16364));
  INVX1 G39925 (.I(W43910), .ZN(O16363));
  INVX1 G39926 (.I(W25197), .ZN(O16362));
  INVX1 G39927 (.I(W29494), .ZN(W47388));
  INVX1 G39928 (.I(W39771), .ZN(W47385));
  INVX1 G39929 (.I(W42199), .ZN(W47384));
  INVX1 G39930 (.I(I222), .ZN(W3593));
  INVX1 G39931 (.I(W36635), .ZN(O16359));
  INVX1 G39932 (.I(W38220), .ZN(O16236));
  INVX1 G39933 (.I(W23569), .ZN(O16357));
  INVX1 G39934 (.I(I904), .ZN(W3597));
  INVX1 G39935 (.I(W3446), .ZN(W3598));
  INVX1 G39936 (.I(I1968), .ZN(W3599));
  INVX1 G39937 (.I(W450), .ZN(W3601));
  INVX1 G39938 (.I(I150), .ZN(W3603));
  INVX1 G39939 (.I(W26), .ZN(W3606));
  INVX1 G39940 (.I(W46210), .ZN(O16349));
  INVX1 G39941 (.I(W1876), .ZN(W3863));
  INVX1 G39942 (.I(I1638), .ZN(W3851));
  INVX1 G39943 (.I(W40114), .ZN(O16114));
  INVX1 G39944 (.I(W31984), .ZN(W47105));
  INVX1 G39945 (.I(I1325), .ZN(W3854));
  INVX1 G39946 (.I(W8355), .ZN(O16112));
  INVX1 G39947 (.I(W3276), .ZN(W3855));
  INVX1 G39948 (.I(W382), .ZN(W3862));
  INVX1 G39949 (.I(W34117), .ZN(O16107));
  INVX1 G39950 (.I(W14050), .ZN(O16106));
  INVX1 G39951 (.I(W213), .ZN(O47));
  INVX1 G39952 (.I(W3277), .ZN(W3865));
  INVX1 G39953 (.I(W3009), .ZN(W3871));
  INVX1 G39954 (.I(W45467), .ZN(W47090));
  INVX1 G39955 (.I(W1764), .ZN(W3872));
  INVX1 G39956 (.I(W2684), .ZN(W3874));
  INVX1 G39957 (.I(W2263), .ZN(W3883));
  INVX1 G39958 (.I(W253), .ZN(W3884));
  INVX1 G39959 (.I(W2413), .ZN(O16092));
  INVX1 G39960 (.I(W39042), .ZN(O16126));
  INVX1 G39961 (.I(W2450), .ZN(W3835));
  INVX1 G39962 (.I(W1245), .ZN(W3837));
  INVX1 G39963 (.I(W1498), .ZN(W3839));
  INVX1 G39964 (.I(W44336), .ZN(O16131));
  INVX1 G39965 (.I(W3473), .ZN(W3840));
  INVX1 G39966 (.I(W35686), .ZN(O16129));
  INVX1 G39967 (.I(W34717), .ZN(W47122));
  INVX1 G39968 (.I(W20141), .ZN(O16127));
  INVX1 G39969 (.I(W817), .ZN(W47120));
  INVX1 G39970 (.I(W3513), .ZN(W3891));
  INVX1 G39971 (.I(W17482), .ZN(O16125));
  INVX1 G39972 (.I(W42889), .ZN(W47117));
  INVX1 G39973 (.I(W2241), .ZN(W3845));
  INVX1 G39974 (.I(W1804), .ZN(W3846));
  INVX1 G39975 (.I(W42187), .ZN(O16121));
  INVX1 G39976 (.I(W43631), .ZN(O16120));
  INVX1 G39977 (.I(W3111), .ZN(W3847));
  INVX1 G39978 (.I(W45262), .ZN(O16118));
  INVX1 G39979 (.I(W2635), .ZN(W3925));
  INVX1 G39980 (.I(I1333), .ZN(W3913));
  INVX1 G39981 (.I(W22641), .ZN(O16066));
  INVX1 G39982 (.I(W2378), .ZN(O16065));
  INVX1 G39983 (.I(W3535), .ZN(O16062));
  INVX1 G39984 (.I(W321), .ZN(W3918));
  INVX1 G39985 (.I(W18310), .ZN(O16060));
  INVX1 G39986 (.I(W2868), .ZN(W3919));
  INVX1 G39987 (.I(W10), .ZN(W3922));
  INVX1 G39988 (.I(W34686), .ZN(O16056));
  INVX1 G39989 (.I(W44667), .ZN(O16069));
  INVX1 G39990 (.I(W2769), .ZN(W3931));
  INVX1 G39991 (.I(W1692), .ZN(W3932));
  INVX1 G39992 (.I(I1980), .ZN(W3933));
  INVX1 G39993 (.I(I1712), .ZN(W3935));
  INVX1 G39994 (.I(W164), .ZN(W3940));
  INVX1 G39995 (.I(I1184), .ZN(W3944));
  INVX1 G39996 (.I(W23029), .ZN(W47027));
  INVX1 G39997 (.I(W32089), .ZN(O16042));
  INVX1 G39998 (.I(W1760), .ZN(W3898));
  INVX1 G39999 (.I(W2027), .ZN(W3892));
  INVX1 G40000 (.I(W6623), .ZN(O16089));
  INVX1 G40001 (.I(W812), .ZN(W3893));
  INVX1 G40002 (.I(W24828), .ZN(O16087));
  INVX1 G40003 (.I(W35375), .ZN(O16086));
  INVX1 G40004 (.I(W40789), .ZN(O16085));
  INVX1 G40005 (.I(W447), .ZN(W3896));
  INVX1 G40006 (.I(W39990), .ZN(O16082));
  INVX1 G40007 (.I(W2555), .ZN(W3833));
  INVX1 G40008 (.I(W2506), .ZN(W3899));
  INVX1 G40009 (.I(W1529), .ZN(W3900));
  INVX1 G40010 (.I(W2959), .ZN(W3905));
  INVX1 G40011 (.I(W24781), .ZN(O16075));
  INVX1 G40012 (.I(W27406), .ZN(O16074));
  INVX1 G40013 (.I(W994), .ZN(W3908));
  INVX1 G40014 (.I(W25233), .ZN(W47057));
  INVX1 G40015 (.I(W1040), .ZN(W3910));
  INVX1 G40016 (.I(I1020), .ZN(W3773));
  INVX1 G40017 (.I(I568), .ZN(W3761));
  INVX1 G40018 (.I(W42771), .ZN(O16207));
  INVX1 G40019 (.I(W2500), .ZN(W3764));
  INVX1 G40020 (.I(W19903), .ZN(O16201));
  INVX1 G40021 (.I(W36772), .ZN(O16197));
  INVX1 G40022 (.I(W26044), .ZN(O16196));
  INVX1 G40023 (.I(W43387), .ZN(O16195));
  INVX1 G40024 (.I(W291), .ZN(W3771));
  INVX1 G40025 (.I(W5352), .ZN(W47195));
  INVX1 G40026 (.I(I1461), .ZN(W3760));
  INVX1 G40027 (.I(W3233), .ZN(W3774));
  INVX1 G40028 (.I(W37267), .ZN(O16190));
  INVX1 G40029 (.I(W19094), .ZN(O16189));
  INVX1 G40030 (.I(W3386), .ZN(O16188));
  INVX1 G40031 (.I(I78), .ZN(W3775));
  INVX1 G40032 (.I(I1389), .ZN(W3781));
  INVX1 G40033 (.I(W593), .ZN(W3782));
  INVX1 G40034 (.I(W43291), .ZN(O16183));
  INVX1 G40035 (.I(I564), .ZN(W3750));
  INVX1 G40036 (.I(I1626), .ZN(W3730));
  INVX1 G40037 (.I(W2217), .ZN(W3732));
  INVX1 G40038 (.I(W1658), .ZN(W3733));
  INVX1 G40039 (.I(W20902), .ZN(O16232));
  INVX1 G40040 (.I(W1578), .ZN(W3736));
  INVX1 G40041 (.I(W11884), .ZN(O16229));
  INVX1 G40042 (.I(I1488), .ZN(W3740));
  INVX1 G40043 (.I(W1096), .ZN(W3745));
  INVX1 G40044 (.I(W1096), .ZN(W47227));
  INVX1 G40045 (.I(W1270), .ZN(W3786));
  INVX1 G40046 (.I(W35293), .ZN(O16218));
  INVX1 G40047 (.I(W1853), .ZN(O16217));
  INVX1 G40048 (.I(I172), .ZN(W3751));
  INVX1 G40049 (.I(W3374), .ZN(W3754));
  INVX1 G40050 (.I(W23008), .ZN(O16213));
  INVX1 G40051 (.I(W19008), .ZN(W47216));
  INVX1 G40052 (.I(W949), .ZN(W3757));
  INVX1 G40053 (.I(W32278), .ZN(O16211));
  INVX1 G40054 (.I(W23948), .ZN(O16145));
  INVX1 G40055 (.I(W15372), .ZN(O16157));
  INVX1 G40056 (.I(W72), .ZN(W3820));
  INVX1 G40057 (.I(W1710), .ZN(W3822));
  INVX1 G40058 (.I(W9209), .ZN(O16152));
  INVX1 G40059 (.I(W41382), .ZN(O16149));
  INVX1 G40060 (.I(W24144), .ZN(W47145));
  INVX1 G40061 (.I(W2059), .ZN(W3827));
  INVX1 G40062 (.I(W34360), .ZN(O16147));
  INVX1 G40063 (.I(W2467), .ZN(W3829));
  INVX1 G40064 (.I(W46966), .ZN(O16158));
  INVX1 G40065 (.I(W43224), .ZN(O16144));
  INVX1 G40066 (.I(W35722), .ZN(O16143));
  INVX1 G40067 (.I(W13720), .ZN(O16141));
  INVX1 G40068 (.I(W10842), .ZN(O16140));
  INVX1 G40069 (.I(W982), .ZN(O16139));
  INVX1 G40070 (.I(W42074), .ZN(O16138));
  INVX1 G40071 (.I(W2193), .ZN(W3831));
  INVX1 G40072 (.I(I786), .ZN(W3832));
  INVX1 G40073 (.I(W409), .ZN(W3804));
  INVX1 G40074 (.I(W1045), .ZN(W3787));
  INVX1 G40075 (.I(W3281), .ZN(W3790));
  INVX1 G40076 (.I(W13717), .ZN(O16178));
  INVX1 G40077 (.I(W1927), .ZN(O45));
  INVX1 G40078 (.I(I283), .ZN(W3801));
  INVX1 G40079 (.I(W1331), .ZN(W3802));
  INVX1 G40080 (.I(W7207), .ZN(O16172));
  INVX1 G40081 (.I(I973), .ZN(W3803));
  INVX1 G40082 (.I(W17958), .ZN(W46582));
  INVX1 G40083 (.I(I1344), .ZN(W3805));
  INVX1 G40084 (.I(W8398), .ZN(O16168));
  INVX1 G40085 (.I(I1822), .ZN(W3807));
  INVX1 G40086 (.I(I1612), .ZN(W3808));
  INVX1 G40087 (.I(W12459), .ZN(O16165));
  INVX1 G40088 (.I(W3341), .ZN(W3810));
  INVX1 G40089 (.I(I797), .ZN(W3814));
  INVX1 G40090 (.I(W4346), .ZN(O16159));
  INVX1 G40091 (.I(W40556), .ZN(O15196));
  INVX1 G40092 (.I(I655), .ZN(W4950));
  INVX1 G40093 (.I(W19705), .ZN(O15204));
  INVX1 G40094 (.I(W2553), .ZN(W4951));
  INVX1 G40095 (.I(W8373), .ZN(W46030));
  INVX1 G40096 (.I(W4293), .ZN(W46029));
  INVX1 G40097 (.I(W2637), .ZN(W4952));
  INVX1 G40098 (.I(W171), .ZN(W46025));
  INVX1 G40099 (.I(I1372), .ZN(O15199));
  INVX1 G40100 (.I(W22885), .ZN(O15198));
  INVX1 G40101 (.I(W4626), .ZN(W4948));
  INVX1 G40102 (.I(W17688), .ZN(O15195));
  INVX1 G40103 (.I(W16373), .ZN(O15193));
  INVX1 G40104 (.I(W29322), .ZN(O15189));
  INVX1 G40105 (.I(W3589), .ZN(O69));
  INVX1 G40106 (.I(W12537), .ZN(O15186));
  INVX1 G40107 (.I(I446), .ZN(W4963));
  INVX1 G40108 (.I(W1399), .ZN(W4964));
  INVX1 G40109 (.I(W45286), .ZN(O15183));
  INVX1 G40110 (.I(W41370), .ZN(O15218));
  INVX1 G40111 (.I(W43460), .ZN(O15227));
  INVX1 G40112 (.I(W3472), .ZN(W4921));
  INVX1 G40113 (.I(W33316), .ZN(O15226));
  INVX1 G40114 (.I(W2845), .ZN(W4922));
  INVX1 G40115 (.I(W3378), .ZN(W4923));
  INVX1 G40116 (.I(W2759), .ZN(W4924));
  INVX1 G40117 (.I(W11108), .ZN(O15222));
  INVX1 G40118 (.I(W11144), .ZN(O15221));
  INVX1 G40119 (.I(W2964), .ZN(O15220));
  INVX1 G40120 (.I(W38816), .ZN(O15181));
  INVX1 G40121 (.I(W455), .ZN(W4932));
  INVX1 G40122 (.I(I1592), .ZN(W4935));
  INVX1 G40123 (.I(I1907), .ZN(W4936));
  INVX1 G40124 (.I(W2119), .ZN(W4938));
  INVX1 G40125 (.I(W187), .ZN(W4941));
  INVX1 G40126 (.I(W399), .ZN(W4944));
  INVX1 G40127 (.I(W20199), .ZN(W46036));
  INVX1 G40128 (.I(W40137), .ZN(O15207));
  INVX1 G40129 (.I(W2887), .ZN(W5003));
  INVX1 G40130 (.I(W2273), .ZN(W4996));
  INVX1 G40131 (.I(W207), .ZN(W4997));
  INVX1 G40132 (.I(W941), .ZN(W4999));
  INVX1 G40133 (.I(W6431), .ZN(O15153));
  INVX1 G40134 (.I(W30003), .ZN(O15152));
  INVX1 G40135 (.I(W1188), .ZN(W5000));
  INVX1 G40136 (.I(W1801), .ZN(O15150));
  INVX1 G40137 (.I(W31499), .ZN(O15149));
  INVX1 G40138 (.I(W12127), .ZN(W45964));
  INVX1 G40139 (.I(W37333), .ZN(O15158));
  INVX1 G40140 (.I(W45674), .ZN(O15147));
  INVX1 G40141 (.I(W32275), .ZN(O15146));
  INVX1 G40142 (.I(W1731), .ZN(W5004));
  INVX1 G40143 (.I(I1622), .ZN(W5008));
  INVX1 G40144 (.I(W45251), .ZN(O15142));
  INVX1 G40145 (.I(W40474), .ZN(O15139));
  INVX1 G40146 (.I(W227), .ZN(W45953));
  INVX1 G40147 (.I(I292), .ZN(W5013));
  INVX1 G40148 (.I(W3004), .ZN(W4974));
  INVX1 G40149 (.I(W28629), .ZN(W46005));
  INVX1 G40150 (.I(W12954), .ZN(O15180));
  INVX1 G40151 (.I(I1490), .ZN(W4967));
  INVX1 G40152 (.I(W29904), .ZN(W45999));
  INVX1 G40153 (.I(W30161), .ZN(O15175));
  INVX1 G40154 (.I(W1527), .ZN(W4971));
  INVX1 G40155 (.I(W41106), .ZN(O15172));
  INVX1 G40156 (.I(W312), .ZN(W4973));
  INVX1 G40157 (.I(W33535), .ZN(O15228));
  INVX1 G40158 (.I(W36890), .ZN(O15169));
  INVX1 G40159 (.I(W24715), .ZN(O15166));
  INVX1 G40160 (.I(W4920), .ZN(W4984));
  INVX1 G40161 (.I(W19771), .ZN(O15162));
  INVX1 G40162 (.I(W2536), .ZN(O15161));
  INVX1 G40163 (.I(W4631), .ZN(W4986));
  INVX1 G40164 (.I(I329), .ZN(W4991));
  INVX1 G40165 (.I(W846), .ZN(W4992));
  INVX1 G40166 (.I(W45532), .ZN(O15280));
  INVX1 G40167 (.I(I1331), .ZN(W4860));
  INVX1 G40168 (.I(W2402), .ZN(W4861));
  INVX1 G40169 (.I(W27), .ZN(W46137));
  INVX1 G40170 (.I(W14257), .ZN(O15288));
  INVX1 G40171 (.I(I178), .ZN(W4862));
  INVX1 G40172 (.I(W30509), .ZN(O15285));
  INVX1 G40173 (.I(W11948), .ZN(O15283));
  INVX1 G40174 (.I(W3225), .ZN(W4867));
  INVX1 G40175 (.I(W3422), .ZN(W4868));
  INVX1 G40176 (.I(W3790), .ZN(W4857));
  INVX1 G40177 (.I(W41173), .ZN(O15279));
  INVX1 G40178 (.I(W6184), .ZN(O15277));
  INVX1 G40179 (.I(W19962), .ZN(W46122));
  INVX1 G40180 (.I(W5624), .ZN(W46121));
  INVX1 G40181 (.I(W41883), .ZN(W46119));
  INVX1 G40182 (.I(W21778), .ZN(O15275));
  INVX1 G40183 (.I(W26564), .ZN(O15274));
  INVX1 G40184 (.I(W1561), .ZN(W4878));
  INVX1 G40185 (.I(I988), .ZN(W4844));
  INVX1 G40186 (.I(W17890), .ZN(O15316));
  INVX1 G40187 (.I(W3679), .ZN(W4836));
  INVX1 G40188 (.I(W23743), .ZN(O15314));
  INVX1 G40189 (.I(W2253), .ZN(O15313));
  INVX1 G40190 (.I(W6533), .ZN(O15311));
  INVX1 G40191 (.I(I1425), .ZN(W4839));
  INVX1 G40192 (.I(W37224), .ZN(O15308));
  INVX1 G40193 (.I(W19303), .ZN(O15305));
  INVX1 G40194 (.I(W20531), .ZN(O15304));
  INVX1 G40195 (.I(W1550), .ZN(W4879));
  INVX1 G40196 (.I(W23337), .ZN(O15301));
  INVX1 G40197 (.I(W4820), .ZN(W4847));
  INVX1 G40198 (.I(W1975), .ZN(W4848));
  INVX1 G40199 (.I(W3875), .ZN(W4849));
  INVX1 G40200 (.I(W818), .ZN(W4850));
  INVX1 G40201 (.I(W909), .ZN(W4853));
  INVX1 G40202 (.I(W4341), .ZN(W4854));
  INVX1 G40203 (.I(W2977), .ZN(W4856));
  INVX1 G40204 (.I(W1998), .ZN(W4914));
  INVX1 G40205 (.I(W2300), .ZN(W4905));
  INVX1 G40206 (.I(W32909), .ZN(O15248));
  INVX1 G40207 (.I(W8048), .ZN(O15247));
  INVX1 G40208 (.I(W5352), .ZN(O15246));
  INVX1 G40209 (.I(W356), .ZN(W4906));
  INVX1 G40210 (.I(W1018), .ZN(W4907));
  INVX1 G40211 (.I(W30732), .ZN(O15244));
  INVX1 G40212 (.I(W40307), .ZN(O15243));
  INVX1 G40213 (.I(W4565), .ZN(W4913));
  INVX1 G40214 (.I(W10048), .ZN(O15250));
  INVX1 G40215 (.I(W2051), .ZN(O15239));
  INVX1 G40216 (.I(W4541), .ZN(W4917));
  INVX1 G40217 (.I(W11214), .ZN(O15236));
  INVX1 G40218 (.I(W24425), .ZN(O15234));
  INVX1 G40219 (.I(W19032), .ZN(O15233));
  INVX1 G40220 (.I(I895), .ZN(O15232));
  INVX1 G40221 (.I(W16807), .ZN(O15230));
  INVX1 G40222 (.I(W11430), .ZN(O15229));
  INVX1 G40223 (.I(W3731), .ZN(W4893));
  INVX1 G40224 (.I(I558), .ZN(W4881));
  INVX1 G40225 (.I(W3963), .ZN(W4882));
  INVX1 G40226 (.I(W3163), .ZN(O15268));
  INVX1 G40227 (.I(I656), .ZN(W4887));
  INVX1 G40228 (.I(W7365), .ZN(O15265));
  INVX1 G40229 (.I(W40639), .ZN(O15264));
  INVX1 G40230 (.I(W18740), .ZN(O15263));
  INVX1 G40231 (.I(I1704), .ZN(W4890));
  INVX1 G40232 (.I(W23367), .ZN(O15137));
  INVX1 G40233 (.I(W3983), .ZN(W4894));
  INVX1 G40234 (.I(W21065), .ZN(O15259));
  INVX1 G40235 (.I(W12530), .ZN(O15258));
  INVX1 G40236 (.I(W31461), .ZN(O15257));
  INVX1 G40237 (.I(W4628), .ZN(W4896));
  INVX1 G40238 (.I(I330), .ZN(W4898));
  INVX1 G40239 (.I(W1493), .ZN(W4899));
  INVX1 G40240 (.I(W15373), .ZN(W46091));
  INVX1 G40241 (.I(W3063), .ZN(W5162));
  INVX1 G40242 (.I(W4223), .ZN(W5147));
  INVX1 G40243 (.I(W2981), .ZN(O74));
  INVX1 G40244 (.I(W45083), .ZN(W45811));
  INVX1 G40245 (.I(W3708), .ZN(W5154));
  INVX1 G40246 (.I(W10624), .ZN(W12659));
  INVX1 G40247 (.I(W19744), .ZN(O15025));
  INVX1 G40248 (.I(I694), .ZN(W5158));
  INVX1 G40249 (.I(W44884), .ZN(O15023));
  INVX1 G40250 (.I(W19480), .ZN(O15022));
  INVX1 G40251 (.I(W4654), .ZN(W5143));
  INVX1 G40252 (.I(W43845), .ZN(O15019));
  INVX1 G40253 (.I(W4007), .ZN(W5163));
  INVX1 G40254 (.I(W21489), .ZN(O15017));
  INVX1 G40255 (.I(W18429), .ZN(O15014));
  INVX1 G40256 (.I(W12035), .ZN(O15012));
  INVX1 G40257 (.I(W2276), .ZN(W5169));
  INVX1 G40258 (.I(W1119), .ZN(O77));
  INVX1 G40259 (.I(W1398), .ZN(W5174));
  INVX1 G40260 (.I(W1179), .ZN(W5129));
  INVX1 G40261 (.I(W8903), .ZN(W45845));
  INVX1 G40262 (.I(W13), .ZN(W5120));
  INVX1 G40263 (.I(W9579), .ZN(O15052));
  INVX1 G40264 (.I(W33105), .ZN(O15051));
  INVX1 G40265 (.I(W17830), .ZN(W45841));
  INVX1 G40266 (.I(W26493), .ZN(O15049));
  INVX1 G40267 (.I(W22354), .ZN(O15048));
  INVX1 G40268 (.I(W30403), .ZN(O15045));
  INVX1 G40269 (.I(W21321), .ZN(O15044));
  INVX1 G40270 (.I(W2134), .ZN(W5175));
  INVX1 G40271 (.I(W13540), .ZN(O15042));
  INVX1 G40272 (.I(W15891), .ZN(O15038));
  INVX1 G40273 (.I(W4627), .ZN(W5135));
  INVX1 G40274 (.I(I1314), .ZN(W5138));
  INVX1 G40275 (.I(W4634), .ZN(W5139));
  INVX1 G40276 (.I(I1942), .ZN(O15034));
  INVX1 G40277 (.I(W37504), .ZN(O15033));
  INVX1 G40278 (.I(I72), .ZN(W5141));
  INVX1 G40279 (.I(W1004), .ZN(O14975));
  INVX1 G40280 (.I(W35174), .ZN(O14985));
  INVX1 G40281 (.I(W3198), .ZN(W5195));
  INVX1 G40282 (.I(W20160), .ZN(W45758));
  INVX1 G40283 (.I(W1848), .ZN(W5198));
  INVX1 G40284 (.I(W12764), .ZN(O14979));
  INVX1 G40285 (.I(W2244), .ZN(W5202));
  INVX1 G40286 (.I(W1157), .ZN(W45751));
  INVX1 G40287 (.I(W24060), .ZN(O14977));
  INVX1 G40288 (.I(W13672), .ZN(O14976));
  INVX1 G40289 (.I(W5117), .ZN(W5194));
  INVX1 G40290 (.I(W354), .ZN(W5204));
  INVX1 G40291 (.I(W3885), .ZN(W5206));
  INVX1 G40292 (.I(I902), .ZN(W5207));
  INVX1 G40293 (.I(W10609), .ZN(O14968));
  INVX1 G40294 (.I(W26026), .ZN(O14967));
  INVX1 G40295 (.I(W41576), .ZN(O14966));
  INVX1 G40296 (.I(W3271), .ZN(W5210));
  INVX1 G40297 (.I(W19779), .ZN(O14963));
  INVX1 G40298 (.I(W38174), .ZN(O14995));
  INVX1 G40299 (.I(I117), .ZN(O15006));
  INVX1 G40300 (.I(W909), .ZN(W5178));
  INVX1 G40301 (.I(W40016), .ZN(O15002));
  INVX1 G40302 (.I(W3859), .ZN(W5179));
  INVX1 G40303 (.I(W21764), .ZN(O15000));
  INVX1 G40304 (.I(W2437), .ZN(O14999));
  INVX1 G40305 (.I(I1492), .ZN(W45776));
  INVX1 G40306 (.I(W7197), .ZN(O14996));
  INVX1 G40307 (.I(W23319), .ZN(O15054));
  INVX1 G40308 (.I(W3643), .ZN(W5185));
  INVX1 G40309 (.I(W27989), .ZN(W45771));
  INVX1 G40310 (.I(W2177), .ZN(W5186));
  INVX1 G40311 (.I(W12806), .ZN(O14992));
  INVX1 G40312 (.I(W3401), .ZN(W5189));
  INVX1 G40313 (.I(W22995), .ZN(W45766));
  INVX1 G40314 (.I(W135), .ZN(W5191));
  INVX1 G40315 (.I(W23246), .ZN(O14987));
  INVX1 G40316 (.I(W4839), .ZN(W5049));
  INVX1 G40317 (.I(W38002), .ZN(O15114));
  INVX1 G40318 (.I(W553), .ZN(W5035));
  INVX1 G40319 (.I(W17162), .ZN(W45918));
  INVX1 G40320 (.I(W31), .ZN(W5036));
  INVX1 G40321 (.I(W10239), .ZN(O15111));
  INVX1 G40322 (.I(W4085), .ZN(W5044));
  INVX1 G40323 (.I(W2529), .ZN(W5045));
  INVX1 G40324 (.I(W3737), .ZN(W5046));
  INVX1 G40325 (.I(W10989), .ZN(O15105));
  INVX1 G40326 (.I(W19078), .ZN(W45922));
  INVX1 G40327 (.I(I1189), .ZN(W5053));
  INVX1 G40328 (.I(W3241), .ZN(W5055));
  INVX1 G40329 (.I(W896), .ZN(W5056));
  INVX1 G40330 (.I(W1783), .ZN(W5058));
  INVX1 G40331 (.I(W764), .ZN(O15099));
  INVX1 G40332 (.I(W1569), .ZN(W5064));
  INVX1 G40333 (.I(W757), .ZN(W5065));
  INVX1 G40334 (.I(W20642), .ZN(O15095));
  INVX1 G40335 (.I(W12494), .ZN(O15122));
  INVX1 G40336 (.I(W8926), .ZN(O15136));
  INVX1 G40337 (.I(W2336), .ZN(W5017));
  INVX1 G40338 (.I(W16506), .ZN(O15133));
  INVX1 G40339 (.I(W26317), .ZN(O15131));
  INVX1 G40340 (.I(I995), .ZN(O15130));
  INVX1 G40341 (.I(W40616), .ZN(O15129));
  INVX1 G40342 (.I(I762), .ZN(W5020));
  INVX1 G40343 (.I(W4556), .ZN(W5023));
  INVX1 G40344 (.I(W321), .ZN(W5025));
  INVX1 G40345 (.I(W29263), .ZN(O15094));
  INVX1 G40346 (.I(W22985), .ZN(O15120));
  INVX1 G40347 (.I(W285), .ZN(W5029));
  INVX1 G40348 (.I(W27728), .ZN(O15117));
  INVX1 G40349 (.I(W1369), .ZN(W5032));
  INVX1 G40350 (.I(W2385), .ZN(W5033));
  INVX1 G40351 (.I(W10625), .ZN(W45925));
  INVX1 G40352 (.I(W3649), .ZN(W45924));
  INVX1 G40353 (.I(W17287), .ZN(W45923));
  INVX1 G40354 (.I(W4010), .ZN(W5103));
  INVX1 G40355 (.I(W27804), .ZN(O15072));
  INVX1 G40356 (.I(W25909), .ZN(O15071));
  INVX1 G40357 (.I(W30201), .ZN(W45867));
  INVX1 G40358 (.I(W21129), .ZN(O15070));
  INVX1 G40359 (.I(W27656), .ZN(O15069));
  INVX1 G40360 (.I(W42831), .ZN(O15067));
  INVX1 G40361 (.I(W1237), .ZN(W5093));
  INVX1 G40362 (.I(W21), .ZN(W5094));
  INVX1 G40363 (.I(I1278), .ZN(W5098));
  INVX1 G40364 (.I(W39611), .ZN(O15073));
  INVX1 G40365 (.I(W153), .ZN(W5104));
  INVX1 G40366 (.I(W36886), .ZN(O15061));
  INVX1 G40367 (.I(W4639), .ZN(W5107));
  INVX1 G40368 (.I(I1825), .ZN(W5109));
  INVX1 G40369 (.I(I421), .ZN(W5110));
  INVX1 G40370 (.I(W2700), .ZN(W5117));
  INVX1 G40371 (.I(W4906), .ZN(W5118));
  INVX1 G40372 (.I(I61), .ZN(W5119));
  INVX1 G40373 (.I(W35710), .ZN(O15084));
  INVX1 G40374 (.I(W31563), .ZN(W45895));
  INVX1 G40375 (.I(I245), .ZN(W5070));
  INVX1 G40376 (.I(W2042), .ZN(W5075));
  INVX1 G40377 (.I(W3447), .ZN(O15088));
  INVX1 G40378 (.I(W12544), .ZN(O15087));
  INVX1 G40379 (.I(W35693), .ZN(O15085));
  INVX1 G40380 (.I(W29061), .ZN(W45884));
  INVX1 G40381 (.I(W16124), .ZN(W45883));
  INVX1 G40382 (.I(W3369), .ZN(O15317));
  INVX1 G40383 (.I(I1414), .ZN(W5078));
  INVX1 G40384 (.I(I776), .ZN(W5079));
  INVX1 G40385 (.I(W3488), .ZN(W5080));
  INVX1 G40386 (.I(I610), .ZN(W5082));
  INVX1 G40387 (.I(W1898), .ZN(W5083));
  INVX1 G40388 (.I(W25073), .ZN(O15078));
  INVX1 G40389 (.I(I587), .ZN(W5088));
  INVX1 G40390 (.I(I1256), .ZN(O15074));
  INVX1 G40391 (.I(I454), .ZN(W4597));
  INVX1 G40392 (.I(W2820), .ZN(W4586));
  INVX1 G40393 (.I(W59), .ZN(W4587));
  INVX1 G40394 (.I(W2986), .ZN(W4589));
  INVX1 G40395 (.I(W4148), .ZN(W4591));
  INVX1 G40396 (.I(W6027), .ZN(O15544));
  INVX1 G40397 (.I(I1626), .ZN(W4594));
  INVX1 G40398 (.I(I1717), .ZN(W4595));
  INVX1 G40399 (.I(I266), .ZN(O61));
  INVX1 G40400 (.I(W16194), .ZN(O15540));
  INVX1 G40401 (.I(I1759), .ZN(O15551));
  INVX1 G40402 (.I(W40089), .ZN(O15537));
  INVX1 G40403 (.I(W4383), .ZN(W4600));
  INVX1 G40404 (.I(I1224), .ZN(W4611));
  INVX1 G40405 (.I(W289), .ZN(W4613));
  INVX1 G40406 (.I(W10411), .ZN(O15532));
  INVX1 G40407 (.I(I1756), .ZN(W4614));
  INVX1 G40408 (.I(W366), .ZN(O15530));
  INVX1 G40409 (.I(W605), .ZN(W4615));
  INVX1 G40410 (.I(W1426), .ZN(W4570));
  INVX1 G40411 (.I(W2239), .ZN(W4559));
  INVX1 G40412 (.I(I79), .ZN(O15572));
  INVX1 G40413 (.I(W1070), .ZN(W4560));
  INVX1 G40414 (.I(W2620), .ZN(W4561));
  INVX1 G40415 (.I(I1212), .ZN(W4566));
  INVX1 G40416 (.I(W25413), .ZN(W46459));
  INVX1 G40417 (.I(W25344), .ZN(O15566));
  INVX1 G40418 (.I(I1578), .ZN(W4568));
  INVX1 G40419 (.I(W7429), .ZN(O15563));
  INVX1 G40420 (.I(I643), .ZN(W4617));
  INVX1 G40421 (.I(W1706), .ZN(W4571));
  INVX1 G40422 (.I(W38424), .ZN(O15560));
  INVX1 G40423 (.I(W2530), .ZN(W4572));
  INVX1 G40424 (.I(W403), .ZN(W4573));
  INVX1 G40425 (.I(W41851), .ZN(O15557));
  INVX1 G40426 (.I(W1392), .ZN(W4578));
  INVX1 G40427 (.I(W3576), .ZN(W4581));
  INVX1 G40428 (.I(W36861), .ZN(W46443));
  INVX1 G40429 (.I(W4476), .ZN(W4655));
  INVX1 G40430 (.I(W6887), .ZN(O15506));
  INVX1 G40431 (.I(W213), .ZN(W4647));
  INVX1 G40432 (.I(W4615), .ZN(W4648));
  INVX1 G40433 (.I(W4561), .ZN(W4650));
  INVX1 G40434 (.I(W4286), .ZN(W4651));
  INVX1 G40435 (.I(W100), .ZN(W4653));
  INVX1 G40436 (.I(W205), .ZN(W4654));
  INVX1 G40437 (.I(I1075), .ZN(O15498));
  INVX1 G40438 (.I(W7673), .ZN(O15497));
  INVX1 G40439 (.I(W1486), .ZN(W4643));
  INVX1 G40440 (.I(W24944), .ZN(O15494));
  INVX1 G40441 (.I(W1405), .ZN(W4657));
  INVX1 G40442 (.I(W13016), .ZN(W46377));
  INVX1 G40443 (.I(W20435), .ZN(O15493));
  INVX1 G40444 (.I(W3065), .ZN(W4658));
  INVX1 G40445 (.I(W2520), .ZN(W4660));
  INVX1 G40446 (.I(W158), .ZN(W4662));
  INVX1 G40447 (.I(I1854), .ZN(W4664));
  INVX1 G40448 (.I(W41978), .ZN(O15518));
  INVX1 G40449 (.I(W1769), .ZN(W4619));
  INVX1 G40450 (.I(I166), .ZN(O15527));
  INVX1 G40451 (.I(W2654), .ZN(W4623));
  INVX1 G40452 (.I(W19231), .ZN(W46411));
  INVX1 G40453 (.I(W9695), .ZN(O15524));
  INVX1 G40454 (.I(W656), .ZN(W4625));
  INVX1 G40455 (.I(I102), .ZN(W4629));
  INVX1 G40456 (.I(W551), .ZN(W4631));
  INVX1 G40457 (.I(W1834), .ZN(W4557));
  INVX1 G40458 (.I(W2718), .ZN(W46402));
  INVX1 G40459 (.I(W41002), .ZN(O15516));
  INVX1 G40460 (.I(W2444), .ZN(W4636));
  INVX1 G40461 (.I(I392), .ZN(W4638));
  INVX1 G40462 (.I(W45836), .ZN(O15512));
  INVX1 G40463 (.I(W2214), .ZN(W4639));
  INVX1 G40464 (.I(W39171), .ZN(O15510));
  INVX1 G40465 (.I(W1717), .ZN(W4641));
  INVX1 G40466 (.I(W341), .ZN(W4486));
  INVX1 G40467 (.I(I1870), .ZN(W4457));
  INVX1 G40468 (.I(I712), .ZN(W4463));
  INVX1 G40469 (.I(W4187), .ZN(W4474));
  INVX1 G40470 (.I(W26523), .ZN(W46546));
  INVX1 G40471 (.I(I562), .ZN(W4476));
  INVX1 G40472 (.I(I1770), .ZN(W4477));
  INVX1 G40473 (.I(W1327), .ZN(W4480));
  INVX1 G40474 (.I(W16439), .ZN(O15636));
  INVX1 G40475 (.I(W24650), .ZN(O15635));
  INVX1 G40476 (.I(W17264), .ZN(O15648));
  INVX1 G40477 (.I(I686), .ZN(O15631));
  INVX1 G40478 (.I(I1149), .ZN(W4488));
  INVX1 G40479 (.I(W40695), .ZN(O15628));
  INVX1 G40480 (.I(W3154), .ZN(W4490));
  INVX1 G40481 (.I(W11983), .ZN(O15626));
  INVX1 G40482 (.I(W19663), .ZN(O15624));
  INVX1 G40483 (.I(W26595), .ZN(O15622));
  INVX1 G40484 (.I(W28091), .ZN(O15621));
  INVX1 G40485 (.I(I1914), .ZN(W4445));
  INVX1 G40486 (.I(W1112), .ZN(W4427));
  INVX1 G40487 (.I(W4040), .ZN(W4429));
  INVX1 G40488 (.I(I102), .ZN(W4430));
  INVX1 G40489 (.I(W3891), .ZN(W4431));
  INVX1 G40490 (.I(W19684), .ZN(O15666));
  INVX1 G40491 (.I(W2292), .ZN(O15665));
  INVX1 G40492 (.I(I362), .ZN(W4434));
  INVX1 G40493 (.I(W3639), .ZN(W4438));
  INVX1 G40494 (.I(W3403), .ZN(W4440));
  INVX1 G40495 (.I(W7277), .ZN(O15619));
  INVX1 G40496 (.I(W1182), .ZN(W4446));
  INVX1 G40497 (.I(W43369), .ZN(O15656));
  INVX1 G40498 (.I(W13610), .ZN(O15655));
  INVX1 G40499 (.I(W13441), .ZN(O15654));
  INVX1 G40500 (.I(W1811), .ZN(W4447));
  INVX1 G40501 (.I(W32483), .ZN(W46560));
  INVX1 G40502 (.I(W1128), .ZN(O15651));
  INVX1 G40503 (.I(W2611), .ZN(W4455));
  INVX1 G40504 (.I(W30165), .ZN(O15585));
  INVX1 G40505 (.I(W2751), .ZN(W4531));
  INVX1 G40506 (.I(W1429), .ZN(W4534));
  INVX1 G40507 (.I(I576), .ZN(W4536));
  INVX1 G40508 (.I(W3653), .ZN(W46489));
  INVX1 G40509 (.I(W5322), .ZN(O15590));
  INVX1 G40510 (.I(W20020), .ZN(O15589));
  INVX1 G40511 (.I(W17539), .ZN(O15588));
  INVX1 G40512 (.I(W43976), .ZN(O15587));
  INVX1 G40513 (.I(W3112), .ZN(W4540));
  INVX1 G40514 (.I(W2384), .ZN(O59));
  INVX1 G40515 (.I(W30405), .ZN(W46480));
  INVX1 G40516 (.I(W43793), .ZN(O15582));
  INVX1 G40517 (.I(I1934), .ZN(W4546));
  INVX1 G40518 (.I(W38389), .ZN(O15580));
  INVX1 G40519 (.I(W1048), .ZN(W4549));
  INVX1 G40520 (.I(W8135), .ZN(O15579));
  INVX1 G40521 (.I(W306), .ZN(W4550));
  INVX1 G40522 (.I(I445), .ZN(W4553));
  INVX1 G40523 (.I(W46078), .ZN(W46509));
  INVX1 G40524 (.I(W518), .ZN(W4498));
  INVX1 G40525 (.I(W41434), .ZN(O15617));
  INVX1 G40526 (.I(W3446), .ZN(W4499));
  INVX1 G40527 (.I(W5274), .ZN(W46518));
  INVX1 G40528 (.I(I1164), .ZN(W4507));
  INVX1 G40529 (.I(W1954), .ZN(W4508));
  INVX1 G40530 (.I(W38751), .ZN(W46512));
  INVX1 G40531 (.I(I32), .ZN(W4510));
  INVX1 G40532 (.I(W2748), .ZN(O15488));
  INVX1 G40533 (.I(W33367), .ZN(O15609));
  INVX1 G40534 (.I(W2139), .ZN(W4518));
  INVX1 G40535 (.I(W2030), .ZN(W4519));
  INVX1 G40536 (.I(W2014), .ZN(W4521));
  INVX1 G40537 (.I(W3977), .ZN(W4523));
  INVX1 G40538 (.I(W4165), .ZN(W4524));
  INVX1 G40539 (.I(W4084), .ZN(W4526));
  INVX1 G40540 (.I(W2739), .ZN(W4528));
  INVX1 G40541 (.I(W4424), .ZN(W4790));
  INVX1 G40542 (.I(W282), .ZN(W4782));
  INVX1 G40543 (.I(I485), .ZN(W4783));
  INVX1 G40544 (.I(I1343), .ZN(W4785));
  INVX1 G40545 (.I(W27324), .ZN(O15372));
  INVX1 G40546 (.I(W41365), .ZN(O15371));
  INVX1 G40547 (.I(W9092), .ZN(O15370));
  INVX1 G40548 (.I(W26527), .ZN(W46233));
  INVX1 G40549 (.I(W2110), .ZN(W4787));
  INVX1 G40550 (.I(W569), .ZN(W4789));
  INVX1 G40551 (.I(I888), .ZN(W4780));
  INVX1 G40552 (.I(W614), .ZN(W4796));
  INVX1 G40553 (.I(W10581), .ZN(O15363));
  INVX1 G40554 (.I(W20226), .ZN(O15362));
  INVX1 G40555 (.I(W42518), .ZN(O15361));
  INVX1 G40556 (.I(W27049), .ZN(O15360));
  INVX1 G40557 (.I(W3424), .ZN(W4800));
  INVX1 G40558 (.I(W992), .ZN(W4801));
  INVX1 G40559 (.I(W11047), .ZN(W46215));
  INVX1 G40560 (.I(W25695), .ZN(O15386));
  INVX1 G40561 (.I(W8414), .ZN(O15402));
  INVX1 G40562 (.I(W2634), .ZN(W4755));
  INVX1 G40563 (.I(W1273), .ZN(W4758));
  INVX1 G40564 (.I(W22180), .ZN(O15396));
  INVX1 G40565 (.I(W41261), .ZN(O15395));
  INVX1 G40566 (.I(W219), .ZN(W4760));
  INVX1 G40567 (.I(W3364), .ZN(W4761));
  INVX1 G40568 (.I(W3268), .ZN(W4764));
  INVX1 G40569 (.I(W44529), .ZN(O15390));
  INVX1 G40570 (.I(W29656), .ZN(O15356));
  INVX1 G40571 (.I(W19008), .ZN(O15385));
  INVX1 G40572 (.I(I786), .ZN(W4769));
  INVX1 G40573 (.I(I188), .ZN(W4772));
  INVX1 G40574 (.I(W4672), .ZN(W4774));
  INVX1 G40575 (.I(W3357), .ZN(W4775));
  INVX1 G40576 (.I(W291), .ZN(W4776));
  INVX1 G40577 (.I(W10429), .ZN(O15378));
  INVX1 G40578 (.I(W16934), .ZN(O15376));
  INVX1 G40579 (.I(W34493), .ZN(W46176));
  INVX1 G40580 (.I(I737), .ZN(W4822));
  INVX1 G40581 (.I(W3069), .ZN(W4823));
  INVX1 G40582 (.I(W6890), .ZN(O15333));
  INVX1 G40583 (.I(W3147), .ZN(W4826));
  INVX1 G40584 (.I(W21141), .ZN(O15331));
  INVX1 G40585 (.I(W15140), .ZN(O15329));
  INVX1 G40586 (.I(W40927), .ZN(O15328));
  INVX1 G40587 (.I(W25527), .ZN(O15327));
  INVX1 G40588 (.I(W9937), .ZN(O15326));
  INVX1 G40589 (.I(W23833), .ZN(O15337));
  INVX1 G40590 (.I(W30843), .ZN(O15324));
  INVX1 G40591 (.I(W467), .ZN(O15323));
  INVX1 G40592 (.I(W1780), .ZN(W4829));
  INVX1 G40593 (.I(W34534), .ZN(O15321));
  INVX1 G40594 (.I(W3854), .ZN(W4830));
  INVX1 G40595 (.I(W31636), .ZN(O15319));
  INVX1 G40596 (.I(I1523), .ZN(W4831));
  INVX1 G40597 (.I(W28156), .ZN(W46168));
  INVX1 G40598 (.I(W8746), .ZN(O15347));
  INVX1 G40599 (.I(W3673), .ZN(W4803));
  INVX1 G40600 (.I(W37479), .ZN(O15355));
  INVX1 G40601 (.I(W3019), .ZN(W4805));
  INVX1 G40602 (.I(W38281), .ZN(O15354));
  INVX1 G40603 (.I(W41805), .ZN(O15353));
  INVX1 G40604 (.I(W1667), .ZN(W4808));
  INVX1 G40605 (.I(W4706), .ZN(W4812));
  INVX1 G40606 (.I(W27305), .ZN(W46203));
  INVX1 G40607 (.I(W3061), .ZN(W4753));
  INVX1 G40608 (.I(I1842), .ZN(W4815));
  INVX1 G40609 (.I(W13614), .ZN(O15345));
  INVX1 G40610 (.I(W6102), .ZN(W46197));
  INVX1 G40611 (.I(I1339), .ZN(W4817));
  INVX1 G40612 (.I(W43251), .ZN(W46193));
  INVX1 G40613 (.I(W29195), .ZN(O15340));
  INVX1 G40614 (.I(I1526), .ZN(W4821));
  INVX1 G40615 (.I(W11198), .ZN(O15338));
  INVX1 G40616 (.I(W10742), .ZN(O15455));
  INVX1 G40617 (.I(W10589), .ZN(O15466));
  INVX1 G40618 (.I(I1301), .ZN(W4694));
  INVX1 G40619 (.I(W43643), .ZN(O15462));
  INVX1 G40620 (.I(W4246), .ZN(W4701));
  INVX1 G40621 (.I(I1266), .ZN(W4702));
  INVX1 G40622 (.I(W354), .ZN(W4704));
  INVX1 G40623 (.I(W34992), .ZN(O15458));
  INVX1 G40624 (.I(W1333), .ZN(W4708));
  INVX1 G40625 (.I(W1868), .ZN(W4709));
  INVX1 G40626 (.I(W40845), .ZN(O15467));
  INVX1 G40627 (.I(W28113), .ZN(O15454));
  INVX1 G40628 (.I(W82), .ZN(W4710));
  INVX1 G40629 (.I(W3730), .ZN(W4711));
  INVX1 G40630 (.I(W45884), .ZN(O15451));
  INVX1 G40631 (.I(I24), .ZN(W4714));
  INVX1 G40632 (.I(W1637), .ZN(O15449));
  INVX1 G40633 (.I(W366), .ZN(W4715));
  INVX1 G40634 (.I(W21945), .ZN(O15447));
  INVX1 G40635 (.I(W21035), .ZN(W46355));
  INVX1 G40636 (.I(I1457), .ZN(W4666));
  INVX1 G40637 (.I(W27020), .ZN(O15486));
  INVX1 G40638 (.I(W2400), .ZN(O15485));
  INVX1 G40639 (.I(W1261), .ZN(W4677));
  INVX1 G40640 (.I(W13874), .ZN(O15481));
  INVX1 G40641 (.I(W117), .ZN(W4679));
  INVX1 G40642 (.I(W395), .ZN(W4681));
  INVX1 G40643 (.I(W4054), .ZN(W46357));
  INVX1 G40644 (.I(W12710), .ZN(O15478));
  INVX1 G40645 (.I(W6190), .ZN(O15446));
  INVX1 G40646 (.I(W21536), .ZN(W46353));
  INVX1 G40647 (.I(W45704), .ZN(O15476));
  INVX1 G40648 (.I(W1935), .ZN(W4684));
  INVX1 G40649 (.I(W3948), .ZN(W4689));
  INVX1 G40650 (.I(W252), .ZN(W4690));
  INVX1 G40651 (.I(W38555), .ZN(O15470));
  INVX1 G40652 (.I(I683), .ZN(W4692));
  INVX1 G40653 (.I(W1379), .ZN(W4693));
  INVX1 G40654 (.I(W4330), .ZN(W4745));
  INVX1 G40655 (.I(W28267), .ZN(O15422));
  INVX1 G40656 (.I(W1888), .ZN(W4734));
  INVX1 G40657 (.I(W3668), .ZN(W4735));
  INVX1 G40658 (.I(W3189), .ZN(W4737));
  INVX1 G40659 (.I(I380), .ZN(W4739));
  INVX1 G40660 (.I(W45445), .ZN(O15416));
  INVX1 G40661 (.I(W5805), .ZN(O15414));
  INVX1 G40662 (.I(W32462), .ZN(W46282));
  INVX1 G40663 (.I(W3922), .ZN(W4743));
  INVX1 G40664 (.I(W3111), .ZN(W4733));
  INVX1 G40665 (.I(W16922), .ZN(O15411));
  INVX1 G40666 (.I(W792), .ZN(W4748));
  INVX1 G40667 (.I(W20595), .ZN(W46277));
  INVX1 G40668 (.I(W4431), .ZN(W4749));
  INVX1 G40669 (.I(W36021), .ZN(O15408));
  INVX1 G40670 (.I(W45278), .ZN(O15406));
  INVX1 G40671 (.I(W904), .ZN(W4751));
  INVX1 G40672 (.I(W5272), .ZN(O15404));
  INVX1 G40673 (.I(W22940), .ZN(O15432));
  INVX1 G40674 (.I(W15736), .ZN(W46317));
  INVX1 G40675 (.I(W21069), .ZN(O15445));
  INVX1 G40676 (.I(W34932), .ZN(O15444));
  INVX1 G40677 (.I(W4750), .ZN(W46313));
  INVX1 G40678 (.I(W14660), .ZN(O15442));
  INVX1 G40679 (.I(W16269), .ZN(O15435));
  INVX1 G40680 (.I(W31452), .ZN(O15434));
  INVX1 G40681 (.I(W4060), .ZN(W4726));
  INVX1 G40682 (.I(W1234), .ZN(W43917));
  INVX1 G40683 (.I(W2615), .ZN(W4727));
  INVX1 G40684 (.I(W1010), .ZN(O15430));
  INVX1 G40685 (.I(I1118), .ZN(W4729));
  INVX1 G40686 (.I(W43766), .ZN(O15429));
  INVX1 G40687 (.I(W39764), .ZN(O15428));
  INVX1 G40688 (.I(W27478), .ZN(O15427));
  INVX1 G40689 (.I(W24668), .ZN(O15426));
  INVX1 G40690 (.I(W4692), .ZN(W4730));
  INVX1 G40691 (.I(W8299), .ZN(O1987));
  INVX1 G40692 (.I(W1388), .ZN(O5335));
  INVX1 G40693 (.I(W19596), .ZN(W20337));
  INVX1 G40694 (.I(W5102), .ZN(W20338));
  INVX1 G40695 (.I(I348), .ZN(O5334));
  INVX1 G40696 (.I(W2920), .ZN(W20339));
  INVX1 G40697 (.I(W18639), .ZN(O5333));
  INVX1 G40698 (.I(W7668), .ZN(W20345));
  INVX1 G40699 (.I(W4999), .ZN(O1982));
  INVX1 G40700 (.I(W16899), .ZN(O1983));
  INVX1 G40701 (.I(W13545), .ZN(O1986));
  INVX1 G40702 (.I(W5666), .ZN(W20334));
  INVX1 G40703 (.I(W10843), .ZN(O1989));
  INVX1 G40704 (.I(I36), .ZN(W30428));
  INVX1 G40705 (.I(W3066), .ZN(W20362));
  INVX1 G40706 (.I(W657), .ZN(W30424));
  INVX1 G40707 (.I(W6071), .ZN(W20366));
  INVX1 G40708 (.I(W10742), .ZN(W20367));
  INVX1 G40709 (.I(W8858), .ZN(O1991));
  INVX1 G40710 (.I(W3764), .ZN(W20370));
  INVX1 G40711 (.I(W10183), .ZN(O1992));
  INVX1 G40712 (.I(W14194), .ZN(W20318));
  INVX1 G40713 (.I(W29170), .ZN(O5354));
  INVX1 G40714 (.I(W11621), .ZN(W20310));
  INVX1 G40715 (.I(W28837), .ZN(W30472));
  INVX1 G40716 (.I(W6868), .ZN(O1973));
  INVX1 G40717 (.I(W12051), .ZN(W20312));
  INVX1 G40718 (.I(W13027), .ZN(W30468));
  INVX1 G40719 (.I(W9466), .ZN(O1974));
  INVX1 G40720 (.I(W12160), .ZN(W20315));
  INVX1 G40721 (.I(W11723), .ZN(W30465));
  INVX1 G40722 (.I(W1354), .ZN(O1993));
  INVX1 G40723 (.I(W29355), .ZN(W30461));
  INVX1 G40724 (.I(W12803), .ZN(O5346));
  INVX1 G40725 (.I(W15281), .ZN(W20323));
  INVX1 G40726 (.I(W9395), .ZN(W20327));
  INVX1 G40727 (.I(W9533), .ZN(W30454));
  INVX1 G40728 (.I(I85), .ZN(O5341));
  INVX1 G40729 (.I(W23603), .ZN(O5339));
  INVX1 G40730 (.I(W12928), .ZN(O5338));
  INVX1 G40731 (.I(W4164), .ZN(O1976));
  INVX1 G40732 (.I(W16431), .ZN(O5304));
  INVX1 G40733 (.I(W14653), .ZN(O5311));
  INVX1 G40734 (.I(W1946), .ZN(O2000));
  INVX1 G40735 (.I(W20167), .ZN(W20402));
  INVX1 G40736 (.I(W25074), .ZN(O5309));
  INVX1 G40737 (.I(W2809), .ZN(W20405));
  INVX1 G40738 (.I(W6465), .ZN(W20406));
  INVX1 G40739 (.I(W1293), .ZN(W30381));
  INVX1 G40740 (.I(W8804), .ZN(W30380));
  INVX1 G40741 (.I(W15501), .ZN(W20413));
  INVX1 G40742 (.I(W29785), .ZN(W30391));
  INVX1 G40743 (.I(W18217), .ZN(O2005));
  INVX1 G40744 (.I(W21154), .ZN(W30375));
  INVX1 G40745 (.I(W6716), .ZN(W30374));
  INVX1 G40746 (.I(W3056), .ZN(W30372));
  INVX1 G40747 (.I(W5819), .ZN(O2006));
  INVX1 G40748 (.I(W4458), .ZN(O5302));
  INVX1 G40749 (.I(W10863), .ZN(W20419));
  INVX1 G40750 (.I(I408), .ZN(O5300));
  INVX1 G40751 (.I(W14229), .ZN(W20420));
  INVX1 G40752 (.I(W4555), .ZN(W20385));
  INVX1 G40753 (.I(W20513), .ZN(O5324));
  INVX1 G40754 (.I(W7763), .ZN(O5323));
  INVX1 G40755 (.I(W9374), .ZN(W30414));
  INVX1 G40756 (.I(W14278), .ZN(W30413));
  INVX1 G40757 (.I(W6219), .ZN(W20378));
  INVX1 G40758 (.I(W2146), .ZN(W20380));
  INVX1 G40759 (.I(W28718), .ZN(O5321));
  INVX1 G40760 (.I(W21635), .ZN(O5320));
  INVX1 G40761 (.I(W20293), .ZN(W20384));
  INVX1 G40762 (.I(W9031), .ZN(W20309));
  INVX1 G40763 (.I(I1820), .ZN(W30405));
  INVX1 G40764 (.I(W17867), .ZN(O5319));
  INVX1 G40765 (.I(W13302), .ZN(W30403));
  INVX1 G40766 (.I(W10117), .ZN(W30402));
  INVX1 G40767 (.I(W4081), .ZN(W20387));
  INVX1 G40768 (.I(W4395), .ZN(O5315));
  INVX1 G40769 (.I(W16679), .ZN(W20391));
  INVX1 G40770 (.I(W15459), .ZN(W20393));
  INVX1 G40771 (.I(W18693), .ZN(W20399));
  INVX1 G40772 (.I(W16488), .ZN(W20252));
  INVX1 G40773 (.I(W16351), .ZN(W20235));
  INVX1 G40774 (.I(W928), .ZN(W30561));
  INVX1 G40775 (.I(W15231), .ZN(W20236));
  INVX1 G40776 (.I(I907), .ZN(W30557));
  INVX1 G40777 (.I(W18570), .ZN(W30554));
  INVX1 G40778 (.I(W10262), .ZN(W20244));
  INVX1 G40779 (.I(W16570), .ZN(W20248));
  INVX1 G40780 (.I(W17104), .ZN(W20251));
  INVX1 G40781 (.I(W12034), .ZN(W30548));
  INVX1 G40782 (.I(W19549), .ZN(W30547));
  INVX1 G40783 (.I(W18509), .ZN(O5396));
  INVX1 G40784 (.I(W889), .ZN(W20254));
  INVX1 G40785 (.I(W17965), .ZN(W30543));
  INVX1 G40786 (.I(W14719), .ZN(O1964));
  INVX1 G40787 (.I(W20676), .ZN(O5386));
  INVX1 G40788 (.I(W2437), .ZN(W20256));
  INVX1 G40789 (.I(W8706), .ZN(O5385));
  INVX1 G40790 (.I(W18798), .ZN(W30538));
  INVX1 G40791 (.I(W7288), .ZN(W20259));
  INVX1 G40792 (.I(W7940), .ZN(O5383));
  INVX1 G40793 (.I(W3031), .ZN(W20224));
  INVX1 G40794 (.I(W26976), .ZN(O5406));
  INVX1 G40795 (.I(W13917), .ZN(W30588));
  INVX1 G40796 (.I(W19611), .ZN(W30587));
  INVX1 G40797 (.I(W3239), .ZN(O5404));
  INVX1 G40798 (.I(W11009), .ZN(W20211));
  INVX1 G40799 (.I(W5719), .ZN(W20215));
  INVX1 G40800 (.I(I872), .ZN(W20219));
  INVX1 G40801 (.I(W6934), .ZN(W20221));
  INVX1 G40802 (.I(W2313), .ZN(W20223));
  INVX1 G40803 (.I(W10078), .ZN(W20264));
  INVX1 G40804 (.I(W27923), .ZN(W30574));
  INVX1 G40805 (.I(W13096), .ZN(W20225));
  INVX1 G40806 (.I(W2268), .ZN(W30572));
  INVX1 G40807 (.I(W13206), .ZN(O5399));
  INVX1 G40808 (.I(W22633), .ZN(W30570));
  INVX1 G40809 (.I(W1120), .ZN(W20228));
  INVX1 G40810 (.I(W9831), .ZN(W20230));
  INVX1 G40811 (.I(I613), .ZN(W30567));
  INVX1 G40812 (.I(W9521), .ZN(W30566));
  INVX1 G40813 (.I(W15174), .ZN(W20296));
  INVX1 G40814 (.I(W5109), .ZN(W20282));
  INVX1 G40815 (.I(W2214), .ZN(O1968));
  INVX1 G40816 (.I(W14512), .ZN(O5366));
  INVX1 G40817 (.I(W1559), .ZN(W30503));
  INVX1 G40818 (.I(W2375), .ZN(W20288));
  INVX1 G40819 (.I(W3756), .ZN(W30501));
  INVX1 G40820 (.I(W408), .ZN(W30499));
  INVX1 G40821 (.I(W18027), .ZN(W30497));
  INVX1 G40822 (.I(W25854), .ZN(W30496));
  INVX1 G40823 (.I(W1620), .ZN(W30508));
  INVX1 G40824 (.I(W1289), .ZN(W20297));
  INVX1 G40825 (.I(W7259), .ZN(O5362));
  INVX1 G40826 (.I(W15615), .ZN(O5361));
  INVX1 G40827 (.I(I466), .ZN(W20302));
  INVX1 G40828 (.I(W25767), .ZN(O5357));
  INVX1 G40829 (.I(W23021), .ZN(O5356));
  INVX1 G40830 (.I(W2831), .ZN(O1972));
  INVX1 G40831 (.I(W20862), .ZN(O5355));
  INVX1 G40832 (.I(W20787), .ZN(W30476));
  INVX1 G40833 (.I(W2374), .ZN(W20272));
  INVX1 G40834 (.I(W19475), .ZN(W20265));
  INVX1 G40835 (.I(W5384), .ZN(W30530));
  INVX1 G40836 (.I(W12463), .ZN(W30529));
  INVX1 G40837 (.I(W7937), .ZN(W20267));
  INVX1 G40838 (.I(W28990), .ZN(O5379));
  INVX1 G40839 (.I(W14308), .ZN(W20270));
  INVX1 G40840 (.I(W1046), .ZN(O1966));
  INVX1 G40841 (.I(I1668), .ZN(W30524));
  INVX1 G40842 (.I(W2017), .ZN(O5378));
  INVX1 G40843 (.I(W11556), .ZN(O2008));
  INVX1 G40844 (.I(W19652), .ZN(O5377));
  INVX1 G40845 (.I(W7172), .ZN(W20273));
  INVX1 G40846 (.I(W7308), .ZN(W20274));
  INVX1 G40847 (.I(W25260), .ZN(O5374));
  INVX1 G40848 (.I(W2163), .ZN(W20276));
  INVX1 G40849 (.I(W23970), .ZN(W30514));
  INVX1 G40850 (.I(W19638), .ZN(O5371));
  INVX1 G40851 (.I(W10253), .ZN(W20280));
  INVX1 G40852 (.I(W19173), .ZN(O5368));
  INVX1 G40853 (.I(W6211), .ZN(W20603));
  INVX1 G40854 (.I(W18191), .ZN(O5230));
  INVX1 G40855 (.I(W4542), .ZN(W20588));
  INVX1 G40856 (.I(W20650), .ZN(O5228));
  INVX1 G40857 (.I(I1112), .ZN(O5226));
  INVX1 G40858 (.I(W5883), .ZN(W20596));
  INVX1 G40859 (.I(W4963), .ZN(W30196));
  INVX1 G40860 (.I(W5579), .ZN(W30193));
  INVX1 G40861 (.I(W3870), .ZN(W20599));
  INVX1 G40862 (.I(W14389), .ZN(O5222));
  INVX1 G40863 (.I(W7861), .ZN(W20602));
  INVX1 G40864 (.I(W16001), .ZN(O2038));
  INVX1 G40865 (.I(W18849), .ZN(O2041));
  INVX1 G40866 (.I(W18063), .ZN(O2042));
  INVX1 G40867 (.I(W12998), .ZN(W30183));
  INVX1 G40868 (.I(W5242), .ZN(O5217));
  INVX1 G40869 (.I(W5350), .ZN(W20608));
  INVX1 G40870 (.I(W18602), .ZN(W20611));
  INVX1 G40871 (.I(W9106), .ZN(O2043));
  INVX1 G40872 (.I(W13045), .ZN(O5214));
  INVX1 G40873 (.I(W10476), .ZN(W20616));
  INVX1 G40874 (.I(W3904), .ZN(O2033));
  INVX1 G40875 (.I(W14131), .ZN(O2028));
  INVX1 G40876 (.I(W1373), .ZN(O2029));
  INVX1 G40877 (.I(W12631), .ZN(O2030));
  INVX1 G40878 (.I(W28821), .ZN(W30232));
  INVX1 G40879 (.I(W28831), .ZN(W30227));
  INVX1 G40880 (.I(W24335), .ZN(O5241));
  INVX1 G40881 (.I(W1189), .ZN(O2032));
  INVX1 G40882 (.I(I910), .ZN(W20566));
  INVX1 G40883 (.I(W12667), .ZN(O5240));
  INVX1 G40884 (.I(W15117), .ZN(W20617));
  INVX1 G40885 (.I(W305), .ZN(O2034));
  INVX1 G40886 (.I(W6946), .ZN(O5237));
  INVX1 G40887 (.I(W2965), .ZN(W20572));
  INVX1 G40888 (.I(I1700), .ZN(O2036));
  INVX1 G40889 (.I(W3155), .ZN(W20576));
  INVX1 G40890 (.I(W3397), .ZN(O5234));
  INVX1 G40891 (.I(W16826), .ZN(W20580));
  INVX1 G40892 (.I(W13382), .ZN(W20582));
  INVX1 G40893 (.I(W7328), .ZN(W20584));
  INVX1 G40894 (.I(W3845), .ZN(W30132));
  INVX1 G40895 (.I(I1274), .ZN(W30144));
  INVX1 G40896 (.I(W19821), .ZN(O5202));
  INVX1 G40897 (.I(W28089), .ZN(W30142));
  INVX1 G40898 (.I(W1484), .ZN(W20637));
  INVX1 G40899 (.I(W12417), .ZN(W20638));
  INVX1 G40900 (.I(W6947), .ZN(W30139));
  INVX1 G40901 (.I(W4824), .ZN(W20642));
  INVX1 G40902 (.I(W13175), .ZN(O2049));
  INVX1 G40903 (.I(W12665), .ZN(W20650));
  INVX1 G40904 (.I(W19783), .ZN(W20635));
  INVX1 G40905 (.I(W9301), .ZN(W20651));
  INVX1 G40906 (.I(W12750), .ZN(O5198));
  INVX1 G40907 (.I(W13324), .ZN(W30128));
  INVX1 G40908 (.I(W26225), .ZN(O5197));
  INVX1 G40909 (.I(W19180), .ZN(O2051));
  INVX1 G40910 (.I(W2863), .ZN(W20659));
  INVX1 G40911 (.I(I79), .ZN(W30121));
  INVX1 G40912 (.I(W5594), .ZN(W30120));
  INVX1 G40913 (.I(W19995), .ZN(W30119));
  INVX1 G40914 (.I(W10717), .ZN(O2045));
  INVX1 G40915 (.I(W17814), .ZN(W30170));
  INVX1 G40916 (.I(W9540), .ZN(W20620));
  INVX1 G40917 (.I(W1819), .ZN(O5211));
  INVX1 G40918 (.I(W8067), .ZN(W30167));
  INVX1 G40919 (.I(W13523), .ZN(W30165));
  INVX1 G40920 (.I(W28873), .ZN(W30164));
  INVX1 G40921 (.I(W17038), .ZN(O5210));
  INVX1 G40922 (.I(W17075), .ZN(W20624));
  INVX1 G40923 (.I(W10091), .ZN(W30161));
  INVX1 G40924 (.I(W9174), .ZN(W20554));
  INVX1 G40925 (.I(W15577), .ZN(W20627));
  INVX1 G40926 (.I(W28791), .ZN(O5207));
  INVX1 G40927 (.I(W19725), .ZN(O2046));
  INVX1 G40928 (.I(W13311), .ZN(O2047));
  INVX1 G40929 (.I(W21317), .ZN(O5205));
  INVX1 G40930 (.I(W11536), .ZN(O5204));
  INVX1 G40931 (.I(W9405), .ZN(W30151));
  INVX1 G40932 (.I(W14583), .ZN(W20632));
  INVX1 G40933 (.I(W6348), .ZN(O5203));
  INVX1 G40934 (.I(W25588), .ZN(W30312));
  INVX1 G40935 (.I(W7255), .ZN(O5288));
  INVX1 G40936 (.I(W6602), .ZN(W20466));
  INVX1 G40937 (.I(W26294), .ZN(O5287));
  INVX1 G40938 (.I(W29132), .ZN(W30328));
  INVX1 G40939 (.I(W8409), .ZN(W20469));
  INVX1 G40940 (.I(W11255), .ZN(W30320));
  INVX1 G40941 (.I(W15390), .ZN(W20484));
  INVX1 G40942 (.I(W18540), .ZN(W20485));
  INVX1 G40943 (.I(W22747), .ZN(O5281));
  INVX1 G40944 (.I(W4288), .ZN(W20463));
  INVX1 G40945 (.I(W6109), .ZN(O5280));
  INVX1 G40946 (.I(W24019), .ZN(W30310));
  INVX1 G40947 (.I(W13619), .ZN(W30309));
  INVX1 G40948 (.I(W18403), .ZN(O2016));
  INVX1 G40949 (.I(I166), .ZN(W20488));
  INVX1 G40950 (.I(W4587), .ZN(W30304));
  INVX1 G40951 (.I(W6877), .ZN(W20492));
  INVX1 G40952 (.I(W22576), .ZN(O5278));
  INVX1 G40953 (.I(W11462), .ZN(W20494));
  INVX1 G40954 (.I(W7928), .ZN(W20445));
  INVX1 G40955 (.I(W7558), .ZN(W20425));
  INVX1 G40956 (.I(W11831), .ZN(W20426));
  INVX1 G40957 (.I(W14944), .ZN(W20427));
  INVX1 G40958 (.I(W19542), .ZN(W30357));
  INVX1 G40959 (.I(W12639), .ZN(W20438));
  INVX1 G40960 (.I(W8319), .ZN(W20439));
  INVX1 G40961 (.I(W18549), .ZN(W20443));
  INVX1 G40962 (.I(W4398), .ZN(W30351));
  INVX1 G40963 (.I(W1934), .ZN(O2010));
  INVX1 G40964 (.I(W478), .ZN(W20495));
  INVX1 G40965 (.I(W26309), .ZN(W30346));
  INVX1 G40966 (.I(W25680), .ZN(W30345));
  INVX1 G40967 (.I(W17372), .ZN(W20453));
  INVX1 G40968 (.I(W4801), .ZN(W30343));
  INVX1 G40969 (.I(W12073), .ZN(W20455));
  INVX1 G40970 (.I(W8547), .ZN(W20456));
  INVX1 G40971 (.I(W9523), .ZN(W20460));
  INVX1 G40972 (.I(W21091), .ZN(O5290));
  INVX1 G40973 (.I(W17624), .ZN(O2014));
  INVX1 G40974 (.I(W2094), .ZN(O2025));
  INVX1 G40975 (.I(W29945), .ZN(W30261));
  INVX1 G40976 (.I(W785), .ZN(W20533));
  INVX1 G40977 (.I(W14921), .ZN(W20534));
  INVX1 G40978 (.I(W20821), .ZN(O5258));
  INVX1 G40979 (.I(W3441), .ZN(O5257));
  INVX1 G40980 (.I(W12065), .ZN(W20537));
  INVX1 G40981 (.I(W26967), .ZN(O5256));
  INVX1 G40982 (.I(W15634), .ZN(W20538));
  INVX1 G40983 (.I(W5791), .ZN(W30252));
  INVX1 G40984 (.I(W6110), .ZN(W20527));
  INVX1 G40985 (.I(W209), .ZN(W30248));
  INVX1 G40986 (.I(W20357), .ZN(W20542));
  INVX1 G40987 (.I(W19525), .ZN(W20543));
  INVX1 G40988 (.I(W15022), .ZN(O2026));
  INVX1 G40989 (.I(I1927), .ZN(W30243));
  INVX1 G40990 (.I(W18258), .ZN(W20546));
  INVX1 G40991 (.I(I1459), .ZN(W20547));
  INVX1 G40992 (.I(W1393), .ZN(W20550));
  INVX1 G40993 (.I(W16351), .ZN(O5247));
  INVX1 G40994 (.I(W14257), .ZN(O5265));
  INVX1 G40995 (.I(W12424), .ZN(O5274));
  INVX1 G40996 (.I(W12424), .ZN(W30291));
  INVX1 G40997 (.I(W23518), .ZN(O5272));
  INVX1 G40998 (.I(W18631), .ZN(W30289));
  INVX1 G40999 (.I(W14075), .ZN(W20505));
  INVX1 G41000 (.I(W27624), .ZN(O5269));
  INVX1 G41001 (.I(W573), .ZN(O5268));
  INVX1 G41002 (.I(W6586), .ZN(W20508));
  INVX1 G41003 (.I(W12186), .ZN(W20510));
  INVX1 G41004 (.I(W11947), .ZN(W20209));
  INVX1 G41005 (.I(W11774), .ZN(O5264));
  INVX1 G41006 (.I(W19580), .ZN(O5263));
  INVX1 G41007 (.I(I1865), .ZN(W20511));
  INVX1 G41008 (.I(W14896), .ZN(W30273));
  INVX1 G41009 (.I(W19103), .ZN(W30272));
  INVX1 G41010 (.I(W14509), .ZN(W20515));
  INVX1 G41011 (.I(W13959), .ZN(W20524));
  INVX1 G41012 (.I(W19646), .ZN(W20526));
  INVX1 G41013 (.I(I68), .ZN(W30266));
  INVX1 G41014 (.I(W22149), .ZN(W30900));
  INVX1 G41015 (.I(W5895), .ZN(O5550));
  INVX1 G41016 (.I(W8513), .ZN(W30913));
  INVX1 G41017 (.I(W17215), .ZN(W30912));
  INVX1 G41018 (.I(W23363), .ZN(W30911));
  INVX1 G41019 (.I(W6715), .ZN(W30910));
  INVX1 G41020 (.I(W23065), .ZN(O5549));
  INVX1 G41021 (.I(W12205), .ZN(W30908));
  INVX1 G41022 (.I(W14031), .ZN(W30905));
  INVX1 G41023 (.I(W10569), .ZN(O5546));
  INVX1 G41024 (.I(W3135), .ZN(W19921));
  INVX1 G41025 (.I(W4464), .ZN(W19911));
  INVX1 G41026 (.I(W3569), .ZN(O5542));
  INVX1 G41027 (.I(W7873), .ZN(O5540));
  INVX1 G41028 (.I(W6247), .ZN(W19927));
  INVX1 G41029 (.I(W2300), .ZN(W30893));
  INVX1 G41030 (.I(W29695), .ZN(O5538));
  INVX1 G41031 (.I(W14166), .ZN(O5537));
  INVX1 G41032 (.I(W19502), .ZN(W19935));
  INVX1 G41033 (.I(W24063), .ZN(W30888));
  INVX1 G41034 (.I(W3306), .ZN(W19937));
  INVX1 G41035 (.I(W16565), .ZN(W30932));
  INVX1 G41036 (.I(W26179), .ZN(O5565));
  INVX1 G41037 (.I(W2412), .ZN(W19885));
  INVX1 G41038 (.I(W16607), .ZN(W19888));
  INVX1 G41039 (.I(W16195), .ZN(W19891));
  INVX1 G41040 (.I(W1102), .ZN(W19892));
  INVX1 G41041 (.I(W5136), .ZN(W19894));
  INVX1 G41042 (.I(W1361), .ZN(W30935));
  INVX1 G41043 (.I(W16236), .ZN(O1878));
  INVX1 G41044 (.I(W17609), .ZN(W30933));
  INVX1 G41045 (.I(W2938), .ZN(O1891));
  INVX1 G41046 (.I(W17655), .ZN(W19899));
  INVX1 G41047 (.I(W12401), .ZN(W19904));
  INVX1 G41048 (.I(W11193), .ZN(O5555));
  INVX1 G41049 (.I(W10527), .ZN(W30925));
  INVX1 G41050 (.I(W8766), .ZN(W19905));
  INVX1 G41051 (.I(W9337), .ZN(W19906));
  INVX1 G41052 (.I(W2826), .ZN(W19907));
  INVX1 G41053 (.I(W23899), .ZN(O5552));
  INVX1 G41054 (.I(W6995), .ZN(W19910));
  INVX1 G41055 (.I(W12000), .ZN(O5517));
  INVX1 G41056 (.I(W14138), .ZN(W19973));
  INVX1 G41057 (.I(I1503), .ZN(W19976));
  INVX1 G41058 (.I(I1264), .ZN(W19977));
  INVX1 G41059 (.I(W9931), .ZN(O1902));
  INVX1 G41060 (.I(W4662), .ZN(W30844));
  INVX1 G41061 (.I(W8555), .ZN(W30842));
  INVX1 G41062 (.I(W24324), .ZN(O5520));
  INVX1 G41063 (.I(W23185), .ZN(O5519));
  INVX1 G41064 (.I(W9451), .ZN(O1904));
  INVX1 G41065 (.I(W28322), .ZN(W30850));
  INVX1 G41066 (.I(W542), .ZN(O5516));
  INVX1 G41067 (.I(W10804), .ZN(W19983));
  INVX1 G41068 (.I(W2169), .ZN(W19984));
  INVX1 G41069 (.I(W8122), .ZN(W19986));
  INVX1 G41070 (.I(W12504), .ZN(W30832));
  INVX1 G41071 (.I(W16657), .ZN(W19987));
  INVX1 G41072 (.I(W13171), .ZN(W19988));
  INVX1 G41073 (.I(I1296), .ZN(W19990));
  INVX1 G41074 (.I(W25988), .ZN(W30827));
  INVX1 G41075 (.I(W16898), .ZN(W19957));
  INVX1 G41076 (.I(W13494), .ZN(W19943));
  INVX1 G41077 (.I(W30030), .ZN(O5531));
  INVX1 G41078 (.I(W13115), .ZN(O5530));
  INVX1 G41079 (.I(W15099), .ZN(W30876));
  INVX1 G41080 (.I(W14485), .ZN(W30874));
  INVX1 G41081 (.I(I811), .ZN(W30873));
  INVX1 G41082 (.I(W18780), .ZN(O5528));
  INVX1 G41083 (.I(W10067), .ZN(W19950));
  INVX1 G41084 (.I(W4437), .ZN(W19951));
  INVX1 G41085 (.I(W18726), .ZN(W19883));
  INVX1 G41086 (.I(W15104), .ZN(O5526));
  INVX1 G41087 (.I(W10320), .ZN(O1895));
  INVX1 G41088 (.I(W265), .ZN(W30862));
  INVX1 G41089 (.I(W19441), .ZN(O1897));
  INVX1 G41090 (.I(W28196), .ZN(W30857));
  INVX1 G41091 (.I(W184), .ZN(O1899));
  INVX1 G41092 (.I(W653), .ZN(W30853));
  INVX1 G41093 (.I(W16075), .ZN(O1901));
  INVX1 G41094 (.I(I1806), .ZN(W30851));
  INVX1 G41095 (.I(W22041), .ZN(W31023));
  INVX1 G41096 (.I(I723), .ZN(W31034));
  INVX1 G41097 (.I(W6818), .ZN(O1858));
  INVX1 G41098 (.I(I642), .ZN(W19801));
  INVX1 G41099 (.I(W11595), .ZN(O1859));
  INVX1 G41100 (.I(I1448), .ZN(O5610));
  INVX1 G41101 (.I(W10146), .ZN(W31027));
  INVX1 G41102 (.I(W19512), .ZN(W19804));
  INVX1 G41103 (.I(I1772), .ZN(W31025));
  INVX1 G41104 (.I(W6521), .ZN(O5608));
  INVX1 G41105 (.I(W6917), .ZN(W31036));
  INVX1 G41106 (.I(W19638), .ZN(W31019));
  INVX1 G41107 (.I(W3295), .ZN(W31018));
  INVX1 G41108 (.I(W30259), .ZN(O5606));
  INVX1 G41109 (.I(W13195), .ZN(W31015));
  INVX1 G41110 (.I(W19182), .ZN(O5605));
  INVX1 G41111 (.I(W6499), .ZN(W19810));
  INVX1 G41112 (.I(W16865), .ZN(W19811));
  INVX1 G41113 (.I(W10108), .ZN(W19812));
  INVX1 G41114 (.I(W13400), .ZN(W19823));
  INVX1 G41115 (.I(W2613), .ZN(O5623));
  INVX1 G41116 (.I(W30201), .ZN(W31058));
  INVX1 G41117 (.I(W5911), .ZN(W19782));
  INVX1 G41118 (.I(W2620), .ZN(W31055));
  INVX1 G41119 (.I(W16519), .ZN(W31054));
  INVX1 G41120 (.I(W93), .ZN(O1851));
  INVX1 G41121 (.I(W12516), .ZN(W31052));
  INVX1 G41122 (.I(W12751), .ZN(O1852));
  INVX1 G41123 (.I(W6747), .ZN(W19789));
  INVX1 G41124 (.I(W5027), .ZN(W19790));
  INVX1 G41125 (.I(W15191), .ZN(W19827));
  INVX1 G41126 (.I(W2908), .ZN(O5622));
  INVX1 G41127 (.I(W7129), .ZN(W19791));
  INVX1 G41128 (.I(W1497), .ZN(W19794));
  INVX1 G41129 (.I(W13807), .ZN(O1854));
  INVX1 G41130 (.I(W8284), .ZN(W31041));
  INVX1 G41131 (.I(W8924), .ZN(O1856));
  INVX1 G41132 (.I(W1990), .ZN(O5617));
  INVX1 G41133 (.I(I1634), .ZN(W31038));
  INVX1 G41134 (.I(W411), .ZN(O5616));
  INVX1 G41135 (.I(W3968), .ZN(O5576));
  INVX1 G41136 (.I(W22799), .ZN(O5583));
  INVX1 G41137 (.I(W16255), .ZN(W19849));
  INVX1 G41138 (.I(W14860), .ZN(W19851));
  INVX1 G41139 (.I(W15809), .ZN(W19854));
  INVX1 G41140 (.I(W9396), .ZN(W19856));
  INVX1 G41141 (.I(W28908), .ZN(O5580));
  INVX1 G41142 (.I(I1199), .ZN(O1868));
  INVX1 G41143 (.I(W1123), .ZN(O5578));
  INVX1 G41144 (.I(W1894), .ZN(W19860));
  INVX1 G41145 (.I(W7156), .ZN(W19846));
  INVX1 G41146 (.I(W3031), .ZN(W19863));
  INVX1 G41147 (.I(W14153), .ZN(W19864));
  INVX1 G41148 (.I(W19593), .ZN(W19868));
  INVX1 G41149 (.I(W8932), .ZN(O1872));
  INVX1 G41150 (.I(W15293), .ZN(W19871));
  INVX1 G41151 (.I(W897), .ZN(O1873));
  INVX1 G41152 (.I(W25010), .ZN(W30952));
  INVX1 G41153 (.I(W22085), .ZN(O5569));
  INVX1 G41154 (.I(W16262), .ZN(W19881));
  INVX1 G41155 (.I(W19286), .ZN(O1867));
  INVX1 G41156 (.I(W25695), .ZN(O5600));
  INVX1 G41157 (.I(W26556), .ZN(O5599));
  INVX1 G41158 (.I(W10712), .ZN(O5595));
  INVX1 G41159 (.I(I1049), .ZN(W30997));
  INVX1 G41160 (.I(W1281), .ZN(W19835));
  INVX1 G41161 (.I(W6341), .ZN(O1866));
  INVX1 G41162 (.I(W27321), .ZN(O5594));
  INVX1 G41163 (.I(W550), .ZN(W19841));
  INVX1 G41164 (.I(W8145), .ZN(W30991));
  INVX1 G41165 (.I(W14882), .ZN(W19992));
  INVX1 G41166 (.I(W20163), .ZN(O5590));
  INVX1 G41167 (.I(I57), .ZN(O5589));
  INVX1 G41168 (.I(W24418), .ZN(O5588));
  INVX1 G41169 (.I(W21759), .ZN(W30985));
  INVX1 G41170 (.I(W26106), .ZN(W30983));
  INVX1 G41171 (.I(W12844), .ZN(O5586));
  INVX1 G41172 (.I(W19972), .ZN(O5585));
  INVX1 G41173 (.I(W17191), .ZN(W19845));
  INVX1 G41174 (.I(W26401), .ZN(O5584));
  INVX1 G41175 (.I(W18763), .ZN(W20140));
  INVX1 G41176 (.I(W14905), .ZN(O5450));
  INVX1 G41177 (.I(W5294), .ZN(O5448));
  INVX1 G41178 (.I(W13754), .ZN(W20123));
  INVX1 G41179 (.I(I1159), .ZN(O1933));
  INVX1 G41180 (.I(W15018), .ZN(W30672));
  INVX1 G41181 (.I(W9022), .ZN(W20132));
  INVX1 G41182 (.I(W8143), .ZN(O5443));
  INVX1 G41183 (.I(W6395), .ZN(O1936));
  INVX1 G41184 (.I(W9874), .ZN(O1937));
  INVX1 G41185 (.I(W14651), .ZN(W20139));
  INVX1 G41186 (.I(W5999), .ZN(O5451));
  INVX1 G41187 (.I(W3573), .ZN(W20141));
  INVX1 G41188 (.I(W7303), .ZN(O1938));
  INVX1 G41189 (.I(W1264), .ZN(W20148));
  INVX1 G41190 (.I(W2469), .ZN(O5436));
  INVX1 G41191 (.I(W4115), .ZN(W20150));
  INVX1 G41192 (.I(W11218), .ZN(W30654));
  INVX1 G41193 (.I(W22218), .ZN(W30653));
  INVX1 G41194 (.I(W3289), .ZN(O5434));
  INVX1 G41195 (.I(W2599), .ZN(W20153));
  INVX1 G41196 (.I(W22560), .ZN(W30691));
  INVX1 G41197 (.I(W11250), .ZN(O1927));
  INVX1 G41198 (.I(W19414), .ZN(O5457));
  INVX1 G41199 (.I(W18086), .ZN(W30700));
  INVX1 G41200 (.I(W2691), .ZN(W30699));
  INVX1 G41201 (.I(W14873), .ZN(W20107));
  INVX1 G41202 (.I(I752), .ZN(W20110));
  INVX1 G41203 (.I(W14336), .ZN(O5454));
  INVX1 G41204 (.I(W18666), .ZN(O5452));
  INVX1 G41205 (.I(W13795), .ZN(W20113));
  INVX1 G41206 (.I(W1293), .ZN(O1941));
  INVX1 G41207 (.I(W17130), .ZN(W20114));
  INVX1 G41208 (.I(W3410), .ZN(W30689));
  INVX1 G41209 (.I(W2107), .ZN(W30688));
  INVX1 G41210 (.I(W28777), .ZN(W30687));
  INVX1 G41211 (.I(W4510), .ZN(W30686));
  INVX1 G41212 (.I(W12340), .ZN(W20115));
  INVX1 G41213 (.I(W2230), .ZN(W30684));
  INVX1 G41214 (.I(W18241), .ZN(W20117));
  INVX1 G41215 (.I(W27228), .ZN(W30682));
  INVX1 G41216 (.I(W23400), .ZN(O5412));
  INVX1 G41217 (.I(W1860), .ZN(W20183));
  INVX1 G41218 (.I(W24281), .ZN(W30617));
  INVX1 G41219 (.I(W19770), .ZN(W20184));
  INVX1 G41220 (.I(W11748), .ZN(W20187));
  INVX1 G41221 (.I(W12738), .ZN(W20188));
  INVX1 G41222 (.I(W11705), .ZN(W20189));
  INVX1 G41223 (.I(W15876), .ZN(W20191));
  INVX1 G41224 (.I(W9698), .ZN(W30607));
  INVX1 G41225 (.I(W12373), .ZN(W30606));
  INVX1 G41226 (.I(W7993), .ZN(W30619));
  INVX1 G41227 (.I(I753), .ZN(W20195));
  INVX1 G41228 (.I(W12797), .ZN(W30603));
  INVX1 G41229 (.I(I184), .ZN(O1950));
  INVX1 G41230 (.I(W6388), .ZN(W20198));
  INVX1 G41231 (.I(W1249), .ZN(W20199));
  INVX1 G41232 (.I(W6556), .ZN(W30597));
  INVX1 G41233 (.I(W3935), .ZN(O5407));
  INVX1 G41234 (.I(W14092), .ZN(O1953));
  INVX1 G41235 (.I(W2097), .ZN(O1955));
  INVX1 G41236 (.I(W2565), .ZN(W20168));
  INVX1 G41237 (.I(W14509), .ZN(W20155));
  INVX1 G41238 (.I(W14335), .ZN(W20158));
  INVX1 G41239 (.I(W14972), .ZN(W20159));
  INVX1 G41240 (.I(W15333), .ZN(W30642));
  INVX1 G41241 (.I(W21009), .ZN(O5426));
  INVX1 G41242 (.I(W15834), .ZN(W20161));
  INVX1 G41243 (.I(W11853), .ZN(W20165));
  INVX1 G41244 (.I(W11625), .ZN(O5423));
  INVX1 G41245 (.I(W18685), .ZN(O1945));
  INVX1 G41246 (.I(I1704), .ZN(W30704));
  INVX1 G41247 (.I(I1730), .ZN(W20170));
  INVX1 G41248 (.I(W11419), .ZN(W30631));
  INVX1 G41249 (.I(W3538), .ZN(O1947));
  INVX1 G41250 (.I(W19842), .ZN(O5420));
  INVX1 G41251 (.I(W19828), .ZN(W20179));
  INVX1 G41252 (.I(W121), .ZN(O5418));
  INVX1 G41253 (.I(W4826), .ZN(W30623));
  INVX1 G41254 (.I(W11302), .ZN(W20180));
  INVX1 G41255 (.I(W3289), .ZN(W20181));
  INVX1 G41256 (.I(W17898), .ZN(O5487));
  INVX1 G41257 (.I(W10765), .ZN(W20015));
  INVX1 G41258 (.I(W10835), .ZN(O5492));
  INVX1 G41259 (.I(I1894), .ZN(W20018));
  INVX1 G41260 (.I(W26896), .ZN(W30786));
  INVX1 G41261 (.I(W3386), .ZN(W20026));
  INVX1 G41262 (.I(W14405), .ZN(W20027));
  INVX1 G41263 (.I(W2461), .ZN(W20028));
  INVX1 G41264 (.I(W318), .ZN(W20030));
  INVX1 G41265 (.I(W17079), .ZN(W20033));
  INVX1 G41266 (.I(W13943), .ZN(W30797));
  INVX1 G41267 (.I(W8574), .ZN(O5485));
  INVX1 G41268 (.I(W6987), .ZN(W20036));
  INVX1 G41269 (.I(W6603), .ZN(W20040));
  INVX1 G41270 (.I(W26147), .ZN(W30771));
  INVX1 G41271 (.I(W7099), .ZN(W20042));
  INVX1 G41272 (.I(W12723), .ZN(O1913));
  INVX1 G41273 (.I(W11946), .ZN(O5481));
  INVX1 G41274 (.I(W26211), .ZN(O5480));
  INVX1 G41275 (.I(W16643), .ZN(W20052));
  INVX1 G41276 (.I(W15340), .ZN(W20010));
  INVX1 G41277 (.I(W10184), .ZN(W19993));
  INVX1 G41278 (.I(W1895), .ZN(O5508));
  INVX1 G41279 (.I(W27475), .ZN(W30822));
  INVX1 G41280 (.I(W7680), .ZN(W20000));
  INVX1 G41281 (.I(W12704), .ZN(W20002));
  INVX1 G41282 (.I(W2428), .ZN(W30818));
  INVX1 G41283 (.I(W15341), .ZN(O1906));
  INVX1 G41284 (.I(W2575), .ZN(O1907));
  INVX1 G41285 (.I(W10721), .ZN(W20007));
  INVX1 G41286 (.I(W8566), .ZN(W30759));
  INVX1 G41287 (.I(W21827), .ZN(O5500));
  INVX1 G41288 (.I(W19825), .ZN(O5499));
  INVX1 G41289 (.I(W16681), .ZN(W30806));
  INVX1 G41290 (.I(W8567), .ZN(W20012));
  INVX1 G41291 (.I(W27067), .ZN(W30804));
  INVX1 G41292 (.I(W29101), .ZN(W30802));
  INVX1 G41293 (.I(W24399), .ZN(O5497));
  INVX1 G41294 (.I(W11476), .ZN(O5496));
  INVX1 G41295 (.I(W17287), .ZN(O5495));
  INVX1 G41296 (.I(W64), .ZN(W20092));
  INVX1 G41297 (.I(W18685), .ZN(O1923));
  INVX1 G41298 (.I(W11311), .ZN(O1924));
  INVX1 G41299 (.I(W12429), .ZN(W30726));
  INVX1 G41300 (.I(W27586), .ZN(W30724));
  INVX1 G41301 (.I(W23728), .ZN(O5465));
  INVX1 G41302 (.I(W23288), .ZN(W30722));
  INVX1 G41303 (.I(W28941), .ZN(O5464));
  INVX1 G41304 (.I(W3561), .ZN(W20089));
  INVX1 G41305 (.I(W18132), .ZN(W20090));
  INVX1 G41306 (.I(W17108), .ZN(W20080));
  INVX1 G41307 (.I(W3959), .ZN(W20094));
  INVX1 G41308 (.I(W10742), .ZN(W30715));
  INVX1 G41309 (.I(I1398), .ZN(O5461));
  INVX1 G41310 (.I(W18034), .ZN(W30712));
  INVX1 G41311 (.I(W13178), .ZN(W20096));
  INVX1 G41312 (.I(W12245), .ZN(W20098));
  INVX1 G41313 (.I(I500), .ZN(W30708));
  INVX1 G41314 (.I(W7248), .ZN(W20100));
  INVX1 G41315 (.I(W93), .ZN(W20101));
  INVX1 G41316 (.I(I620), .ZN(W20068));
  INVX1 G41317 (.I(W3862), .ZN(W30758));
  INVX1 G41318 (.I(W20546), .ZN(W30756));
  INVX1 G41319 (.I(W29495), .ZN(O5478));
  INVX1 G41320 (.I(W13135), .ZN(W30753));
  INVX1 G41321 (.I(W280), .ZN(W30752));
  INVX1 G41322 (.I(W1010), .ZN(W20063));
  INVX1 G41323 (.I(W6100), .ZN(W20065));
  INVX1 G41324 (.I(I1883), .ZN(W20066));
  INVX1 G41325 (.I(W18518), .ZN(O1920));
  INVX1 G41326 (.I(W10567), .ZN(W20663));
  INVX1 G41327 (.I(W22630), .ZN(W30742));
  INVX1 G41328 (.I(W2698), .ZN(W20069));
  INVX1 G41329 (.I(I1353), .ZN(W20071));
  INVX1 G41330 (.I(W19134), .ZN(W20072));
  INVX1 G41331 (.I(W27676), .ZN(W30738));
  INVX1 G41332 (.I(W19805), .ZN(W30735));
  INVX1 G41333 (.I(W13211), .ZN(O1921));
  INVX1 G41334 (.I(W15409), .ZN(W30732));
  INVX1 G41335 (.I(W25555), .ZN(O5468));
  INVX1 G41336 (.I(W13882), .ZN(W21299));
  INVX1 G41337 (.I(W21215), .ZN(O2202));
  INVX1 G41338 (.I(W9841), .ZN(O2203));
  INVX1 G41339 (.I(W23707), .ZN(W29481));
  INVX1 G41340 (.I(W16899), .ZN(W21288));
  INVX1 G41341 (.I(I723), .ZN(O4915));
  INVX1 G41342 (.I(W7564), .ZN(O2204));
  INVX1 G41343 (.I(W26790), .ZN(W29475));
  INVX1 G41344 (.I(W16047), .ZN(O4912));
  INVX1 G41345 (.I(W29388), .ZN(O4911));
  INVX1 G41346 (.I(W14556), .ZN(O4910));
  INVX1 G41347 (.I(W9795), .ZN(W21279));
  INVX1 G41348 (.I(W6204), .ZN(O2208));
  INVX1 G41349 (.I(W10424), .ZN(O2209));
  INVX1 G41350 (.I(W25207), .ZN(O4905));
  INVX1 G41351 (.I(W71), .ZN(W21309));
  INVX1 G41352 (.I(W16754), .ZN(O4903));
  INVX1 G41353 (.I(W7844), .ZN(W29458));
  INVX1 G41354 (.I(I471), .ZN(O2212));
  INVX1 G41355 (.I(W7976), .ZN(O2213));
  INVX1 G41356 (.I(W9608), .ZN(W21314));
  INVX1 G41357 (.I(W19889), .ZN(W21260));
  INVX1 G41358 (.I(W9366), .ZN(W21248));
  INVX1 G41359 (.I(W20582), .ZN(W29512));
  INVX1 G41360 (.I(W8863), .ZN(W21251));
  INVX1 G41361 (.I(W4450), .ZN(W21252));
  INVX1 G41362 (.I(W10946), .ZN(O4925));
  INVX1 G41363 (.I(W4639), .ZN(W21256));
  INVX1 G41364 (.I(W24696), .ZN(O4924));
  INVX1 G41365 (.I(W3508), .ZN(W29504));
  INVX1 G41366 (.I(W29107), .ZN(W29502));
  INVX1 G41367 (.I(W11166), .ZN(W21316));
  INVX1 G41368 (.I(W12027), .ZN(W21263));
  INVX1 G41369 (.I(W19608), .ZN(W21265));
  INVX1 G41370 (.I(W15646), .ZN(W29494));
  INVX1 G41371 (.I(W18326), .ZN(W29493));
  INVX1 G41372 (.I(W25725), .ZN(O4920));
  INVX1 G41373 (.I(W18481), .ZN(O2198));
  INVX1 G41374 (.I(W9187), .ZN(W29489));
  INVX1 G41375 (.I(I540), .ZN(W21277));
  INVX1 G41376 (.I(W8893), .ZN(W29486));
  INVX1 G41377 (.I(W11964), .ZN(W21367));
  INVX1 G41378 (.I(W12469), .ZN(O4885));
  INVX1 G41379 (.I(I422), .ZN(O2222));
  INVX1 G41380 (.I(W1903), .ZN(O2223));
  INVX1 G41381 (.I(W17044), .ZN(O2225));
  INVX1 G41382 (.I(W17090), .ZN(W21363));
  INVX1 G41383 (.I(W5919), .ZN(O4882));
  INVX1 G41384 (.I(W4184), .ZN(W21365));
  INVX1 G41385 (.I(W11095), .ZN(O2226));
  INVX1 G41386 (.I(W10369), .ZN(O4878));
  INVX1 G41387 (.I(W26367), .ZN(W29425));
  INVX1 G41388 (.I(W20669), .ZN(W29409));
  INVX1 G41389 (.I(W6849), .ZN(W29408));
  INVX1 G41390 (.I(W11664), .ZN(W21368));
  INVX1 G41391 (.I(W28692), .ZN(W29406));
  INVX1 G41392 (.I(W11390), .ZN(W21371));
  INVX1 G41393 (.I(W5717), .ZN(W29402));
  INVX1 G41394 (.I(W8586), .ZN(W21375));
  INVX1 G41395 (.I(W12970), .ZN(W21377));
  INVX1 G41396 (.I(W6976), .ZN(W29397));
  INVX1 G41397 (.I(W11989), .ZN(W21328));
  INVX1 G41398 (.I(W1613), .ZN(W21317));
  INVX1 G41399 (.I(W9675), .ZN(O2214));
  INVX1 G41400 (.I(W6019), .ZN(W21319));
  INVX1 G41401 (.I(W10282), .ZN(W21320));
  INVX1 G41402 (.I(W8600), .ZN(O2215));
  INVX1 G41403 (.I(W18323), .ZN(W21323));
  INVX1 G41404 (.I(W3838), .ZN(W21324));
  INVX1 G41405 (.I(W19868), .ZN(W21325));
  INVX1 G41406 (.I(W370), .ZN(W21326));
  INVX1 G41407 (.I(W15866), .ZN(W21247));
  INVX1 G41408 (.I(I928), .ZN(W29439));
  INVX1 G41409 (.I(W12862), .ZN(O2217));
  INVX1 G41410 (.I(W4121), .ZN(O2218));
  INVX1 G41411 (.I(W8445), .ZN(W21341));
  INVX1 G41412 (.I(W7692), .ZN(O4888));
  INVX1 G41413 (.I(W27448), .ZN(O4887));
  INVX1 G41414 (.I(W8844), .ZN(O2219));
  INVX1 G41415 (.I(W10849), .ZN(W21348));
  INVX1 G41416 (.I(W19228), .ZN(W21349));
  INVX1 G41417 (.I(W4129), .ZN(W21178));
  INVX1 G41418 (.I(W559), .ZN(O2168));
  INVX1 G41419 (.I(W16627), .ZN(W29599));
  INVX1 G41420 (.I(W1644), .ZN(O2169));
  INVX1 G41421 (.I(W19111), .ZN(O4964));
  INVX1 G41422 (.I(W11398), .ZN(O4963));
  INVX1 G41423 (.I(W21007), .ZN(O2171));
  INVX1 G41424 (.I(W18917), .ZN(W29588));
  INVX1 G41425 (.I(W19765), .ZN(W29587));
  INVX1 G41426 (.I(W3031), .ZN(W29586));
  INVX1 G41427 (.I(W1497), .ZN(O2167));
  INVX1 G41428 (.I(W5876), .ZN(W29584));
  INVX1 G41429 (.I(W17334), .ZN(W29580));
  INVX1 G41430 (.I(W586), .ZN(W21182));
  INVX1 G41431 (.I(W16176), .ZN(W21184));
  INVX1 G41432 (.I(W6818), .ZN(W29576));
  INVX1 G41433 (.I(W1874), .ZN(W29575));
  INVX1 G41434 (.I(W20108), .ZN(O2173));
  INVX1 G41435 (.I(W21092), .ZN(W29573));
  INVX1 G41436 (.I(I85), .ZN(W21187));
  INVX1 G41437 (.I(W2344), .ZN(W21146));
  INVX1 G41438 (.I(W1485), .ZN(O4981));
  INVX1 G41439 (.I(W14514), .ZN(W29630));
  INVX1 G41440 (.I(W8751), .ZN(W21135));
  INVX1 G41441 (.I(W3904), .ZN(W29627));
  INVX1 G41442 (.I(W6519), .ZN(O2157));
  INVX1 G41443 (.I(W624), .ZN(O2159));
  INVX1 G41444 (.I(W20938), .ZN(W21140));
  INVX1 G41445 (.I(W8411), .ZN(W29621));
  INVX1 G41446 (.I(W11275), .ZN(O4976));
  INVX1 G41447 (.I(W12829), .ZN(W29571));
  INVX1 G41448 (.I(W12151), .ZN(W21148));
  INVX1 G41449 (.I(W15868), .ZN(O2162));
  INVX1 G41450 (.I(W14736), .ZN(W21153));
  INVX1 G41451 (.I(W8974), .ZN(W21154));
  INVX1 G41452 (.I(W16412), .ZN(O4971));
  INVX1 G41453 (.I(W3782), .ZN(W29608));
  INVX1 G41454 (.I(W7598), .ZN(O4969));
  INVX1 G41455 (.I(I1428), .ZN(O4968));
  INVX1 G41456 (.I(W13623), .ZN(O2165));
  INVX1 G41457 (.I(W2246), .ZN(W21238));
  INVX1 G41458 (.I(W16578), .ZN(W21223));
  INVX1 G41459 (.I(W1622), .ZN(O2188));
  INVX1 G41460 (.I(W8939), .ZN(W21230));
  INVX1 G41461 (.I(W20584), .ZN(W29534));
  INVX1 G41462 (.I(W19965), .ZN(O2190));
  INVX1 G41463 (.I(W25242), .ZN(O4940));
  INVX1 G41464 (.I(W10859), .ZN(W21233));
  INVX1 G41465 (.I(W13708), .ZN(W29530));
  INVX1 G41466 (.I(W18083), .ZN(W21237));
  INVX1 G41467 (.I(W9379), .ZN(W21222));
  INVX1 G41468 (.I(W3778), .ZN(W29526));
  INVX1 G41469 (.I(W7259), .ZN(W21240));
  INVX1 G41470 (.I(W827), .ZN(W29523));
  INVX1 G41471 (.I(W16532), .ZN(O4934));
  INVX1 G41472 (.I(W2132), .ZN(W29521));
  INVX1 G41473 (.I(W13856), .ZN(O4933));
  INVX1 G41474 (.I(W19098), .ZN(W21242));
  INVX1 G41475 (.I(W991), .ZN(W21244));
  INVX1 G41476 (.I(W20451), .ZN(W21246));
  INVX1 G41477 (.I(W15303), .ZN(W21207));
  INVX1 G41478 (.I(W5884), .ZN(O2176));
  INVX1 G41479 (.I(W5114), .ZN(O2178));
  INVX1 G41480 (.I(W19121), .ZN(W21195));
  INVX1 G41481 (.I(I237), .ZN(O4953));
  INVX1 G41482 (.I(W9677), .ZN(W21199));
  INVX1 G41483 (.I(W8134), .ZN(W29562));
  INVX1 G41484 (.I(I1370), .ZN(W21202));
  INVX1 G41485 (.I(W26074), .ZN(W29558));
  INVX1 G41486 (.I(W8062), .ZN(W29557));
  INVX1 G41487 (.I(W7994), .ZN(O4871));
  INVX1 G41488 (.I(W9780), .ZN(W21209));
  INVX1 G41489 (.I(W20985), .ZN(O4947));
  INVX1 G41490 (.I(W14400), .ZN(W21210));
  INVX1 G41491 (.I(W11893), .ZN(W29549));
  INVX1 G41492 (.I(W3124), .ZN(O2184));
  INVX1 G41493 (.I(W26416), .ZN(W29547));
  INVX1 G41494 (.I(W5214), .ZN(W21215));
  INVX1 G41495 (.I(W4618), .ZN(W21217));
  INVX1 G41496 (.I(W4106), .ZN(O4945));
  INVX1 G41497 (.I(W13228), .ZN(W21522));
  INVX1 G41498 (.I(W9988), .ZN(W21512));
  INVX1 G41499 (.I(W10858), .ZN(O2267));
  INVX1 G41500 (.I(W5038), .ZN(O2268));
  INVX1 G41501 (.I(W21856), .ZN(O4808));
  INVX1 G41502 (.I(W7947), .ZN(W21516));
  INVX1 G41503 (.I(W5809), .ZN(W21518));
  INVX1 G41504 (.I(W17645), .ZN(W21520));
  INVX1 G41505 (.I(W26602), .ZN(W29255));
  INVX1 G41506 (.I(W23067), .ZN(O4806));
  INVX1 G41507 (.I(W27596), .ZN(O4805));
  INVX1 G41508 (.I(W13381), .ZN(O2265));
  INVX1 G41509 (.I(W15095), .ZN(W29249));
  INVX1 G41510 (.I(W13067), .ZN(W21526));
  INVX1 G41511 (.I(W25645), .ZN(W29247));
  INVX1 G41512 (.I(W16367), .ZN(W21527));
  INVX1 G41513 (.I(W4309), .ZN(O2272));
  INVX1 G41514 (.I(W14077), .ZN(W21535));
  INVX1 G41515 (.I(W457), .ZN(W29242));
  INVX1 G41516 (.I(W17435), .ZN(O2274));
  INVX1 G41517 (.I(W21264), .ZN(W21540));
  INVX1 G41518 (.I(W4823), .ZN(W21493));
  INVX1 G41519 (.I(W15683), .ZN(W21486));
  INVX1 G41520 (.I(W16180), .ZN(W29290));
  INVX1 G41521 (.I(W268), .ZN(O2257));
  INVX1 G41522 (.I(W14308), .ZN(O4817));
  INVX1 G41523 (.I(W3078), .ZN(W21489));
  INVX1 G41524 (.I(W3235), .ZN(W21492));
  INVX1 G41525 (.I(W18390), .ZN(O4816));
  INVX1 G41526 (.I(W2301), .ZN(W29284));
  INVX1 G41527 (.I(W29222), .ZN(W29283));
  INVX1 G41528 (.I(I1301), .ZN(O4801));
  INVX1 G41529 (.I(W20423), .ZN(W21495));
  INVX1 G41530 (.I(W12370), .ZN(W29279));
  INVX1 G41531 (.I(W14811), .ZN(W29278));
  INVX1 G41532 (.I(W12980), .ZN(O2259));
  INVX1 G41533 (.I(W10193), .ZN(W21499));
  INVX1 G41534 (.I(W5306), .ZN(O2262));
  INVX1 G41535 (.I(W21615), .ZN(O4813));
  INVX1 G41536 (.I(W11082), .ZN(W21505));
  INVX1 G41537 (.I(W5312), .ZN(W21507));
  INVX1 G41538 (.I(W14342), .ZN(W21584));
  INVX1 G41539 (.I(W6919), .ZN(W29211));
  INVX1 G41540 (.I(W5446), .ZN(W21567));
  INVX1 G41541 (.I(W16048), .ZN(W21569));
  INVX1 G41542 (.I(W1969), .ZN(O2284));
  INVX1 G41543 (.I(W3407), .ZN(O2286));
  INVX1 G41544 (.I(W10549), .ZN(W29200));
  INVX1 G41545 (.I(I267), .ZN(O4787));
  INVX1 G41546 (.I(W2390), .ZN(W21582));
  INVX1 G41547 (.I(W8853), .ZN(W21583));
  INVX1 G41548 (.I(I1672), .ZN(W29212));
  INVX1 G41549 (.I(I1507), .ZN(W29195));
  INVX1 G41550 (.I(I698), .ZN(O2287));
  INVX1 G41551 (.I(W15635), .ZN(W29190));
  INVX1 G41552 (.I(W16738), .ZN(O2288));
  INVX1 G41553 (.I(W7148), .ZN(O2289));
  INVX1 G41554 (.I(W6637), .ZN(O2290));
  INVX1 G41555 (.I(I640), .ZN(W21598));
  INVX1 G41556 (.I(I1375), .ZN(W21599));
  INVX1 G41557 (.I(I365), .ZN(O4781));
  INVX1 G41558 (.I(W10944), .ZN(W21550));
  INVX1 G41559 (.I(W27726), .ZN(O4799));
  INVX1 G41560 (.I(W13194), .ZN(W29231));
  INVX1 G41561 (.I(W15604), .ZN(O2275));
  INVX1 G41562 (.I(W9795), .ZN(O2276));
  INVX1 G41563 (.I(W3027), .ZN(O2277));
  INVX1 G41564 (.I(W7901), .ZN(W21549));
  INVX1 G41565 (.I(W14460), .ZN(O4794));
  INVX1 G41566 (.I(W23729), .ZN(W29225));
  INVX1 G41567 (.I(W25954), .ZN(W29224));
  INVX1 G41568 (.I(W9619), .ZN(O4820));
  INVX1 G41569 (.I(W2285), .ZN(O2278));
  INVX1 G41570 (.I(W10357), .ZN(W21553));
  INVX1 G41571 (.I(W5096), .ZN(W21554));
  INVX1 G41572 (.I(W11966), .ZN(O2279));
  INVX1 G41573 (.I(W11251), .ZN(W21557));
  INVX1 G41574 (.I(W13798), .ZN(W21560));
  INVX1 G41575 (.I(W17224), .ZN(O2280));
  INVX1 G41576 (.I(W6613), .ZN(O4790));
  INVX1 G41577 (.I(W23770), .ZN(W29213));
  INVX1 G41578 (.I(W7690), .ZN(W21423));
  INVX1 G41579 (.I(W1479), .ZN(W29366));
  INVX1 G41580 (.I(W9821), .ZN(O2238));
  INVX1 G41581 (.I(W4725), .ZN(O4858));
  INVX1 G41582 (.I(W11190), .ZN(W21411));
  INVX1 G41583 (.I(W25736), .ZN(W29361));
  INVX1 G41584 (.I(W3931), .ZN(W21412));
  INVX1 G41585 (.I(W9774), .ZN(W21417));
  INVX1 G41586 (.I(W4279), .ZN(O2241));
  INVX1 G41587 (.I(W15247), .ZN(W21420));
  INVX1 G41588 (.I(W1212), .ZN(W29368));
  INVX1 G41589 (.I(W8485), .ZN(O2243));
  INVX1 G41590 (.I(W20607), .ZN(O4853));
  INVX1 G41591 (.I(W21170), .ZN(O2244));
  INVX1 G41592 (.I(W13861), .ZN(O4851));
  INVX1 G41593 (.I(W11684), .ZN(W21432));
  INVX1 G41594 (.I(W18130), .ZN(W21433));
  INVX1 G41595 (.I(W7675), .ZN(W29346));
  INVX1 G41596 (.I(W13428), .ZN(O4847));
  INVX1 G41597 (.I(W10754), .ZN(W21435));
  INVX1 G41598 (.I(W7815), .ZN(O2235));
  INVX1 G41599 (.I(W7466), .ZN(W21382));
  INVX1 G41600 (.I(W5618), .ZN(W21383));
  INVX1 G41601 (.I(W9992), .ZN(O2229));
  INVX1 G41602 (.I(W18725), .ZN(W21386));
  INVX1 G41603 (.I(W5242), .ZN(O2232));
  INVX1 G41604 (.I(W28757), .ZN(W29388));
  INVX1 G41605 (.I(W8951), .ZN(W21392));
  INVX1 G41606 (.I(W350), .ZN(O4868));
  INVX1 G41607 (.I(W3855), .ZN(W21395));
  INVX1 G41608 (.I(I1030), .ZN(W21437));
  INVX1 G41609 (.I(W27326), .ZN(W29381));
  INVX1 G41610 (.I(W2127), .ZN(W29380));
  INVX1 G41611 (.I(W10313), .ZN(W29379));
  INVX1 G41612 (.I(W4423), .ZN(W21401));
  INVX1 G41613 (.I(W19113), .ZN(O4863));
  INVX1 G41614 (.I(W3624), .ZN(W21406));
  INVX1 G41615 (.I(W19130), .ZN(O4862));
  INVX1 G41616 (.I(W5878), .ZN(W21407));
  INVX1 G41617 (.I(W21721), .ZN(O4861));
  INVX1 G41618 (.I(W422), .ZN(W21475));
  INVX1 G41619 (.I(W22815), .ZN(O4830));
  INVX1 G41620 (.I(W23738), .ZN(W29316));
  INVX1 G41621 (.I(W10746), .ZN(W29310));
  INVX1 G41622 (.I(W6090), .ZN(O2251));
  INVX1 G41623 (.I(W17539), .ZN(W21471));
  INVX1 G41624 (.I(W8858), .ZN(O4826));
  INVX1 G41625 (.I(W23524), .ZN(O4825));
  INVX1 G41626 (.I(W5157), .ZN(W21473));
  INVX1 G41627 (.I(W21225), .ZN(O2253));
  INVX1 G41628 (.I(I813), .ZN(W29318));
  INVX1 G41629 (.I(W9002), .ZN(W21476));
  INVX1 G41630 (.I(W16982), .ZN(W21478));
  INVX1 G41631 (.I(W24159), .ZN(W29300));
  INVX1 G41632 (.I(W3726), .ZN(W21479));
  INVX1 G41633 (.I(I781), .ZN(O2255));
  INVX1 G41634 (.I(W19702), .ZN(W21482));
  INVX1 G41635 (.I(W7694), .ZN(W21483));
  INVX1 G41636 (.I(W20215), .ZN(W21484));
  INVX1 G41637 (.I(W16251), .ZN(O2256));
  INVX1 G41638 (.I(W21351), .ZN(W21451));
  INVX1 G41639 (.I(W14656), .ZN(O2245));
  INVX1 G41640 (.I(W2666), .ZN(W21440));
  INVX1 G41641 (.I(W3937), .ZN(W21442));
  INVX1 G41642 (.I(W16909), .ZN(O4841));
  INVX1 G41643 (.I(W17140), .ZN(W21443));
  INVX1 G41644 (.I(W18402), .ZN(O4840));
  INVX1 G41645 (.I(W381), .ZN(W29334));
  INVX1 G41646 (.I(W15520), .ZN(O2247));
  INVX1 G41647 (.I(W20885), .ZN(W21450));
  INVX1 G41648 (.I(W19302), .ZN(W21130));
  INVX1 G41649 (.I(W13769), .ZN(O4838));
  INVX1 G41650 (.I(I917), .ZN(W21452));
  INVX1 G41651 (.I(W4540), .ZN(W21453));
  INVX1 G41652 (.I(W18475), .ZN(O4836));
  INVX1 G41653 (.I(W4429), .ZN(W21458));
  INVX1 G41654 (.I(I481), .ZN(O4833));
  INVX1 G41655 (.I(W10781), .ZN(W21460));
  INVX1 G41656 (.I(W3156), .ZN(W21461));
  INVX1 G41657 (.I(W831), .ZN(O2249));
  INVX1 G41658 (.I(W17623), .ZN(W20806));
  INVX1 G41659 (.I(W21239), .ZN(O5130));
  INVX1 G41660 (.I(W23852), .ZN(W29966));
  INVX1 G41661 (.I(W13567), .ZN(W20795));
  INVX1 G41662 (.I(W4124), .ZN(W20797));
  INVX1 G41663 (.I(W11043), .ZN(O5128));
  INVX1 G41664 (.I(W17026), .ZN(O5127));
  INVX1 G41665 (.I(W5514), .ZN(W20798));
  INVX1 G41666 (.I(W8296), .ZN(W20799));
  INVX1 G41667 (.I(W14588), .ZN(W20804));
  INVX1 G41668 (.I(W4480), .ZN(W29957));
  INVX1 G41669 (.I(W7667), .ZN(W20793));
  INVX1 G41670 (.I(W20519), .ZN(W20807));
  INVX1 G41671 (.I(W4788), .ZN(O2086));
  INVX1 G41672 (.I(W5973), .ZN(W20811));
  INVX1 G41673 (.I(W23223), .ZN(O5124));
  INVX1 G41674 (.I(W8688), .ZN(O5122));
  INVX1 G41675 (.I(W14154), .ZN(W29947));
  INVX1 G41676 (.I(W21004), .ZN(O5120));
  INVX1 G41677 (.I(W292), .ZN(W20829));
  INVX1 G41678 (.I(W9687), .ZN(W20830));
  INVX1 G41679 (.I(W21596), .ZN(W29978));
  INVX1 G41680 (.I(W4879), .ZN(O2079));
  INVX1 G41681 (.I(W23404), .ZN(W29988));
  INVX1 G41682 (.I(W18179), .ZN(W29987));
  INVX1 G41683 (.I(W19468), .ZN(W29986));
  INVX1 G41684 (.I(W14666), .ZN(O5141));
  INVX1 G41685 (.I(W15326), .ZN(W20782));
  INVX1 G41686 (.I(W15630), .ZN(O2083));
  INVX1 G41687 (.I(W11866), .ZN(W20787));
  INVX1 G41688 (.I(W119), .ZN(O5138));
  INVX1 G41689 (.I(W415), .ZN(W29940));
  INVX1 G41690 (.I(I1880), .ZN(W20788));
  INVX1 G41691 (.I(W17831), .ZN(O2084));
  INVX1 G41692 (.I(W20577), .ZN(O5137));
  INVX1 G41693 (.I(W12776), .ZN(O5136));
  INVX1 G41694 (.I(W28709), .ZN(O5135));
  INVX1 G41695 (.I(W16788), .ZN(W20790));
  INVX1 G41696 (.I(W13249), .ZN(W29971));
  INVX1 G41697 (.I(W7876), .ZN(W20791));
  INVX1 G41698 (.I(W18228), .ZN(O5132));
  INVX1 G41699 (.I(W6079), .ZN(W20868));
  INVX1 G41700 (.I(W11657), .ZN(W20861));
  INVX1 G41701 (.I(W6807), .ZN(W20862));
  INVX1 G41702 (.I(W24121), .ZN(O5102));
  INVX1 G41703 (.I(W3758), .ZN(W20863));
  INVX1 G41704 (.I(W8918), .ZN(O2101));
  INVX1 G41705 (.I(W4), .ZN(O5100));
  INVX1 G41706 (.I(W5127), .ZN(W20865));
  INVX1 G41707 (.I(I1529), .ZN(O2103));
  INVX1 G41708 (.I(W717), .ZN(W29900));
  INVX1 G41709 (.I(W22816), .ZN(O5104));
  INVX1 G41710 (.I(W29239), .ZN(W29898));
  INVX1 G41711 (.I(W8513), .ZN(O5098));
  INVX1 G41712 (.I(W15265), .ZN(W29895));
  INVX1 G41713 (.I(W7337), .ZN(W20871));
  INVX1 G41714 (.I(W1299), .ZN(W20872));
  INVX1 G41715 (.I(W8783), .ZN(W20873));
  INVX1 G41716 (.I(W3858), .ZN(O5096));
  INVX1 G41717 (.I(W27997), .ZN(O5095));
  INVX1 G41718 (.I(W4408), .ZN(W20879));
  INVX1 G41719 (.I(W14961), .ZN(W29923));
  INVX1 G41720 (.I(W853), .ZN(W29939));
  INVX1 G41721 (.I(W19688), .ZN(O2095));
  INVX1 G41722 (.I(W4519), .ZN(W20836));
  INVX1 G41723 (.I(W15988), .ZN(W20837));
  INVX1 G41724 (.I(W11008), .ZN(W20839));
  INVX1 G41725 (.I(W8869), .ZN(W20840));
  INVX1 G41726 (.I(W26406), .ZN(W29926));
  INVX1 G41727 (.I(W2952), .ZN(W29925));
  INVX1 G41728 (.I(W22875), .ZN(W29924));
  INVX1 G41729 (.I(W18048), .ZN(O2078));
  INVX1 G41730 (.I(I1876), .ZN(O2099));
  INVX1 G41731 (.I(W7899), .ZN(W20852));
  INVX1 G41732 (.I(W20911), .ZN(O5109));
  INVX1 G41733 (.I(W4788), .ZN(O2100));
  INVX1 G41734 (.I(W1942), .ZN(W29916));
  INVX1 G41735 (.I(W8441), .ZN(O5107));
  INVX1 G41736 (.I(W14249), .ZN(W20856));
  INVX1 G41737 (.I(W19574), .ZN(W20858));
  INVX1 G41738 (.I(W4346), .ZN(O5105));
  INVX1 G41739 (.I(W10940), .ZN(W30076));
  INVX1 G41740 (.I(W8572), .ZN(W20690));
  INVX1 G41741 (.I(W1467), .ZN(W30086));
  INVX1 G41742 (.I(W10516), .ZN(W30085));
  INVX1 G41743 (.I(W29742), .ZN(W30084));
  INVX1 G41744 (.I(W19159), .ZN(W30083));
  INVX1 G41745 (.I(I276), .ZN(W20692));
  INVX1 G41746 (.I(W14969), .ZN(O2059));
  INVX1 G41747 (.I(I43), .ZN(O5182));
  INVX1 G41748 (.I(W13135), .ZN(W30077));
  INVX1 G41749 (.I(W19564), .ZN(W20689));
  INVX1 G41750 (.I(W1456), .ZN(W20696));
  INVX1 G41751 (.I(W7623), .ZN(W20698));
  INVX1 G41752 (.I(W1550), .ZN(W20700));
  INVX1 G41753 (.I(W7801), .ZN(W30070));
  INVX1 G41754 (.I(W11506), .ZN(W20701));
  INVX1 G41755 (.I(W27084), .ZN(W30067));
  INVX1 G41756 (.I(W335), .ZN(W20708));
  INVX1 G41757 (.I(W23749), .ZN(O5176));
  INVX1 G41758 (.I(W17532), .ZN(O5175));
  INVX1 G41759 (.I(W11648), .ZN(W30105));
  INVX1 G41760 (.I(W16344), .ZN(O5194));
  INVX1 G41761 (.I(W7648), .ZN(W30116));
  INVX1 G41762 (.I(W2819), .ZN(W20668));
  INVX1 G41763 (.I(W8510), .ZN(O2053));
  INVX1 G41764 (.I(W22462), .ZN(W30111));
  INVX1 G41765 (.I(I1075), .ZN(W20671));
  INVX1 G41766 (.I(W10731), .ZN(W20672));
  INVX1 G41767 (.I(W20018), .ZN(W30108));
  INVX1 G41768 (.I(W18654), .ZN(W20675));
  INVX1 G41769 (.I(W27364), .ZN(W30060));
  INVX1 G41770 (.I(W17682), .ZN(W20676));
  INVX1 G41771 (.I(W16663), .ZN(O5189));
  INVX1 G41772 (.I(I1256), .ZN(W30100));
  INVX1 G41773 (.I(W21120), .ZN(W30098));
  INVX1 G41774 (.I(W8878), .ZN(W30097));
  INVX1 G41775 (.I(W17847), .ZN(W30096));
  INVX1 G41776 (.I(W9495), .ZN(W20685));
  INVX1 G41777 (.I(W14753), .ZN(W30093));
  INVX1 G41778 (.I(W22468), .ZN(W30091));
  INVX1 G41779 (.I(W3457), .ZN(W30009));
  INVX1 G41780 (.I(W6614), .ZN(W20741));
  INVX1 G41781 (.I(W15662), .ZN(W20748));
  INVX1 G41782 (.I(W7475), .ZN(W20751));
  INVX1 G41783 (.I(W12230), .ZN(W20752));
  INVX1 G41784 (.I(W19849), .ZN(W20753));
  INVX1 G41785 (.I(W21423), .ZN(W30017));
  INVX1 G41786 (.I(W19368), .ZN(W30014));
  INVX1 G41787 (.I(W1171), .ZN(W20756));
  INVX1 G41788 (.I(W19682), .ZN(W30011));
  INVX1 G41789 (.I(I682), .ZN(W30028));
  INVX1 G41790 (.I(W23356), .ZN(W30007));
  INVX1 G41791 (.I(I962), .ZN(W20763));
  INVX1 G41792 (.I(W22679), .ZN(W30004));
  INVX1 G41793 (.I(W25731), .ZN(O5149));
  INVX1 G41794 (.I(W13649), .ZN(W20770));
  INVX1 G41795 (.I(I1135), .ZN(O5147));
  INVX1 G41796 (.I(W28313), .ZN(W29997));
  INVX1 G41797 (.I(W27220), .ZN(W29996));
  INVX1 G41798 (.I(W14086), .ZN(W29995));
  INVX1 G41799 (.I(W2631), .ZN(W20724));
  INVX1 G41800 (.I(W6294), .ZN(W30058));
  INVX1 G41801 (.I(W11160), .ZN(O2064));
  INVX1 G41802 (.I(W2365), .ZN(W20717));
  INVX1 G41803 (.I(W21039), .ZN(W30055));
  INVX1 G41804 (.I(W408), .ZN(O5171));
  INVX1 G41805 (.I(W20655), .ZN(O5170));
  INVX1 G41806 (.I(W15543), .ZN(W20721));
  INVX1 G41807 (.I(I861), .ZN(O5169));
  INVX1 G41808 (.I(W8081), .ZN(W20723));
  INVX1 G41809 (.I(W6202), .ZN(W20882));
  INVX1 G41810 (.I(W21244), .ZN(W30045));
  INVX1 G41811 (.I(W18721), .ZN(O5166));
  INVX1 G41812 (.I(W3469), .ZN(W30042));
  INVX1 G41813 (.I(I432), .ZN(W30040));
  INVX1 G41814 (.I(W3243), .ZN(O5164));
  INVX1 G41815 (.I(W382), .ZN(W30036));
  INVX1 G41816 (.I(W29361), .ZN(O5162));
  INVX1 G41817 (.I(W10023), .ZN(W30032));
  INVX1 G41818 (.I(W29018), .ZN(W30029));
  INVX1 G41819 (.I(W29272), .ZN(W29709));
  INVX1 G41820 (.I(W3661), .ZN(W29724));
  INVX1 G41821 (.I(W19380), .ZN(W21036));
  INVX1 G41822 (.I(W9922), .ZN(W21037));
  INVX1 G41823 (.I(W19341), .ZN(W21038));
  INVX1 G41824 (.I(W18829), .ZN(W29717));
  INVX1 G41825 (.I(W8160), .ZN(W29716));
  INVX1 G41826 (.I(I1825), .ZN(W21044));
  INVX1 G41827 (.I(W248), .ZN(O5014));
  INVX1 G41828 (.I(W19782), .ZN(O5013));
  INVX1 G41829 (.I(W6529), .ZN(W21047));
  INVX1 G41830 (.I(W2735), .ZN(O5017));
  INVX1 G41831 (.I(W19040), .ZN(W21049));
  INVX1 G41832 (.I(W8187), .ZN(W21053));
  INVX1 G41833 (.I(W4053), .ZN(W29704));
  INVX1 G41834 (.I(W16558), .ZN(W29702));
  INVX1 G41835 (.I(W20128), .ZN(O5007));
  INVX1 G41836 (.I(I57), .ZN(W21061));
  INVX1 G41837 (.I(W4027), .ZN(W21065));
  INVX1 G41838 (.I(W13455), .ZN(W29693));
  INVX1 G41839 (.I(W6426), .ZN(W21066));
  INVX1 G41840 (.I(W14761), .ZN(O2136));
  INVX1 G41841 (.I(W26734), .ZN(W29757));
  INVX1 G41842 (.I(W15994), .ZN(O5028));
  INVX1 G41843 (.I(W15246), .ZN(W21008));
  INVX1 G41844 (.I(W10748), .ZN(W29753));
  INVX1 G41845 (.I(W11937), .ZN(W21009));
  INVX1 G41846 (.I(W18377), .ZN(W29751));
  INVX1 G41847 (.I(W9877), .ZN(W21010));
  INVX1 G41848 (.I(W6392), .ZN(W29748));
  INVX1 G41849 (.I(W15884), .ZN(W21014));
  INVX1 G41850 (.I(W17644), .ZN(O5005));
  INVX1 G41851 (.I(W24880), .ZN(W29744));
  INVX1 G41852 (.I(W18746), .ZN(W21016));
  INVX1 G41853 (.I(W20529), .ZN(W29742));
  INVX1 G41854 (.I(W9759), .ZN(W21019));
  INVX1 G41855 (.I(W19627), .ZN(O5019));
  INVX1 G41856 (.I(W18612), .ZN(W21025));
  INVX1 G41857 (.I(I559), .ZN(W29734));
  INVX1 G41858 (.I(W5418), .ZN(W21028));
  INVX1 G41859 (.I(W26298), .ZN(W29727));
  INVX1 G41860 (.I(W12088), .ZN(W21119));
  INVX1 G41861 (.I(W22087), .ZN(W29663));
  INVX1 G41862 (.I(W13126), .ZN(W21096));
  INVX1 G41863 (.I(W7294), .ZN(W21099));
  INVX1 G41864 (.I(W4385), .ZN(W21101));
  INVX1 G41865 (.I(W15858), .ZN(W29657));
  INVX1 G41866 (.I(I825), .ZN(W21108));
  INVX1 G41867 (.I(W10538), .ZN(O2153));
  INVX1 G41868 (.I(I1876), .ZN(W21113));
  INVX1 G41869 (.I(W5493), .ZN(O2154));
  INVX1 G41870 (.I(W1164), .ZN(W29665));
  INVX1 G41871 (.I(W7663), .ZN(O4987));
  INVX1 G41872 (.I(W16272), .ZN(W21124));
  INVX1 G41873 (.I(W10348), .ZN(W21125));
  INVX1 G41874 (.I(W14804), .ZN(W21126));
  INVX1 G41875 (.I(W13527), .ZN(O2155));
  INVX1 G41876 (.I(W11224), .ZN(O4984));
  INVX1 G41877 (.I(W19020), .ZN(W21128));
  INVX1 G41878 (.I(W26588), .ZN(W29636));
  INVX1 G41879 (.I(I700), .ZN(W29635));
  INVX1 G41880 (.I(W2591), .ZN(W29677));
  INVX1 G41881 (.I(W13316), .ZN(W21068));
  INVX1 G41882 (.I(W18652), .ZN(W21070));
  INVX1 G41883 (.I(W17988), .ZN(W21071));
  INVX1 G41884 (.I(W12262), .ZN(O2143));
  INVX1 G41885 (.I(W387), .ZN(O5001));
  INVX1 G41886 (.I(W12812), .ZN(W21074));
  INVX1 G41887 (.I(W14472), .ZN(O4999));
  INVX1 G41888 (.I(W6189), .ZN(W29679));
  INVX1 G41889 (.I(W16636), .ZN(W21081));
  INVX1 G41890 (.I(I1166), .ZN(W21004));
  INVX1 G41891 (.I(W7831), .ZN(W21082));
  INVX1 G41892 (.I(W9386), .ZN(W21085));
  INVX1 G41893 (.I(W11694), .ZN(O4997));
  INVX1 G41894 (.I(W9714), .ZN(O4996));
  INVX1 G41895 (.I(W7770), .ZN(W21090));
  INVX1 G41896 (.I(W26175), .ZN(W29669));
  INVX1 G41897 (.I(W19063), .ZN(W21091));
  INVX1 G41898 (.I(W6398), .ZN(W21092));
  INVX1 G41899 (.I(W39), .ZN(W21093));
  INVX1 G41900 (.I(W8423), .ZN(W20925));
  INVX1 G41901 (.I(W4842), .ZN(W20913));
  INVX1 G41902 (.I(W9099), .ZN(W20914));
  INVX1 G41903 (.I(W17897), .ZN(W20915));
  INVX1 G41904 (.I(W14589), .ZN(W29844));
  INVX1 G41905 (.I(W5065), .ZN(W29841));
  INVX1 G41906 (.I(W10388), .ZN(O5074));
  INVX1 G41907 (.I(W5043), .ZN(W20924));
  INVX1 G41908 (.I(W16975), .ZN(O5072));
  INVX1 G41909 (.I(W21153), .ZN(W29837));
  INVX1 G41910 (.I(W8314), .ZN(W29849));
  INVX1 G41911 (.I(W24113), .ZN(O5071));
  INVX1 G41912 (.I(W11759), .ZN(O5069));
  INVX1 G41913 (.I(W1163), .ZN(O2112));
  INVX1 G41914 (.I(W16402), .ZN(W29829));
  INVX1 G41915 (.I(W493), .ZN(W20932));
  INVX1 G41916 (.I(W8236), .ZN(O2113));
  INVX1 G41917 (.I(W13835), .ZN(W20935));
  INVX1 G41918 (.I(W21464), .ZN(W29820));
  INVX1 G41919 (.I(W9032), .ZN(O5061));
  INVX1 G41920 (.I(W8805), .ZN(W20902));
  INVX1 G41921 (.I(W18034), .ZN(W29882));
  INVX1 G41922 (.I(W14920), .ZN(W29880));
  INVX1 G41923 (.I(W11713), .ZN(O5091));
  INVX1 G41924 (.I(W25314), .ZN(O5089));
  INVX1 G41925 (.I(W17067), .ZN(W20894));
  INVX1 G41926 (.I(W18002), .ZN(W20897));
  INVX1 G41927 (.I(W1630), .ZN(W20898));
  INVX1 G41928 (.I(W18008), .ZN(W20899));
  INVX1 G41929 (.I(W13892), .ZN(W20901));
  INVX1 G41930 (.I(W18020), .ZN(O5060));
  INVX1 G41931 (.I(W29620), .ZN(W29861));
  INVX1 G41932 (.I(W15931), .ZN(W20903));
  INVX1 G41933 (.I(W19628), .ZN(W20904));
  INVX1 G41934 (.I(W24509), .ZN(W29857));
  INVX1 G41935 (.I(W13555), .ZN(W20909));
  INVX1 G41936 (.I(W25347), .ZN(O5079));
  INVX1 G41937 (.I(W18789), .ZN(W29852));
  INVX1 G41938 (.I(W14018), .ZN(W20912));
  INVX1 G41939 (.I(W5095), .ZN(W29850));
  INVX1 G41940 (.I(W8142), .ZN(W20991));
  INVX1 G41941 (.I(W9569), .ZN(W29782));
  INVX1 G41942 (.I(I339), .ZN(W29781));
  INVX1 G41943 (.I(W13770), .ZN(W20986));
  INVX1 G41944 (.I(I607), .ZN(O2130));
  INVX1 G41945 (.I(W1262), .ZN(W20988));
  INVX1 G41946 (.I(W15489), .ZN(W20989));
  INVX1 G41947 (.I(W20241), .ZN(W20990));
  INVX1 G41948 (.I(I1178), .ZN(O5037));
  INVX1 G41949 (.I(W28329), .ZN(W29773));
  INVX1 G41950 (.I(W17740), .ZN(O2127));
  INVX1 G41951 (.I(W6595), .ZN(W20992));
  INVX1 G41952 (.I(W20542), .ZN(O2131));
  INVX1 G41953 (.I(W9240), .ZN(O5035));
  INVX1 G41954 (.I(W12065), .ZN(O5033));
  INVX1 G41955 (.I(W2091), .ZN(O5032));
  INVX1 G41956 (.I(I1649), .ZN(W20997));
  INVX1 G41957 (.I(W14473), .ZN(W20999));
  INVX1 G41958 (.I(W7046), .ZN(W21000));
  INVX1 G41959 (.I(W11467), .ZN(W21003));
  INVX1 G41960 (.I(W7578), .ZN(W20959));
  INVX1 G41961 (.I(W21954), .ZN(O5059));
  INVX1 G41962 (.I(W21898), .ZN(W29814));
  INVX1 G41963 (.I(I721), .ZN(W20946));
  INVX1 G41964 (.I(W27184), .ZN(O5055));
  INVX1 G41965 (.I(W247), .ZN(O5054));
  INVX1 G41966 (.I(W17129), .ZN(O2118));
  INVX1 G41967 (.I(W1303), .ZN(W29806));
  INVX1 G41968 (.I(W560), .ZN(W29805));
  INVX1 G41969 (.I(W6852), .ZN(O5053));
  INVX1 G41970 (.I(W16474), .ZN(W19781));
  INVX1 G41971 (.I(W1039), .ZN(W20960));
  INVX1 G41972 (.I(W7674), .ZN(O5050));
  INVX1 G41973 (.I(W18951), .ZN(W20967));
  INVX1 G41974 (.I(W7933), .ZN(W20969));
  INVX1 G41975 (.I(W1256), .ZN(O5045));
  INVX1 G41976 (.I(W12060), .ZN(W20973));
  INVX1 G41977 (.I(W706), .ZN(W20975));
  INVX1 G41978 (.I(W2142), .ZN(O2126));
  INVX1 G41979 (.I(W15144), .ZN(W29785));
  INVX1 G41980 (.I(W8418), .ZN(W18492));
  INVX1 G41981 (.I(I193), .ZN(W18477));
  INVX1 G41982 (.I(W27582), .ZN(W32353));
  INVX1 G41983 (.I(I100), .ZN(W18479));
  INVX1 G41984 (.I(I587), .ZN(W18480));
  INVX1 G41985 (.I(W21037), .ZN(W32349));
  INVX1 G41986 (.I(W13256), .ZN(O6202));
  INVX1 G41987 (.I(W11828), .ZN(W18485));
  INVX1 G41988 (.I(W15526), .ZN(W18487));
  INVX1 G41989 (.I(W11632), .ZN(W18488));
  INVX1 G41990 (.I(W3317), .ZN(W18491));
  INVX1 G41991 (.I(W4273), .ZN(W32355));
  INVX1 G41992 (.I(W16512), .ZN(O6198));
  INVX1 G41993 (.I(W4099), .ZN(W18495));
  INVX1 G41994 (.I(W11220), .ZN(W18497));
  INVX1 G41995 (.I(W2740), .ZN(W18501));
  INVX1 G41996 (.I(W1372), .ZN(W32328));
  INVX1 G41997 (.I(W95), .ZN(O6192));
  INVX1 G41998 (.I(W23800), .ZN(O6191));
  INVX1 G41999 (.I(W5574), .ZN(W18503));
  INVX1 G42000 (.I(W4386), .ZN(W32323));
  INVX1 G42001 (.I(W1058), .ZN(W18471));
  INVX1 G42002 (.I(W2489), .ZN(W18465));
  INVX1 G42003 (.I(W24323), .ZN(O6213));
  INVX1 G42004 (.I(W5570), .ZN(W18467));
  INVX1 G42005 (.I(I639), .ZN(W18468));
  INVX1 G42006 (.I(W22841), .ZN(W32373));
  INVX1 G42007 (.I(W11369), .ZN(W32372));
  INVX1 G42008 (.I(W18516), .ZN(W32371));
  INVX1 G42009 (.I(W28986), .ZN(W32370));
  INVX1 G42010 (.I(W3843), .ZN(W32368));
  INVX1 G42011 (.I(W6809), .ZN(O1575));
  INVX1 G42012 (.I(W17845), .ZN(W18473));
  INVX1 G42013 (.I(W13662), .ZN(W32365));
  INVX1 G42014 (.I(W13869), .ZN(O6211));
  INVX1 G42015 (.I(W1727), .ZN(W18476));
  INVX1 G42016 (.I(W18846), .ZN(O6209));
  INVX1 G42017 (.I(W11695), .ZN(W32359));
  INVX1 G42018 (.I(W28887), .ZN(O6208));
  INVX1 G42019 (.I(W4835), .ZN(O6207));
  INVX1 G42020 (.I(W9965), .ZN(O6206));
  INVX1 G42021 (.I(W16119), .ZN(O1588));
  INVX1 G42022 (.I(W15226), .ZN(W18549));
  INVX1 G42023 (.I(W8989), .ZN(W32283));
  INVX1 G42024 (.I(W1763), .ZN(O1585));
  INVX1 G42025 (.I(W16503), .ZN(W32281));
  INVX1 G42026 (.I(W3265), .ZN(W32280));
  INVX1 G42027 (.I(W7270), .ZN(W32277));
  INVX1 G42028 (.I(W25833), .ZN(W32275));
  INVX1 G42029 (.I(W3210), .ZN(O6171));
  INVX1 G42030 (.I(W2761), .ZN(O6170));
  INVX1 G42031 (.I(W5596), .ZN(W18545));
  INVX1 G42032 (.I(W10617), .ZN(W18564));
  INVX1 G42033 (.I(W1895), .ZN(W18567));
  INVX1 G42034 (.I(W30271), .ZN(W32266));
  INVX1 G42035 (.I(W10683), .ZN(W18570));
  INVX1 G42036 (.I(W11000), .ZN(O1589));
  INVX1 G42037 (.I(W9355), .ZN(W32262));
  INVX1 G42038 (.I(W13457), .ZN(O6166));
  INVX1 G42039 (.I(W13829), .ZN(W18573));
  INVX1 G42040 (.I(W8379), .ZN(W18575));
  INVX1 G42041 (.I(W17690), .ZN(O1579));
  INVX1 G42042 (.I(I1604), .ZN(W18507));
  INVX1 G42043 (.I(W15161), .ZN(W32319));
  INVX1 G42044 (.I(W26680), .ZN(O6188));
  INVX1 G42045 (.I(W10982), .ZN(W18513));
  INVX1 G42046 (.I(W3262), .ZN(W18517));
  INVX1 G42047 (.I(W6079), .ZN(W18518));
  INVX1 G42048 (.I(W14140), .ZN(W18519));
  INVX1 G42049 (.I(W11933), .ZN(W18522));
  INVX1 G42050 (.I(W6782), .ZN(O6183));
  INVX1 G42051 (.I(W733), .ZN(W18464));
  INVX1 G42052 (.I(W13688), .ZN(O1580));
  INVX1 G42053 (.I(W29203), .ZN(W32304));
  INVX1 G42054 (.I(W2646), .ZN(O6182));
  INVX1 G42055 (.I(W26328), .ZN(O6180));
  INVX1 G42056 (.I(W31140), .ZN(O6178));
  INVX1 G42057 (.I(W7328), .ZN(W18533));
  INVX1 G42058 (.I(W23885), .ZN(W32294));
  INVX1 G42059 (.I(W9618), .ZN(W18543));
  INVX1 G42060 (.I(W1826), .ZN(W18544));
  INVX1 G42061 (.I(W950), .ZN(W18404));
  INVX1 G42062 (.I(W927), .ZN(W18391));
  INVX1 G42063 (.I(W29628), .ZN(W32462));
  INVX1 G42064 (.I(W559), .ZN(W18392));
  INVX1 G42065 (.I(W31018), .ZN(W32460));
  INVX1 G42066 (.I(W13578), .ZN(W18393));
  INVX1 G42067 (.I(W2885), .ZN(W32457));
  INVX1 G42068 (.I(W7086), .ZN(W18397));
  INVX1 G42069 (.I(W16634), .ZN(W18399));
  INVX1 G42070 (.I(W31560), .ZN(W32452));
  INVX1 G42071 (.I(W8708), .ZN(W32451));
  INVX1 G42072 (.I(W16477), .ZN(W18390));
  INVX1 G42073 (.I(W16040), .ZN(O6242));
  INVX1 G42074 (.I(W15915), .ZN(O1560));
  INVX1 G42075 (.I(W10306), .ZN(O1561));
  INVX1 G42076 (.I(W10322), .ZN(O1562));
  INVX1 G42077 (.I(W12955), .ZN(W18412));
  INVX1 G42078 (.I(W21800), .ZN(W32442));
  INVX1 G42079 (.I(W1527), .ZN(W18413));
  INVX1 G42080 (.I(W23887), .ZN(W32439));
  INVX1 G42081 (.I(W29517), .ZN(O6238));
  INVX1 G42082 (.I(W6639), .ZN(W18372));
  INVX1 G42083 (.I(W16395), .ZN(O1556));
  INVX1 G42084 (.I(W12880), .ZN(W18366));
  INVX1 G42085 (.I(W12033), .ZN(W32487));
  INVX1 G42086 (.I(W32027), .ZN(O6252));
  INVX1 G42087 (.I(W6493), .ZN(W32485));
  INVX1 G42088 (.I(I447), .ZN(W18367));
  INVX1 G42089 (.I(W1527), .ZN(W18369));
  INVX1 G42090 (.I(W3519), .ZN(O1558));
  INVX1 G42091 (.I(I921), .ZN(W18371));
  INVX1 G42092 (.I(W23982), .ZN(W32437));
  INVX1 G42093 (.I(W8504), .ZN(W18376));
  INVX1 G42094 (.I(W244), .ZN(W18377));
  INVX1 G42095 (.I(W19430), .ZN(W32477));
  INVX1 G42096 (.I(W1709), .ZN(W32476));
  INVX1 G42097 (.I(W8234), .ZN(O6248));
  INVX1 G42098 (.I(W3574), .ZN(W18379));
  INVX1 G42099 (.I(W32365), .ZN(W32472));
  INVX1 G42100 (.I(W7736), .ZN(W18383));
  INVX1 G42101 (.I(W11488), .ZN(W32468));
  INVX1 G42102 (.I(W29738), .ZN(W32392));
  INVX1 G42103 (.I(W232), .ZN(W32405));
  INVX1 G42104 (.I(W5793), .ZN(W32404));
  INVX1 G42105 (.I(W11823), .ZN(W32403));
  INVX1 G42106 (.I(W10951), .ZN(W18445));
  INVX1 G42107 (.I(W21642), .ZN(O6224));
  INVX1 G42108 (.I(W18214), .ZN(W18449));
  INVX1 G42109 (.I(W17803), .ZN(W18452));
  INVX1 G42110 (.I(W9653), .ZN(O6222));
  INVX1 G42111 (.I(I142), .ZN(O6221));
  INVX1 G42112 (.I(W20100), .ZN(W32406));
  INVX1 G42113 (.I(W11800), .ZN(O6220));
  INVX1 G42114 (.I(W10012), .ZN(W18455));
  INVX1 G42115 (.I(W5003), .ZN(W18456));
  INVX1 G42116 (.I(W25510), .ZN(W32388));
  INVX1 G42117 (.I(W17232), .ZN(W32387));
  INVX1 G42118 (.I(W19522), .ZN(O6218));
  INVX1 G42119 (.I(W9352), .ZN(W18460));
  INVX1 G42120 (.I(W25011), .ZN(O6216));
  INVX1 G42121 (.I(W1273), .ZN(W18462));
  INVX1 G42122 (.I(W3879), .ZN(O6233));
  INVX1 G42123 (.I(W10589), .ZN(W18415));
  INVX1 G42124 (.I(W4726), .ZN(O6237));
  INVX1 G42125 (.I(W210), .ZN(W18416));
  INVX1 G42126 (.I(W28038), .ZN(O6236));
  INVX1 G42127 (.I(W8634), .ZN(W18417));
  INVX1 G42128 (.I(W14217), .ZN(O6234));
  INVX1 G42129 (.I(W3699), .ZN(O1563));
  INVX1 G42130 (.I(W12983), .ZN(W18419));
  INVX1 G42131 (.I(W2017), .ZN(W18420));
  INVX1 G42132 (.I(W7692), .ZN(W18576));
  INVX1 G42133 (.I(I540), .ZN(W18426));
  INVX1 G42134 (.I(W16619), .ZN(W18429));
  INVX1 G42135 (.I(W8595), .ZN(W18430));
  INVX1 G42136 (.I(W22994), .ZN(W32420));
  INVX1 G42137 (.I(W17128), .ZN(O6229));
  INVX1 G42138 (.I(W15564), .ZN(W18439));
  INVX1 G42139 (.I(W20610), .ZN(W32411));
  INVX1 G42140 (.I(W13878), .ZN(W32408));
  INVX1 G42141 (.I(W25462), .ZN(W32407));
  INVX1 G42142 (.I(W17013), .ZN(O1642));
  INVX1 G42143 (.I(W11957), .ZN(W18746));
  INVX1 G42144 (.I(W13754), .ZN(W32093));
  INVX1 G42145 (.I(W5950), .ZN(O6088));
  INVX1 G42146 (.I(W11959), .ZN(W18754));
  INVX1 G42147 (.I(W27476), .ZN(O6086));
  INVX1 G42148 (.I(W26745), .ZN(W32086));
  INVX1 G42149 (.I(W7304), .ZN(O1640));
  INVX1 G42150 (.I(W4694), .ZN(O1641));
  INVX1 G42151 (.I(W4636), .ZN(O6082));
  INVX1 G42152 (.I(W9783), .ZN(W18769));
  INVX1 G42153 (.I(W1648), .ZN(W32099));
  INVX1 G42154 (.I(W15075), .ZN(W18772));
  INVX1 G42155 (.I(I1273), .ZN(O1644));
  INVX1 G42156 (.I(W11098), .ZN(W18775));
  INVX1 G42157 (.I(W10481), .ZN(W18776));
  INVX1 G42158 (.I(W20020), .ZN(O6078));
  INVX1 G42159 (.I(W16589), .ZN(O1645));
  INVX1 G42160 (.I(W31247), .ZN(W32065));
  INVX1 G42161 (.I(W3246), .ZN(O1648));
  INVX1 G42162 (.I(W21195), .ZN(O6074));
  INVX1 G42163 (.I(W1087), .ZN(O6097));
  INVX1 G42164 (.I(W6847), .ZN(W18708));
  INVX1 G42165 (.I(W1019), .ZN(W18710));
  INVX1 G42166 (.I(W14865), .ZN(O6102));
  INVX1 G42167 (.I(W14543), .ZN(W18711));
  INVX1 G42168 (.I(W11991), .ZN(O6100));
  INVX1 G42169 (.I(W8290), .ZN(W18712));
  INVX1 G42170 (.I(W11489), .ZN(O1627));
  INVX1 G42171 (.I(W8259), .ZN(O1628));
  INVX1 G42172 (.I(W21589), .ZN(W32119));
  INVX1 G42173 (.I(W24696), .ZN(W32061));
  INVX1 G42174 (.I(W1782), .ZN(W18727));
  INVX1 G42175 (.I(W14509), .ZN(W18731));
  INVX1 G42176 (.I(W6302), .ZN(W18737));
  INVX1 G42177 (.I(W21492), .ZN(O6094));
  INVX1 G42178 (.I(I284), .ZN(W18740));
  INVX1 G42179 (.I(W23286), .ZN(O6092));
  INVX1 G42180 (.I(W3364), .ZN(O1633));
  INVX1 G42181 (.I(W20274), .ZN(W32103));
  INVX1 G42182 (.I(W7200), .ZN(W32100));
  INVX1 G42183 (.I(W2461), .ZN(W18832));
  INVX1 G42184 (.I(W1301), .ZN(O1653));
  INVX1 G42185 (.I(W31619), .ZN(O6062));
  INVX1 G42186 (.I(W3383), .ZN(O1654));
  INVX1 G42187 (.I(W12121), .ZN(W32027));
  INVX1 G42188 (.I(W3946), .ZN(W32026));
  INVX1 G42189 (.I(W867), .ZN(W18830));
  INVX1 G42190 (.I(I742), .ZN(W32022));
  INVX1 G42191 (.I(I1092), .ZN(O6057));
  INVX1 G42192 (.I(W10162), .ZN(O6056));
  INVX1 G42193 (.I(W4048), .ZN(W18821));
  INVX1 G42194 (.I(W7479), .ZN(W32017));
  INVX1 G42195 (.I(W9538), .ZN(W18834));
  INVX1 G42196 (.I(W8303), .ZN(O1658));
  INVX1 G42197 (.I(W13313), .ZN(O1660));
  INVX1 G42198 (.I(W23508), .ZN(O6051));
  INVX1 G42199 (.I(W11774), .ZN(W18841));
  INVX1 G42200 (.I(W22362), .ZN(O6049));
  INVX1 G42201 (.I(W17531), .ZN(W32007));
  INVX1 G42202 (.I(W16043), .ZN(W32006));
  INVX1 G42203 (.I(W10596), .ZN(W18802));
  INVX1 G42204 (.I(W30221), .ZN(W32060));
  INVX1 G42205 (.I(W17268), .ZN(O1649));
  INVX1 G42206 (.I(I758), .ZN(W32057));
  INVX1 G42207 (.I(W25936), .ZN(W32056));
  INVX1 G42208 (.I(W7580), .ZN(O6071));
  INVX1 G42209 (.I(W5817), .ZN(W18798));
  INVX1 G42210 (.I(W12705), .ZN(W18800));
  INVX1 G42211 (.I(W19053), .ZN(W32049));
  INVX1 G42212 (.I(W19287), .ZN(W32048));
  INVX1 G42213 (.I(W5622), .ZN(O1626));
  INVX1 G42214 (.I(W21220), .ZN(W32046));
  INVX1 G42215 (.I(W22007), .ZN(W32042));
  INVX1 G42216 (.I(W16962), .ZN(O1651));
  INVX1 G42217 (.I(W12997), .ZN(W18814));
  INVX1 G42218 (.I(W11931), .ZN(W18815));
  INVX1 G42219 (.I(W6697), .ZN(W18817));
  INVX1 G42220 (.I(W238), .ZN(W18819));
  INVX1 G42221 (.I(W12328), .ZN(W32035));
  INVX1 G42222 (.I(W12092), .ZN(W18820));
  INVX1 G42223 (.I(W5125), .ZN(W18627));
  INVX1 G42224 (.I(W9850), .ZN(W18616));
  INVX1 G42225 (.I(W4975), .ZN(O6150));
  INVX1 G42226 (.I(W8959), .ZN(O6149));
  INVX1 G42227 (.I(W1165), .ZN(W32221));
  INVX1 G42228 (.I(I1726), .ZN(W32220));
  INVX1 G42229 (.I(I1708), .ZN(W18621));
  INVX1 G42230 (.I(W8137), .ZN(W32217));
  INVX1 G42231 (.I(W16939), .ZN(W18623));
  INVX1 G42232 (.I(W1518), .ZN(W18624));
  INVX1 G42233 (.I(W2265), .ZN(O1602));
  INVX1 G42234 (.I(W15592), .ZN(O1607));
  INVX1 G42235 (.I(W28262), .ZN(W32212));
  INVX1 G42236 (.I(W9342), .ZN(W18631));
  INVX1 G42237 (.I(W21627), .ZN(W32209));
  INVX1 G42238 (.I(I1396), .ZN(W32208));
  INVX1 G42239 (.I(W6517), .ZN(O6146));
  INVX1 G42240 (.I(I270), .ZN(W18632));
  INVX1 G42241 (.I(W1157), .ZN(W18634));
  INVX1 G42242 (.I(W31510), .ZN(W32203));
  INVX1 G42243 (.I(W8629), .ZN(W18595));
  INVX1 G42244 (.I(W15133), .ZN(W32256));
  INVX1 G42245 (.I(W17610), .ZN(W18578));
  INVX1 G42246 (.I(I347), .ZN(W18581));
  INVX1 G42247 (.I(W17755), .ZN(O1594));
  INVX1 G42248 (.I(I827), .ZN(W32249));
  INVX1 G42249 (.I(W3431), .ZN(O1596));
  INVX1 G42250 (.I(W22079), .ZN(W32247));
  INVX1 G42251 (.I(W4198), .ZN(O6161));
  INVX1 G42252 (.I(I1400), .ZN(W18593));
  INVX1 G42253 (.I(I1270), .ZN(W18635));
  INVX1 G42254 (.I(I303), .ZN(O1598));
  INVX1 G42255 (.I(W19851), .ZN(O6156));
  INVX1 G42256 (.I(W3629), .ZN(W18600));
  INVX1 G42257 (.I(W14332), .ZN(W32237));
  INVX1 G42258 (.I(W15309), .ZN(O1599));
  INVX1 G42259 (.I(W14468), .ZN(O6155));
  INVX1 G42260 (.I(W16613), .ZN(O1600));
  INVX1 G42261 (.I(W16201), .ZN(W18607));
  INVX1 G42262 (.I(W2671), .ZN(W18608));
  INVX1 G42263 (.I(W4989), .ZN(W18691));
  INVX1 G42264 (.I(W14986), .ZN(W32166));
  INVX1 G42265 (.I(W12109), .ZN(W18672));
  INVX1 G42266 (.I(W3780), .ZN(O6121));
  INVX1 G42267 (.I(W7598), .ZN(W32155));
  INVX1 G42268 (.I(W8384), .ZN(O6119));
  INVX1 G42269 (.I(I602), .ZN(W32153));
  INVX1 G42270 (.I(W21375), .ZN(O6118));
  INVX1 G42271 (.I(W17852), .ZN(W18689));
  INVX1 G42272 (.I(W4060), .ZN(W32149));
  INVX1 G42273 (.I(W22259), .ZN(O6126));
  INVX1 G42274 (.I(W18990), .ZN(O6115));
  INVX1 G42275 (.I(W17099), .ZN(W18695));
  INVX1 G42276 (.I(W12365), .ZN(W18697));
  INVX1 G42277 (.I(W283), .ZN(W18699));
  INVX1 G42278 (.I(W26438), .ZN(W32138));
  INVX1 G42279 (.I(W24306), .ZN(W32136));
  INVX1 G42280 (.I(W20705), .ZN(W32135));
  INVX1 G42281 (.I(W14462), .ZN(W18704));
  INVX1 G42282 (.I(W12538), .ZN(O1625));
  INVX1 G42283 (.I(W11763), .ZN(O1616));
  INVX1 G42284 (.I(W17264), .ZN(W18637));
  INVX1 G42285 (.I(W4386), .ZN(W18639));
  INVX1 G42286 (.I(W16434), .ZN(O6140));
  INVX1 G42287 (.I(W6282), .ZN(W18644));
  INVX1 G42288 (.I(W18187), .ZN(O1612));
  INVX1 G42289 (.I(W1853), .ZN(O6136));
  INVX1 G42290 (.I(W3172), .ZN(W32189));
  INVX1 G42291 (.I(W5752), .ZN(W18649));
  INVX1 G42292 (.I(W11989), .ZN(W32185));
  INVX1 G42293 (.I(I1509), .ZN(W32491));
  INVX1 G42294 (.I(W1201), .ZN(W18656));
  INVX1 G42295 (.I(W6234), .ZN(W18657));
  INVX1 G42296 (.I(W8357), .ZN(W18658));
  INVX1 G42297 (.I(W19487), .ZN(O6132));
  INVX1 G42298 (.I(W13050), .ZN(W32174));
  INVX1 G42299 (.I(W140), .ZN(O6129));
  INVX1 G42300 (.I(W15891), .ZN(W32171));
  INVX1 G42301 (.I(W128), .ZN(W32169));
  INVX1 G42302 (.I(W2791), .ZN(W18671));
  INVX1 G42303 (.I(W11784), .ZN(O6397));
  INVX1 G42304 (.I(W8395), .ZN(W18061));
  INVX1 G42305 (.I(W14056), .ZN(O6406));
  INVX1 G42306 (.I(W11680), .ZN(W18063));
  INVX1 G42307 (.I(W18624), .ZN(W32804));
  INVX1 G42308 (.I(I1610), .ZN(W18064));
  INVX1 G42309 (.I(W18890), .ZN(O6403));
  INVX1 G42310 (.I(W10623), .ZN(W18067));
  INVX1 G42311 (.I(W20258), .ZN(O6401));
  INVX1 G42312 (.I(W25082), .ZN(W32796));
  INVX1 G42313 (.I(W21766), .ZN(W32795));
  INVX1 G42314 (.I(W9838), .ZN(W32809));
  INVX1 G42315 (.I(I1808), .ZN(W18075));
  INVX1 G42316 (.I(W3842), .ZN(W18076));
  INVX1 G42317 (.I(W13199), .ZN(W18077));
  INVX1 G42318 (.I(W16146), .ZN(O6395));
  INVX1 G42319 (.I(W9583), .ZN(O6393));
  INVX1 G42320 (.I(W16372), .ZN(W18081));
  INVX1 G42321 (.I(W9615), .ZN(W18083));
  INVX1 G42322 (.I(W11818), .ZN(W18086));
  INVX1 G42323 (.I(W6786), .ZN(W32776));
  INVX1 G42324 (.I(W17097), .ZN(W32823));
  INVX1 G42325 (.I(W6928), .ZN(W18029));
  INVX1 G42326 (.I(W8117), .ZN(W18034));
  INVX1 G42327 (.I(W13439), .ZN(W18035));
  INVX1 G42328 (.I(W2072), .ZN(W18037));
  INVX1 G42329 (.I(I1134), .ZN(W32832));
  INVX1 G42330 (.I(W24192), .ZN(O6417));
  INVX1 G42331 (.I(W13005), .ZN(O6416));
  INVX1 G42332 (.I(W15243), .ZN(W32826));
  INVX1 G42333 (.I(W19101), .ZN(O6415));
  INVX1 G42334 (.I(W14331), .ZN(O1501));
  INVX1 G42335 (.I(W1731), .ZN(O6414));
  INVX1 G42336 (.I(W130), .ZN(O6413));
  INVX1 G42337 (.I(W25839), .ZN(O6412));
  INVX1 G42338 (.I(W13555), .ZN(W18050));
  INVX1 G42339 (.I(W18725), .ZN(O6410));
  INVX1 G42340 (.I(I253), .ZN(O1490));
  INVX1 G42341 (.I(W30736), .ZN(O6409));
  INVX1 G42342 (.I(I220), .ZN(W18053));
  INVX1 G42343 (.I(W2456), .ZN(W32811));
  INVX1 G42344 (.I(I1370), .ZN(O6375));
  INVX1 G42345 (.I(W13445), .ZN(W32748));
  INVX1 G42346 (.I(W5229), .ZN(O6380));
  INVX1 G42347 (.I(W2215), .ZN(W18115));
  INVX1 G42348 (.I(W6301), .ZN(W32743));
  INVX1 G42349 (.I(W27811), .ZN(O6378));
  INVX1 G42350 (.I(W22524), .ZN(O6377));
  INVX1 G42351 (.I(W25454), .ZN(W32740));
  INVX1 G42352 (.I(W18447), .ZN(O6376));
  INVX1 G42353 (.I(W9175), .ZN(W32738));
  INVX1 G42354 (.I(W14338), .ZN(W32749));
  INVX1 G42355 (.I(W23746), .ZN(O6374));
  INVX1 G42356 (.I(W21999), .ZN(W32734));
  INVX1 G42357 (.I(W9682), .ZN(W18118));
  INVX1 G42358 (.I(W6327), .ZN(O1506));
  INVX1 G42359 (.I(W5765), .ZN(O6371));
  INVX1 G42360 (.I(W3315), .ZN(W18121));
  INVX1 G42361 (.I(W1477), .ZN(W18122));
  INVX1 G42362 (.I(W12507), .ZN(W18125));
  INVX1 G42363 (.I(W17995), .ZN(W18127));
  INVX1 G42364 (.I(W14205), .ZN(W32762));
  INVX1 G42365 (.I(W5680), .ZN(W18093));
  INVX1 G42366 (.I(W8607), .ZN(W18094));
  INVX1 G42367 (.I(W31642), .ZN(W32771));
  INVX1 G42368 (.I(W8323), .ZN(W18095));
  INVX1 G42369 (.I(W3736), .ZN(W18096));
  INVX1 G42370 (.I(W7538), .ZN(W18100));
  INVX1 G42371 (.I(W17617), .ZN(W32765));
  INVX1 G42372 (.I(W31411), .ZN(W32764));
  INVX1 G42373 (.I(W18063), .ZN(W18104));
  INVX1 G42374 (.I(W13085), .ZN(W18028));
  INVX1 G42375 (.I(W17848), .ZN(O6387));
  INVX1 G42376 (.I(W222), .ZN(W18106));
  INVX1 G42377 (.I(W14658), .ZN(O6385));
  INVX1 G42378 (.I(W5727), .ZN(O1502));
  INVX1 G42379 (.I(W15693), .ZN(W32756));
  INVX1 G42380 (.I(W1934), .ZN(W32755));
  INVX1 G42381 (.I(W2384), .ZN(W18108));
  INVX1 G42382 (.I(W12889), .ZN(O6382));
  INVX1 G42383 (.I(W1320), .ZN(W32750));
  INVX1 G42384 (.I(W30170), .ZN(W32920));
  INVX1 G42385 (.I(W8706), .ZN(O1470));
  INVX1 G42386 (.I(W18414), .ZN(O6459));
  INVX1 G42387 (.I(W12772), .ZN(W32928));
  INVX1 G42388 (.I(W8748), .ZN(W17934));
  INVX1 G42389 (.I(W297), .ZN(W17935));
  INVX1 G42390 (.I(W30069), .ZN(W32925));
  INVX1 G42391 (.I(W15728), .ZN(W17938));
  INVX1 G42392 (.I(W14453), .ZN(W17939));
  INVX1 G42393 (.I(I722), .ZN(W32921));
  INVX1 G42394 (.I(W3616), .ZN(W17931));
  INVX1 G42395 (.I(W5444), .ZN(W32919));
  INVX1 G42396 (.I(W31151), .ZN(O6456));
  INVX1 G42397 (.I(W19461), .ZN(O6455));
  INVX1 G42398 (.I(W3035), .ZN(O6454));
  INVX1 G42399 (.I(I495), .ZN(O1473));
  INVX1 G42400 (.I(W533), .ZN(W32914));
  INVX1 G42401 (.I(W27269), .ZN(W32913));
  INVX1 G42402 (.I(W30358), .ZN(W32912));
  INVX1 G42403 (.I(W17712), .ZN(W17946));
  INVX1 G42404 (.I(W22772), .ZN(W32946));
  INVX1 G42405 (.I(W327), .ZN(O1467));
  INVX1 G42406 (.I(W2583), .ZN(W32957));
  INVX1 G42407 (.I(W24429), .ZN(O6472));
  INVX1 G42408 (.I(W8755), .ZN(W17914));
  INVX1 G42409 (.I(W280), .ZN(O6470));
  INVX1 G42410 (.I(W23798), .ZN(W32951));
  INVX1 G42411 (.I(W12015), .ZN(O6468));
  INVX1 G42412 (.I(W15337), .ZN(W17917));
  INVX1 G42413 (.I(W6574), .ZN(W17919));
  INVX1 G42414 (.I(W7201), .ZN(W17949));
  INVX1 G42415 (.I(W10894), .ZN(W32945));
  INVX1 G42416 (.I(W17136), .ZN(W17920));
  INVX1 G42417 (.I(W13429), .ZN(O6466));
  INVX1 G42418 (.I(W6553), .ZN(W17923));
  INVX1 G42419 (.I(W17645), .ZN(W17926));
  INVX1 G42420 (.I(W32367), .ZN(W32936));
  INVX1 G42421 (.I(W5988), .ZN(O6462));
  INVX1 G42422 (.I(W5208), .ZN(W32934));
  INVX1 G42423 (.I(W3864), .ZN(W17930));
  INVX1 G42424 (.I(W8883), .ZN(O6433));
  INVX1 G42425 (.I(W1300), .ZN(O6442));
  INVX1 G42426 (.I(W16228), .ZN(W17996));
  INVX1 G42427 (.I(I1036), .ZN(W32871));
  INVX1 G42428 (.I(W16046), .ZN(W32870));
  INVX1 G42429 (.I(W15960), .ZN(W18002));
  INVX1 G42430 (.I(W13645), .ZN(W18008));
  INVX1 G42431 (.I(W16482), .ZN(O1483));
  INVX1 G42432 (.I(W8166), .ZN(O1486));
  INVX1 G42433 (.I(W30425), .ZN(O6434));
  INVX1 G42434 (.I(W12819), .ZN(W17992));
  INVX1 G42435 (.I(W4303), .ZN(O6432));
  INVX1 G42436 (.I(I163), .ZN(W18021));
  INVX1 G42437 (.I(W25571), .ZN(W32850));
  INVX1 G42438 (.I(I560), .ZN(W18022));
  INVX1 G42439 (.I(W312), .ZN(W18025));
  INVX1 G42440 (.I(I351), .ZN(O6427));
  INVX1 G42441 (.I(W31765), .ZN(W32845));
  INVX1 G42442 (.I(W7883), .ZN(W32844));
  INVX1 G42443 (.I(W14963), .ZN(W32843));
  INVX1 G42444 (.I(W14521), .ZN(O6448));
  INVX1 G42445 (.I(W13073), .ZN(W17952));
  INVX1 G42446 (.I(W24916), .ZN(W32906));
  INVX1 G42447 (.I(W8876), .ZN(W17954));
  INVX1 G42448 (.I(W13324), .ZN(W32900));
  INVX1 G42449 (.I(W8038), .ZN(W17965));
  INVX1 G42450 (.I(W20827), .ZN(W32895));
  INVX1 G42451 (.I(W3398), .ZN(W17971));
  INVX1 G42452 (.I(W2466), .ZN(O1478));
  INVX1 G42453 (.I(W4431), .ZN(W17973));
  INVX1 G42454 (.I(W543), .ZN(O1508));
  INVX1 G42455 (.I(I1362), .ZN(W17974));
  INVX1 G42456 (.I(W5259), .ZN(W17980));
  INVX1 G42457 (.I(W16321), .ZN(W32887));
  INVX1 G42458 (.I(W5519), .ZN(W17984));
  INVX1 G42459 (.I(W5782), .ZN(W17985));
  INVX1 G42460 (.I(W14171), .ZN(W17986));
  INVX1 G42461 (.I(W20180), .ZN(W32882));
  INVX1 G42462 (.I(W4643), .ZN(W32881));
  INVX1 G42463 (.I(W17970), .ZN(O1479));
  INVX1 G42464 (.I(W25706), .ZN(W32576));
  INVX1 G42465 (.I(W11544), .ZN(O6302));
  INVX1 G42466 (.I(W12620), .ZN(W32589));
  INVX1 G42467 (.I(W22529), .ZN(O6301));
  INVX1 G42468 (.I(W9854), .ZN(O6300));
  INVX1 G42469 (.I(W9685), .ZN(O6299));
  INVX1 G42470 (.I(W25246), .ZN(O6298));
  INVX1 G42471 (.I(W5351), .ZN(O1534));
  INVX1 G42472 (.I(W26419), .ZN(O6297));
  INVX1 G42473 (.I(W338), .ZN(O1535));
  INVX1 G42474 (.I(W31263), .ZN(W32577));
  INVX1 G42475 (.I(W1538), .ZN(O1532));
  INVX1 G42476 (.I(W13537), .ZN(W18278));
  INVX1 G42477 (.I(W3648), .ZN(O1538));
  INVX1 G42478 (.I(W15391), .ZN(W18289));
  INVX1 G42479 (.I(W8528), .ZN(O1539));
  INVX1 G42480 (.I(W6941), .ZN(O6291));
  INVX1 G42481 (.I(W9145), .ZN(W18291));
  INVX1 G42482 (.I(W24784), .ZN(O6290));
  INVX1 G42483 (.I(W14155), .ZN(O1540));
  INVX1 G42484 (.I(W7488), .ZN(O1541));
  INVX1 G42485 (.I(W25995), .ZN(W32608));
  INVX1 G42486 (.I(I174), .ZN(W18230));
  INVX1 G42487 (.I(W17121), .ZN(W18231));
  INVX1 G42488 (.I(W8509), .ZN(W32622));
  INVX1 G42489 (.I(W14528), .ZN(W18240));
  INVX1 G42490 (.I(W19810), .ZN(O6316));
  INVX1 G42491 (.I(W24943), .ZN(O6315));
  INVX1 G42492 (.I(I727), .ZN(W18243));
  INVX1 G42493 (.I(W31167), .ZN(O6313));
  INVX1 G42494 (.I(W4667), .ZN(W18244));
  INVX1 G42495 (.I(W6926), .ZN(W18300));
  INVX1 G42496 (.I(W2787), .ZN(O6310));
  INVX1 G42497 (.I(W11398), .ZN(W32606));
  INVX1 G42498 (.I(W9839), .ZN(O1528));
  INVX1 G42499 (.I(I1942), .ZN(W18255));
  INVX1 G42500 (.I(W18186), .ZN(W32600));
  INVX1 G42501 (.I(W18235), .ZN(W18258));
  INVX1 G42502 (.I(W10013), .ZN(W18259));
  INVX1 G42503 (.I(I505), .ZN(W18261));
  INVX1 G42504 (.I(W7821), .ZN(W32592));
  INVX1 G42505 (.I(W22336), .ZN(W32510));
  INVX1 G42506 (.I(W1320), .ZN(W18329));
  INVX1 G42507 (.I(W14928), .ZN(W18332));
  INVX1 G42508 (.I(W11217), .ZN(O1549));
  INVX1 G42509 (.I(W6855), .ZN(W32519));
  INVX1 G42510 (.I(W4148), .ZN(O6266));
  INVX1 G42511 (.I(W30388), .ZN(O6263));
  INVX1 G42512 (.I(W113), .ZN(W32514));
  INVX1 G42513 (.I(W4021), .ZN(W18340));
  INVX1 G42514 (.I(W796), .ZN(W18342));
  INVX1 G42515 (.I(W3717), .ZN(W18326));
  INVX1 G42516 (.I(I1658), .ZN(W18345));
  INVX1 G42517 (.I(W10874), .ZN(O1553));
  INVX1 G42518 (.I(W6754), .ZN(W18349));
  INVX1 G42519 (.I(W13933), .ZN(W32503));
  INVX1 G42520 (.I(W28459), .ZN(W32498));
  INVX1 G42521 (.I(W12115), .ZN(W18357));
  INVX1 G42522 (.I(W6836), .ZN(W18360));
  INVX1 G42523 (.I(W5730), .ZN(W32494));
  INVX1 G42524 (.I(W26308), .ZN(W32492));
  INVX1 G42525 (.I(I898), .ZN(W18305));
  INVX1 G42526 (.I(W25592), .ZN(W32554));
  INVX1 G42527 (.I(W28634), .ZN(W32553));
  INVX1 G42528 (.I(W28840), .ZN(W32552));
  INVX1 G42529 (.I(W11711), .ZN(W18303));
  INVX1 G42530 (.I(I1141), .ZN(O6282));
  INVX1 G42531 (.I(W18728), .ZN(O6281));
  INVX1 G42532 (.I(W12313), .ZN(O6280));
  INVX1 G42533 (.I(W134), .ZN(W18304));
  INVX1 G42534 (.I(W18008), .ZN(W32545));
  INVX1 G42535 (.I(W10077), .ZN(W18229));
  INVX1 G42536 (.I(W4475), .ZN(W18309));
  INVX1 G42537 (.I(W2075), .ZN(W18311));
  INVX1 G42538 (.I(W17570), .ZN(O6274));
  INVX1 G42539 (.I(W15819), .ZN(W18312));
  INVX1 G42540 (.I(W26430), .ZN(W32534));
  INVX1 G42541 (.I(W6928), .ZN(W32531));
  INVX1 G42542 (.I(W12790), .ZN(O1544));
  INVX1 G42543 (.I(W29719), .ZN(W32529));
  INVX1 G42544 (.I(W11933), .ZN(W18321));
  INVX1 G42545 (.I(W10795), .ZN(W18169));
  INVX1 G42546 (.I(W14482), .ZN(O6353));
  INVX1 G42547 (.I(W757), .ZN(W18158));
  INVX1 G42548 (.I(I1167), .ZN(O6352));
  INVX1 G42549 (.I(W14642), .ZN(O6351));
  INVX1 G42550 (.I(W5401), .ZN(W18160));
  INVX1 G42551 (.I(W6264), .ZN(O6350));
  INVX1 G42552 (.I(W18168), .ZN(W32692));
  INVX1 G42553 (.I(W5496), .ZN(W32690));
  INVX1 G42554 (.I(W12975), .ZN(W18167));
  INVX1 G42555 (.I(W17826), .ZN(W18156));
  INVX1 G42556 (.I(W6463), .ZN(O6348));
  INVX1 G42557 (.I(W3747), .ZN(O1514));
  INVX1 G42558 (.I(W11193), .ZN(W18173));
  INVX1 G42559 (.I(W13405), .ZN(W18174));
  INVX1 G42560 (.I(W19150), .ZN(O6345));
  INVX1 G42561 (.I(W18144), .ZN(W18178));
  INVX1 G42562 (.I(W10748), .ZN(W18179));
  INVX1 G42563 (.I(W3172), .ZN(O6342));
  INVX1 G42564 (.I(W23678), .ZN(O6341));
  INVX1 G42565 (.I(W9072), .ZN(W18140));
  INVX1 G42566 (.I(W17196), .ZN(W18130));
  INVX1 G42567 (.I(W14577), .ZN(W18132));
  INVX1 G42568 (.I(W15742), .ZN(W18133));
  INVX1 G42569 (.I(W10630), .ZN(W18134));
  INVX1 G42570 (.I(W14743), .ZN(W18135));
  INVX1 G42571 (.I(W1272), .ZN(W18136));
  INVX1 G42572 (.I(I1824), .ZN(W32716));
  INVX1 G42573 (.I(W27931), .ZN(W32715));
  INVX1 G42574 (.I(W812), .ZN(W32714));
  INVX1 G42575 (.I(W17839), .ZN(O1515));
  INVX1 G42576 (.I(W30738), .ZN(O6361));
  INVX1 G42577 (.I(W32483), .ZN(O6360));
  INVX1 G42578 (.I(W26233), .ZN(W32707));
  INVX1 G42579 (.I(W31820), .ZN(O6359));
  INVX1 G42580 (.I(W14091), .ZN(W18148));
  INVX1 G42581 (.I(W13153), .ZN(W18151));
  INVX1 G42582 (.I(W1795), .ZN(W18153));
  INVX1 G42583 (.I(I1596), .ZN(O6356));
  INVX1 G42584 (.I(W10779), .ZN(W18154));
  INVX1 G42585 (.I(W2810), .ZN(W18215));
  INVX1 G42586 (.I(W3120), .ZN(W18208));
  INVX1 G42587 (.I(W13251), .ZN(O6328));
  INVX1 G42588 (.I(W13983), .ZN(W18210));
  INVX1 G42589 (.I(I991), .ZN(W32643));
  INVX1 G42590 (.I(W18204), .ZN(W18212));
  INVX1 G42591 (.I(W4833), .ZN(W18213));
  INVX1 G42592 (.I(W9378), .ZN(W18214));
  INVX1 G42593 (.I(W31656), .ZN(O6326));
  INVX1 G42594 (.I(W15237), .ZN(O6325));
  INVX1 G42595 (.I(W31964), .ZN(W32649));
  INVX1 G42596 (.I(W17023), .ZN(W18217));
  INVX1 G42597 (.I(W15736), .ZN(O6324));
  INVX1 G42598 (.I(W17829), .ZN(W18220));
  INVX1 G42599 (.I(W1900), .ZN(W18221));
  INVX1 G42600 (.I(W12440), .ZN(O6322));
  INVX1 G42601 (.I(W29718), .ZN(W32630));
  INVX1 G42602 (.I(W9800), .ZN(W18222));
  INVX1 G42603 (.I(W3379), .ZN(W18223));
  INVX1 G42604 (.I(W969), .ZN(O1521));
  INVX1 G42605 (.I(W1952), .ZN(W18192));
  INVX1 G42606 (.I(W7), .ZN(O6339));
  INVX1 G42607 (.I(W6137), .ZN(O6338));
  INVX1 G42608 (.I(W10363), .ZN(W18183));
  INVX1 G42609 (.I(W31941), .ZN(W32672));
  INVX1 G42610 (.I(W27415), .ZN(W32671));
  INVX1 G42611 (.I(W18115), .ZN(O1516));
  INVX1 G42612 (.I(I903), .ZN(O6337));
  INVX1 G42613 (.I(W607), .ZN(O6336));
  INVX1 G42614 (.I(I1310), .ZN(W18191));
  INVX1 G42615 (.I(W23290), .ZN(W32003));
  INVX1 G42616 (.I(W5466), .ZN(W18193));
  INVX1 G42617 (.I(W12613), .ZN(W18194));
  INVX1 G42618 (.I(W12714), .ZN(W18198));
  INVX1 G42619 (.I(W1512), .ZN(W18201));
  INVX1 G42620 (.I(W15923), .ZN(W18202));
  INVX1 G42621 (.I(W24036), .ZN(W32654));
  INVX1 G42622 (.I(W8884), .ZN(O6332));
  INVX1 G42623 (.I(W32399), .ZN(W32651));
  INVX1 G42624 (.I(W7299), .ZN(W18204));
  INVX1 G42625 (.I(I1334), .ZN(O5754));
  INVX1 G42626 (.I(W1428), .ZN(W31382));
  INVX1 G42627 (.I(W12374), .ZN(W19453));
  INVX1 G42628 (.I(I1255), .ZN(O1778));
  INVX1 G42629 (.I(W10125), .ZN(O5758));
  INVX1 G42630 (.I(W4126), .ZN(W31375));
  INVX1 G42631 (.I(W6648), .ZN(W19458));
  INVX1 G42632 (.I(W21368), .ZN(W31370));
  INVX1 G42633 (.I(W12196), .ZN(W19462));
  INVX1 G42634 (.I(W4152), .ZN(W31368));
  INVX1 G42635 (.I(W6968), .ZN(W31367));
  INVX1 G42636 (.I(W18666), .ZN(W19450));
  INVX1 G42637 (.I(W22912), .ZN(O5753));
  INVX1 G42638 (.I(W21209), .ZN(W31363));
  INVX1 G42639 (.I(W15841), .ZN(W19468));
  INVX1 G42640 (.I(W16969), .ZN(W31360));
  INVX1 G42641 (.I(W7839), .ZN(O1780));
  INVX1 G42642 (.I(W11291), .ZN(W31357));
  INVX1 G42643 (.I(W10956), .ZN(W19478));
  INVX1 G42644 (.I(W9917), .ZN(O5749));
  INVX1 G42645 (.I(W15428), .ZN(W19479));
  INVX1 G42646 (.I(W3303), .ZN(O1772));
  INVX1 G42647 (.I(W31114), .ZN(O5776));
  INVX1 G42648 (.I(W351), .ZN(W19417));
  INVX1 G42649 (.I(W28398), .ZN(W31411));
  INVX1 G42650 (.I(W20912), .ZN(O5774));
  INVX1 G42651 (.I(W2831), .ZN(W31409));
  INVX1 G42652 (.I(W8350), .ZN(O1770));
  INVX1 G42653 (.I(W3297), .ZN(W19423));
  INVX1 G42654 (.I(W16225), .ZN(W31402));
  INVX1 G42655 (.I(W12071), .ZN(W19424));
  INVX1 G42656 (.I(W4940), .ZN(W19480));
  INVX1 G42657 (.I(W21180), .ZN(W31398));
  INVX1 G42658 (.I(W7571), .ZN(W19430));
  INVX1 G42659 (.I(W11626), .ZN(O1774));
  INVX1 G42660 (.I(W5709), .ZN(W19436));
  INVX1 G42661 (.I(I1509), .ZN(O5766));
  INVX1 G42662 (.I(I388), .ZN(O5763));
  INVX1 G42663 (.I(W12584), .ZN(W19442));
  INVX1 G42664 (.I(W7168), .ZN(W31387));
  INVX1 G42665 (.I(W18495), .ZN(W31384));
  INVX1 G42666 (.I(W11060), .ZN(O5730));
  INVX1 G42667 (.I(W1083), .ZN(W19516));
  INVX1 G42668 (.I(W3653), .ZN(W19517));
  INVX1 G42669 (.I(W7819), .ZN(W31315));
  INVX1 G42670 (.I(W13640), .ZN(W19519));
  INVX1 G42671 (.I(W9249), .ZN(W31313));
  INVX1 G42672 (.I(W8589), .ZN(O1789));
  INVX1 G42673 (.I(W16943), .ZN(W19522));
  INVX1 G42674 (.I(W18292), .ZN(O5732));
  INVX1 G42675 (.I(W9396), .ZN(O1790));
  INVX1 G42676 (.I(W16467), .ZN(W31318));
  INVX1 G42677 (.I(W10397), .ZN(W19526));
  INVX1 G42678 (.I(W3303), .ZN(W19529));
  INVX1 G42679 (.I(W10390), .ZN(W19531));
  INVX1 G42680 (.I(W3000), .ZN(W31299));
  INVX1 G42681 (.I(W1056), .ZN(W19535));
  INVX1 G42682 (.I(W30420), .ZN(W31297));
  INVX1 G42683 (.I(W9860), .ZN(O5725));
  INVX1 G42684 (.I(W13344), .ZN(W31295));
  INVX1 G42685 (.I(W6568), .ZN(W19536));
  INVX1 G42686 (.I(I1710), .ZN(W19500));
  INVX1 G42687 (.I(W3605), .ZN(W19481));
  INVX1 G42688 (.I(W15921), .ZN(O1781));
  INVX1 G42689 (.I(W5959), .ZN(W19484));
  INVX1 G42690 (.I(W24407), .ZN(O5747));
  INVX1 G42691 (.I(W7529), .ZN(W31344));
  INVX1 G42692 (.I(W27715), .ZN(O5746));
  INVX1 G42693 (.I(W5109), .ZN(W19489));
  INVX1 G42694 (.I(W29222), .ZN(W31338));
  INVX1 G42695 (.I(W11078), .ZN(O1783));
  INVX1 G42696 (.I(W12333), .ZN(O1769));
  INVX1 G42697 (.I(W24299), .ZN(O5741));
  INVX1 G42698 (.I(W4787), .ZN(W19503));
  INVX1 G42699 (.I(W20849), .ZN(O5739));
  INVX1 G42700 (.I(W16437), .ZN(W19504));
  INVX1 G42701 (.I(W21508), .ZN(O5738));
  INVX1 G42702 (.I(W18396), .ZN(W19507));
  INVX1 G42703 (.I(W15390), .ZN(W19512));
  INVX1 G42704 (.I(W8705), .ZN(O5735));
  INVX1 G42705 (.I(W2093), .ZN(W19513));
  INVX1 G42706 (.I(W1099), .ZN(W19333));
  INVX1 G42707 (.I(W1557), .ZN(O5813));
  INVX1 G42708 (.I(W1262), .ZN(W31496));
  INVX1 G42709 (.I(W17813), .ZN(W31494));
  INVX1 G42710 (.I(W25821), .ZN(O5811));
  INVX1 G42711 (.I(W1140), .ZN(W19329));
  INVX1 G42712 (.I(W1726), .ZN(O5810));
  INVX1 G42713 (.I(I1029), .ZN(W31489));
  INVX1 G42714 (.I(W8868), .ZN(W19332));
  INVX1 G42715 (.I(W24998), .ZN(W31486));
  INVX1 G42716 (.I(W2066), .ZN(W19327));
  INVX1 G42717 (.I(W16679), .ZN(W19336));
  INVX1 G42718 (.I(W5447), .ZN(W31482));
  INVX1 G42719 (.I(W16568), .ZN(W31481));
  INVX1 G42720 (.I(W2917), .ZN(W19337));
  INVX1 G42721 (.I(W5380), .ZN(W19338));
  INVX1 G42722 (.I(W1950), .ZN(W19339));
  INVX1 G42723 (.I(W6652), .ZN(W31477));
  INVX1 G42724 (.I(W3166), .ZN(O5804));
  INVX1 G42725 (.I(W14900), .ZN(W19341));
  INVX1 G42726 (.I(W11934), .ZN(W19309));
  INVX1 G42727 (.I(W11168), .ZN(O5825));
  INVX1 G42728 (.I(W3445), .ZN(W19289));
  INVX1 G42729 (.I(W26655), .ZN(W31524));
  INVX1 G42730 (.I(W2543), .ZN(W19292));
  INVX1 G42731 (.I(W28286), .ZN(O5822));
  INVX1 G42732 (.I(W11837), .ZN(W31515));
  INVX1 G42733 (.I(W7065), .ZN(W19306));
  INVX1 G42734 (.I(W10269), .ZN(W31513));
  INVX1 G42735 (.I(W8104), .ZN(W19308));
  INVX1 G42736 (.I(W11650), .ZN(W19350));
  INVX1 G42737 (.I(W29385), .ZN(W31510));
  INVX1 G42738 (.I(W4000), .ZN(W19310));
  INVX1 G42739 (.I(W19082), .ZN(W19313));
  INVX1 G42740 (.I(W10549), .ZN(W19315));
  INVX1 G42741 (.I(W19915), .ZN(W31506));
  INVX1 G42742 (.I(W13135), .ZN(W19321));
  INVX1 G42743 (.I(W3556), .ZN(W19322));
  INVX1 G42744 (.I(W4931), .ZN(W31502));
  INVX1 G42745 (.I(I20), .ZN(W19325));
  INVX1 G42746 (.I(W5545), .ZN(W19404));
  INVX1 G42747 (.I(I1113), .ZN(O5790));
  INVX1 G42748 (.I(W1411), .ZN(O1762));
  INVX1 G42749 (.I(W7078), .ZN(O1763));
  INVX1 G42750 (.I(W13076), .ZN(W31438));
  INVX1 G42751 (.I(W286), .ZN(W19395));
  INVX1 G42752 (.I(W31385), .ZN(O5788));
  INVX1 G42753 (.I(W899), .ZN(W31435));
  INVX1 G42754 (.I(W5375), .ZN(O1764));
  INVX1 G42755 (.I(W17292), .ZN(O1766));
  INVX1 G42756 (.I(W14410), .ZN(W19389));
  INVX1 G42757 (.I(W28278), .ZN(O5783));
  INVX1 G42758 (.I(W7941), .ZN(W19406));
  INVX1 G42759 (.I(W11207), .ZN(W19408));
  INVX1 G42760 (.I(W10960), .ZN(O1767));
  INVX1 G42761 (.I(W3463), .ZN(O1768));
  INVX1 G42762 (.I(W19855), .ZN(O5781));
  INVX1 G42763 (.I(W26747), .ZN(O5779));
  INVX1 G42764 (.I(W27554), .ZN(O5778));
  INVX1 G42765 (.I(I2), .ZN(W31416));
  INVX1 G42766 (.I(W12173), .ZN(W19371));
  INVX1 G42767 (.I(W4455), .ZN(W19352));
  INVX1 G42768 (.I(W4709), .ZN(W19353));
  INVX1 G42769 (.I(W14513), .ZN(O1751));
  INVX1 G42770 (.I(W26734), .ZN(O5802));
  INVX1 G42771 (.I(I875), .ZN(O1752));
  INVX1 G42772 (.I(W30918), .ZN(O5800));
  INVX1 G42773 (.I(W10671), .ZN(W19362));
  INVX1 G42774 (.I(W9537), .ZN(W19363));
  INVX1 G42775 (.I(W14523), .ZN(O5798));
  INVX1 G42776 (.I(W3062), .ZN(W19537));
  INVX1 G42777 (.I(W16343), .ZN(W19375));
  INVX1 G42778 (.I(W16258), .ZN(W31452));
  INVX1 G42779 (.I(W4379), .ZN(W19376));
  INVX1 G42780 (.I(W15479), .ZN(W19379));
  INVX1 G42781 (.I(W18849), .ZN(W19383));
  INVX1 G42782 (.I(W20614), .ZN(W31447));
  INVX1 G42783 (.I(W130), .ZN(O1760));
  INVX1 G42784 (.I(W13320), .ZN(W31445));
  INVX1 G42785 (.I(W16278), .ZN(W19386));
  INVX1 G42786 (.I(W11815), .ZN(O5654));
  INVX1 G42787 (.I(W30583), .ZN(O5661));
  INVX1 G42788 (.I(W17779), .ZN(O1825));
  INVX1 G42789 (.I(I288), .ZN(W19693));
  INVX1 G42790 (.I(W15374), .ZN(O5659));
  INVX1 G42791 (.I(W2204), .ZN(O1826));
  INVX1 G42792 (.I(W13432), .ZN(O1827));
  INVX1 G42793 (.I(W16702), .ZN(W19696));
  INVX1 G42794 (.I(W11656), .ZN(O5657));
  INVX1 G42795 (.I(W14065), .ZN(O5656));
  INVX1 G42796 (.I(W13537), .ZN(O1828));
  INVX1 G42797 (.I(I195), .ZN(O1824));
  INVX1 G42798 (.I(W10047), .ZN(W31133));
  INVX1 G42799 (.I(W15180), .ZN(W31132));
  INVX1 G42800 (.I(W1841), .ZN(O5652));
  INVX1 G42801 (.I(W529), .ZN(W19704));
  INVX1 G42802 (.I(W24708), .ZN(W31128));
  INVX1 G42803 (.I(W7870), .ZN(W19709));
  INVX1 G42804 (.I(W10992), .ZN(O1831));
  INVX1 G42805 (.I(W23621), .ZN(W31123));
  INVX1 G42806 (.I(W21893), .ZN(W31121));
  INVX1 G42807 (.I(W25133), .ZN(O5669));
  INVX1 G42808 (.I(W25029), .ZN(W31178));
  INVX1 G42809 (.I(I1888), .ZN(O1817));
  INVX1 G42810 (.I(W20227), .ZN(W31176));
  INVX1 G42811 (.I(W31031), .ZN(O5673));
  INVX1 G42812 (.I(W19029), .ZN(W19665));
  INVX1 G42813 (.I(W7406), .ZN(W31171));
  INVX1 G42814 (.I(W13963), .ZN(W19670));
  INVX1 G42815 (.I(W17693), .ZN(W31168));
  INVX1 G42816 (.I(W16776), .ZN(W31166));
  INVX1 G42817 (.I(W26066), .ZN(W31120));
  INVX1 G42818 (.I(W5438), .ZN(W19676));
  INVX1 G42819 (.I(W711), .ZN(W31162));
  INVX1 G42820 (.I(W18388), .ZN(W19677));
  INVX1 G42821 (.I(W995), .ZN(W31159));
  INVX1 G42822 (.I(I990), .ZN(W19679));
  INVX1 G42823 (.I(I1894), .ZN(W31155));
  INVX1 G42824 (.I(W3465), .ZN(W31152));
  INVX1 G42825 (.I(W24229), .ZN(W31151));
  INVX1 G42826 (.I(W27439), .ZN(O5664));
  INVX1 G42827 (.I(W8940), .ZN(W31076));
  INVX1 G42828 (.I(W12107), .ZN(O5641));
  INVX1 G42829 (.I(W9184), .ZN(W19738));
  INVX1 G42830 (.I(I1939), .ZN(W19739));
  INVX1 G42831 (.I(W7034), .ZN(W31091));
  INVX1 G42832 (.I(W16654), .ZN(W19740));
  INVX1 G42833 (.I(W19579), .ZN(W31085));
  INVX1 G42834 (.I(W8907), .ZN(O5635));
  INVX1 G42835 (.I(W6368), .ZN(W31078));
  INVX1 G42836 (.I(W15687), .ZN(W19758));
  INVX1 G42837 (.I(I1399), .ZN(O1840));
  INVX1 G42838 (.I(W18637), .ZN(W31074));
  INVX1 G42839 (.I(W16303), .ZN(W19762));
  INVX1 G42840 (.I(W6613), .ZN(O5631));
  INVX1 G42841 (.I(W6671), .ZN(W19766));
  INVX1 G42842 (.I(W19281), .ZN(W19770));
  INVX1 G42843 (.I(W15754), .ZN(W19771));
  INVX1 G42844 (.I(W2758), .ZN(O1849));
  INVX1 G42845 (.I(W8331), .ZN(O5628));
  INVX1 G42846 (.I(W229), .ZN(W19778));
  INVX1 G42847 (.I(W25864), .ZN(O5646));
  INVX1 G42848 (.I(W16779), .ZN(W31119));
  INVX1 G42849 (.I(W7850), .ZN(W31117));
  INVX1 G42850 (.I(W13044), .ZN(W31115));
  INVX1 G42851 (.I(W3905), .ZN(W19716));
  INVX1 G42852 (.I(W20774), .ZN(W31113));
  INVX1 G42853 (.I(W19446), .ZN(W19719));
  INVX1 G42854 (.I(W2643), .ZN(O1833));
  INVX1 G42855 (.I(W7401), .ZN(W19723));
  INVX1 G42856 (.I(W9587), .ZN(W31108));
  INVX1 G42857 (.I(W3827), .ZN(O1816));
  INVX1 G42858 (.I(W6770), .ZN(W31106));
  INVX1 G42859 (.I(W3186), .ZN(O1835));
  INVX1 G42860 (.I(I743), .ZN(O1837));
  INVX1 G42861 (.I(W20925), .ZN(O5645));
  INVX1 G42862 (.I(W19712), .ZN(O1838));
  INVX1 G42863 (.I(W4519), .ZN(W31100));
  INVX1 G42864 (.I(W9406), .ZN(W19732));
  INVX1 G42865 (.I(W5347), .ZN(W19734));
  INVX1 G42866 (.I(W17687), .ZN(W31097));
  INVX1 G42867 (.I(W14093), .ZN(W31247));
  INVX1 G42868 (.I(W6085), .ZN(O1801));
  INVX1 G42869 (.I(W17372), .ZN(W19581));
  INVX1 G42870 (.I(W24996), .ZN(W31257));
  INVX1 G42871 (.I(W29595), .ZN(W31256));
  INVX1 G42872 (.I(W19436), .ZN(W19582));
  INVX1 G42873 (.I(W15905), .ZN(W19583));
  INVX1 G42874 (.I(W30576), .ZN(W31253));
  INVX1 G42875 (.I(W18116), .ZN(O1802));
  INVX1 G42876 (.I(W16375), .ZN(W19587));
  INVX1 G42877 (.I(W2153), .ZN(W31261));
  INVX1 G42878 (.I(W763), .ZN(O5708));
  INVX1 G42879 (.I(W16648), .ZN(W19597));
  INVX1 G42880 (.I(W5043), .ZN(W19598));
  INVX1 G42881 (.I(W1429), .ZN(O1806));
  INVX1 G42882 (.I(W15098), .ZN(W19601));
  INVX1 G42883 (.I(W3693), .ZN(W19602));
  INVX1 G42884 (.I(W16914), .ZN(O5703));
  INVX1 G42885 (.I(I371), .ZN(W19603));
  INVX1 G42886 (.I(W14980), .ZN(W31234));
  INVX1 G42887 (.I(W20839), .ZN(O5717));
  INVX1 G42888 (.I(W26413), .ZN(W31291));
  INVX1 G42889 (.I(W4902), .ZN(O5722));
  INVX1 G42890 (.I(W9075), .ZN(O1794));
  INVX1 G42891 (.I(W2366), .ZN(O5719));
  INVX1 G42892 (.I(W15212), .ZN(W19548));
  INVX1 G42893 (.I(W13388), .ZN(W19549));
  INVX1 G42894 (.I(W16586), .ZN(W31281));
  INVX1 G42895 (.I(W1449), .ZN(W31280));
  INVX1 G42896 (.I(W6606), .ZN(W19552));
  INVX1 G42897 (.I(W18102), .ZN(W19604));
  INVX1 G42898 (.I(W21260), .ZN(O5715));
  INVX1 G42899 (.I(W6369), .ZN(O1798));
  INVX1 G42900 (.I(W28950), .ZN(W31270));
  INVX1 G42901 (.I(W2694), .ZN(W19565));
  INVX1 G42902 (.I(W8857), .ZN(O1800));
  INVX1 G42903 (.I(W7814), .ZN(W31267));
  INVX1 G42904 (.I(W4939), .ZN(W19568));
  INVX1 G42905 (.I(I1256), .ZN(W19573));
  INVX1 G42906 (.I(W11468), .ZN(W19576));
  INVX1 G42907 (.I(W11004), .ZN(W19641));
  INVX1 G42908 (.I(W30317), .ZN(O5688));
  INVX1 G42909 (.I(I695), .ZN(W31202));
  INVX1 G42910 (.I(W29358), .ZN(O5687));
  INVX1 G42911 (.I(W913), .ZN(O5686));
  INVX1 G42912 (.I(W19227), .ZN(O5685));
  INVX1 G42913 (.I(W7088), .ZN(O1811));
  INVX1 G42914 (.I(W16278), .ZN(O5683));
  INVX1 G42915 (.I(W8175), .ZN(W19633));
  INVX1 G42916 (.I(W259), .ZN(W19636));
  INVX1 G42917 (.I(I317), .ZN(W19630));
  INVX1 G42918 (.I(W3470), .ZN(W19643));
  INVX1 G42919 (.I(W9084), .ZN(O5679));
  INVX1 G42920 (.I(W21191), .ZN(O5678));
  INVX1 G42921 (.I(W1126), .ZN(W19644));
  INVX1 G42922 (.I(W9711), .ZN(O5676));
  INVX1 G42923 (.I(W15796), .ZN(W19645));
  INVX1 G42924 (.I(W60), .ZN(W19656));
  INVX1 G42925 (.I(W4921), .ZN(W19657));
  INVX1 G42926 (.I(W3184), .ZN(W19658));
  INVX1 G42927 (.I(W10769), .ZN(O5697));
  INVX1 G42928 (.I(W28922), .ZN(O5701));
  INVX1 G42929 (.I(W7254), .ZN(W31230));
  INVX1 G42930 (.I(W1771), .ZN(W19607));
  INVX1 G42931 (.I(W11508), .ZN(W31228));
  INVX1 G42932 (.I(W29716), .ZN(W31226));
  INVX1 G42933 (.I(W6862), .ZN(W19610));
  INVX1 G42934 (.I(W22687), .ZN(W31223));
  INVX1 G42935 (.I(W20602), .ZN(O5698));
  INVX1 G42936 (.I(W1377), .ZN(W31221));
  INVX1 G42937 (.I(W6441), .ZN(O5826));
  INVX1 G42938 (.I(W26902), .ZN(O5696));
  INVX1 G42939 (.I(W14139), .ZN(O5695));
  INVX1 G42940 (.I(W13845), .ZN(W19614));
  INVX1 G42941 (.I(W13254), .ZN(O1808));
  INVX1 G42942 (.I(W2280), .ZN(O5692));
  INVX1 G42943 (.I(W11232), .ZN(W19617));
  INVX1 G42944 (.I(W15091), .ZN(O5691));
  INVX1 G42945 (.I(W1208), .ZN(W19625));
  INVX1 G42946 (.I(W2401), .ZN(W19626));
  INVX1 G42947 (.I(W23760), .ZN(W31844));
  INVX1 G42948 (.I(W21146), .ZN(O5981));
  INVX1 G42949 (.I(W21730), .ZN(O5980));
  INVX1 G42950 (.I(W7679), .ZN(O5979));
  INVX1 G42951 (.I(W1805), .ZN(O1686));
  INVX1 G42952 (.I(W8967), .ZN(O5977));
  INVX1 G42953 (.I(I1759), .ZN(W18984));
  INVX1 G42954 (.I(W15741), .ZN(W31851));
  INVX1 G42955 (.I(W2416), .ZN(W31850));
  INVX1 G42956 (.I(W10838), .ZN(W31846));
  INVX1 G42957 (.I(W8523), .ZN(W18994));
  INVX1 G42958 (.I(W18863), .ZN(O5982));
  INVX1 G42959 (.I(W4549), .ZN(W19001));
  INVX1 G42960 (.I(W30187), .ZN(W31841));
  INVX1 G42961 (.I(W2209), .ZN(O5972));
  INVX1 G42962 (.I(W26611), .ZN(O5970));
  INVX1 G42963 (.I(W12431), .ZN(W19004));
  INVX1 G42964 (.I(W6466), .ZN(W19005));
  INVX1 G42965 (.I(W6377), .ZN(W19007));
  INVX1 G42966 (.I(I152), .ZN(W19008));
  INVX1 G42967 (.I(W17466), .ZN(O5968));
  INVX1 G42968 (.I(W2610), .ZN(W18968));
  INVX1 G42969 (.I(W16993), .ZN(W31890));
  INVX1 G42970 (.I(W2798), .ZN(W31888));
  INVX1 G42971 (.I(W4689), .ZN(O5997));
  INVX1 G42972 (.I(W17554), .ZN(W31885));
  INVX1 G42973 (.I(W25362), .ZN(W31880));
  INVX1 G42974 (.I(W19093), .ZN(O5994));
  INVX1 G42975 (.I(W18274), .ZN(O5993));
  INVX1 G42976 (.I(W6207), .ZN(W18964));
  INVX1 G42977 (.I(W5159), .ZN(W18967));
  INVX1 G42978 (.I(W28079), .ZN(O5967));
  INVX1 G42979 (.I(W22676), .ZN(W31871));
  INVX1 G42980 (.I(W888), .ZN(O5990));
  INVX1 G42981 (.I(W14622), .ZN(W18972));
  INVX1 G42982 (.I(W30128), .ZN(O5988));
  INVX1 G42983 (.I(W13384), .ZN(O5987));
  INVX1 G42984 (.I(W8541), .ZN(O5986));
  INVX1 G42985 (.I(W11646), .ZN(O5985));
  INVX1 G42986 (.I(W8652), .ZN(W18975));
  INVX1 G42987 (.I(W7957), .ZN(W18976));
  INVX1 G42988 (.I(W4291), .ZN(O5938));
  INVX1 G42989 (.I(W7312), .ZN(W19047));
  INVX1 G42990 (.I(W15509), .ZN(W31793));
  INVX1 G42991 (.I(W4033), .ZN(W19051));
  INVX1 G42992 (.I(W10201), .ZN(W19054));
  INVX1 G42993 (.I(W20769), .ZN(W31788));
  INVX1 G42994 (.I(W15734), .ZN(O5945));
  INVX1 G42995 (.I(W15100), .ZN(W19056));
  INVX1 G42996 (.I(W12788), .ZN(W19058));
  INVX1 G42997 (.I(I1206), .ZN(O5939));
  INVX1 G42998 (.I(W8390), .ZN(O1695));
  INVX1 G42999 (.I(W3599), .ZN(W19066));
  INVX1 G43000 (.I(W25467), .ZN(W31774));
  INVX1 G43001 (.I(W6001), .ZN(W19068));
  INVX1 G43002 (.I(W17767), .ZN(O5936));
  INVX1 G43003 (.I(I626), .ZN(W19071));
  INVX1 G43004 (.I(W29335), .ZN(W31768));
  INVX1 G43005 (.I(W21979), .ZN(O5934));
  INVX1 G43006 (.I(I1475), .ZN(W31765));
  INVX1 G43007 (.I(W18477), .ZN(W19073));
  INVX1 G43008 (.I(W503), .ZN(W19033));
  INVX1 G43009 (.I(W3672), .ZN(W19011));
  INVX1 G43010 (.I(W19415), .ZN(W31829));
  INVX1 G43011 (.I(W29144), .ZN(W31827));
  INVX1 G43012 (.I(W8437), .ZN(O5964));
  INVX1 G43013 (.I(W1932), .ZN(W31820));
  INVX1 G43014 (.I(W20992), .ZN(W31817));
  INVX1 G43015 (.I(W2250), .ZN(W31816));
  INVX1 G43016 (.I(W31016), .ZN(O5960));
  INVX1 G43017 (.I(W3321), .ZN(W19028));
  INVX1 G43018 (.I(W23368), .ZN(W31891));
  INVX1 G43019 (.I(W4590), .ZN(W19036));
  INVX1 G43020 (.I(W17839), .ZN(W19039));
  INVX1 G43021 (.I(W19436), .ZN(O5955));
  INVX1 G43022 (.I(W13783), .ZN(W19040));
  INVX1 G43023 (.I(W23126), .ZN(O5954));
  INVX1 G43024 (.I(W2246), .ZN(O5953));
  INVX1 G43025 (.I(W10787), .ZN(W19042));
  INVX1 G43026 (.I(W10216), .ZN(O5951));
  INVX1 G43027 (.I(W10438), .ZN(W19045));
  INVX1 G43028 (.I(W15360), .ZN(W18886));
  INVX1 G43029 (.I(W6937), .ZN(W18877));
  INVX1 G43030 (.I(W7787), .ZN(O1667));
  INVX1 G43031 (.I(W19709), .ZN(W31971));
  INVX1 G43032 (.I(W15520), .ZN(W31970));
  INVX1 G43033 (.I(W3558), .ZN(W31968));
  INVX1 G43034 (.I(W3867), .ZN(W31967));
  INVX1 G43035 (.I(W325), .ZN(O1669));
  INVX1 G43036 (.I(W1992), .ZN(W18883));
  INVX1 G43037 (.I(I103), .ZN(O1670));
  INVX1 G43038 (.I(W7898), .ZN(O6031));
  INVX1 G43039 (.I(W18474), .ZN(W18888));
  INVX1 G43040 (.I(W23216), .ZN(O6026));
  INVX1 G43041 (.I(W4692), .ZN(W18890));
  INVX1 G43042 (.I(W29124), .ZN(O6025));
  INVX1 G43043 (.I(W31225), .ZN(W31957));
  INVX1 G43044 (.I(I24), .ZN(O6024));
  INVX1 G43045 (.I(W4897), .ZN(W31955));
  INVX1 G43046 (.I(W21342), .ZN(O6023));
  INVX1 G43047 (.I(W11723), .ZN(W31952));
  INVX1 G43048 (.I(W13497), .ZN(W18859));
  INVX1 G43049 (.I(W8194), .ZN(W18846));
  INVX1 G43050 (.I(W3192), .ZN(O6045));
  INVX1 G43051 (.I(W4800), .ZN(O6044));
  INVX1 G43052 (.I(W15318), .ZN(W18849));
  INVX1 G43053 (.I(W26624), .ZN(O6041));
  INVX1 G43054 (.I(W9552), .ZN(W18851));
  INVX1 G43055 (.I(W31243), .ZN(W31994));
  INVX1 G43056 (.I(W1788), .ZN(O1662));
  INVX1 G43057 (.I(W26238), .ZN(O6037));
  INVX1 G43058 (.I(W22248), .ZN(W31950));
  INVX1 G43059 (.I(W20630), .ZN(O6036));
  INVX1 G43060 (.I(W9713), .ZN(W18862));
  INVX1 G43061 (.I(W4573), .ZN(W18863));
  INVX1 G43062 (.I(W10702), .ZN(W18864));
  INVX1 G43063 (.I(W4299), .ZN(W18869));
  INVX1 G43064 (.I(W7086), .ZN(W31980));
  INVX1 G43065 (.I(W5900), .ZN(W18874));
  INVX1 G43066 (.I(W12481), .ZN(W31977));
  INVX1 G43067 (.I(W6575), .ZN(W18876));
  INVX1 G43068 (.I(W15928), .ZN(W31903));
  INVX1 G43069 (.I(W4778), .ZN(O6012));
  INVX1 G43070 (.I(W27405), .ZN(W31920));
  INVX1 G43071 (.I(W511), .ZN(W18929));
  INVX1 G43072 (.I(W5039), .ZN(O6008));
  INVX1 G43073 (.I(W12095), .ZN(W18936));
  INVX1 G43074 (.I(W2681), .ZN(W31911));
  INVX1 G43075 (.I(W8484), .ZN(W18939));
  INVX1 G43076 (.I(W11489), .ZN(W31907));
  INVX1 G43077 (.I(W4762), .ZN(W18943));
  INVX1 G43078 (.I(W11777), .ZN(W18924));
  INVX1 G43079 (.I(W18943), .ZN(W18946));
  INVX1 G43080 (.I(W3799), .ZN(W18947));
  INVX1 G43081 (.I(W14118), .ZN(W18949));
  INVX1 G43082 (.I(W19716), .ZN(W31898));
  INVX1 G43083 (.I(W5776), .ZN(W18950));
  INVX1 G43084 (.I(W4356), .ZN(W18951));
  INVX1 G43085 (.I(W27923), .ZN(O6001));
  INVX1 G43086 (.I(W23693), .ZN(W31894));
  INVX1 G43087 (.I(W18526), .ZN(O6000));
  INVX1 G43088 (.I(W6537), .ZN(W18906));
  INVX1 G43089 (.I(W17864), .ZN(W31949));
  INVX1 G43090 (.I(W10643), .ZN(W18898));
  INVX1 G43091 (.I(W4867), .ZN(W18899));
  INVX1 G43092 (.I(W1288), .ZN(W18900));
  INVX1 G43093 (.I(W19664), .ZN(W31944));
  INVX1 G43094 (.I(W5595), .ZN(O6019));
  INVX1 G43095 (.I(I467), .ZN(O6018));
  INVX1 G43096 (.I(W2036), .ZN(O1675));
  INVX1 G43097 (.I(W19176), .ZN(W31940));
  INVX1 G43098 (.I(W2698), .ZN(O1699));
  INVX1 G43099 (.I(W24926), .ZN(W31937));
  INVX1 G43100 (.I(W9378), .ZN(W18911));
  INVX1 G43101 (.I(W4316), .ZN(W31933));
  INVX1 G43102 (.I(W10542), .ZN(O1677));
  INVX1 G43103 (.I(W30035), .ZN(O6015));
  INVX1 G43104 (.I(W25494), .ZN(W31930));
  INVX1 G43105 (.I(W9743), .ZN(W18915));
  INVX1 G43106 (.I(W11579), .ZN(W18918));
  INVX1 G43107 (.I(W19207), .ZN(W31924));
  INVX1 G43108 (.I(W12308), .ZN(W31596));
  INVX1 G43109 (.I(W3613), .ZN(W31613));
  INVX1 G43110 (.I(W11346), .ZN(W19223));
  INVX1 G43111 (.I(W14595), .ZN(O1729));
  INVX1 G43112 (.I(W21945), .ZN(W31609));
  INVX1 G43113 (.I(W10046), .ZN(W19228));
  INVX1 G43114 (.I(W24183), .ZN(W31604));
  INVX1 G43115 (.I(W8133), .ZN(W19233));
  INVX1 G43116 (.I(W30100), .ZN(W31600));
  INVX1 G43117 (.I(W9644), .ZN(W19238));
  INVX1 G43118 (.I(W8445), .ZN(O5853));
  INVX1 G43119 (.I(W1706), .ZN(W19221));
  INVX1 G43120 (.I(W514), .ZN(W31595));
  INVX1 G43121 (.I(W9821), .ZN(W19242));
  INVX1 G43122 (.I(W10426), .ZN(O5851));
  INVX1 G43123 (.I(I1593), .ZN(O1733));
  INVX1 G43124 (.I(W31308), .ZN(O5848));
  INVX1 G43125 (.I(W15439), .ZN(W31587));
  INVX1 G43126 (.I(W21278), .ZN(W31586));
  INVX1 G43127 (.I(W681), .ZN(W31585));
  INVX1 G43128 (.I(W25297), .ZN(W31584));
  INVX1 G43129 (.I(W1984), .ZN(W19209));
  INVX1 G43130 (.I(W25054), .ZN(W31644));
  INVX1 G43131 (.I(W4091), .ZN(W19195));
  INVX1 G43132 (.I(I1079), .ZN(W31642));
  INVX1 G43133 (.I(W15927), .ZN(O5870));
  INVX1 G43134 (.I(W751), .ZN(O5869));
  INVX1 G43135 (.I(W17253), .ZN(W31637));
  INVX1 G43136 (.I(W8114), .ZN(W19205));
  INVX1 G43137 (.I(W155), .ZN(O1725));
  INVX1 G43138 (.I(W10264), .ZN(W19207));
  INVX1 G43139 (.I(W26334), .ZN(W31583));
  INVX1 G43140 (.I(W1972), .ZN(O5865));
  INVX1 G43141 (.I(W2701), .ZN(O5864));
  INVX1 G43142 (.I(W13746), .ZN(W19214));
  INVX1 G43143 (.I(W13462), .ZN(O5863));
  INVX1 G43144 (.I(W7914), .ZN(W19215));
  INVX1 G43145 (.I(W14773), .ZN(W31621));
  INVX1 G43146 (.I(W31093), .ZN(W31619));
  INVX1 G43147 (.I(W13309), .ZN(W31617));
  INVX1 G43148 (.I(W2692), .ZN(W31616));
  INVX1 G43149 (.I(W20308), .ZN(W31545));
  INVX1 G43150 (.I(W3526), .ZN(W31557));
  INVX1 G43151 (.I(W5759), .ZN(W31556));
  INVX1 G43152 (.I(W3189), .ZN(W19264));
  INVX1 G43153 (.I(W20050), .ZN(O5838));
  INVX1 G43154 (.I(W11097), .ZN(O1737));
  INVX1 G43155 (.I(W4383), .ZN(W19268));
  INVX1 G43156 (.I(W10515), .ZN(O5835));
  INVX1 G43157 (.I(W14845), .ZN(W19271));
  INVX1 G43158 (.I(W3478), .ZN(W19273));
  INVX1 G43159 (.I(W28669), .ZN(W31559));
  INVX1 G43160 (.I(W17101), .ZN(O1739));
  INVX1 G43161 (.I(W11591), .ZN(O1740));
  INVX1 G43162 (.I(W29249), .ZN(W31542));
  INVX1 G43163 (.I(W27467), .ZN(W31541));
  INVX1 G43164 (.I(W20367), .ZN(W31540));
  INVX1 G43165 (.I(W27389), .ZN(O5830));
  INVX1 G43166 (.I(W12249), .ZN(O5829));
  INVX1 G43167 (.I(W16705), .ZN(W31535));
  INVX1 G43168 (.I(W22827), .ZN(W31534));
  INVX1 G43169 (.I(W20200), .ZN(O5842));
  INVX1 G43170 (.I(W1327), .ZN(W19249));
  INVX1 G43171 (.I(W13799), .ZN(W19251));
  INVX1 G43172 (.I(W16907), .ZN(W19254));
  INVX1 G43173 (.I(W13239), .ZN(W19255));
  INVX1 G43174 (.I(W10983), .ZN(W31576));
  INVX1 G43175 (.I(W27609), .ZN(O5844));
  INVX1 G43176 (.I(W12359), .ZN(O5843));
  INVX1 G43177 (.I(W23177), .ZN(W31573));
  INVX1 G43178 (.I(W7160), .ZN(W31572));
  INVX1 G43179 (.I(W25168), .ZN(O5872));
  INVX1 G43180 (.I(W23396), .ZN(W31570));
  INVX1 G43181 (.I(W21758), .ZN(W31569));
  INVX1 G43182 (.I(W14502), .ZN(W19260));
  INVX1 G43183 (.I(W23370), .ZN(O5841));
  INVX1 G43184 (.I(W3499), .ZN(W31564));
  INVX1 G43185 (.I(W9707), .ZN(W31563));
  INVX1 G43186 (.I(W12831), .ZN(W19262));
  INVX1 G43187 (.I(W15104), .ZN(O5840));
  INVX1 G43188 (.I(W21535), .ZN(W31560));
  INVX1 G43189 (.I(W23823), .ZN(W31717));
  INVX1 G43190 (.I(W14973), .ZN(W19105));
  INVX1 G43191 (.I(W14701), .ZN(W19106));
  INVX1 G43192 (.I(W13178), .ZN(W19107));
  INVX1 G43193 (.I(W13387), .ZN(W19110));
  INVX1 G43194 (.I(W13680), .ZN(W19111));
  INVX1 G43195 (.I(W13891), .ZN(W31724));
  INVX1 G43196 (.I(W24503), .ZN(O5911));
  INVX1 G43197 (.I(I1709), .ZN(O5910));
  INVX1 G43198 (.I(I257), .ZN(W19120));
  INVX1 G43199 (.I(W26005), .ZN(W31733));
  INVX1 G43200 (.I(W15898), .ZN(W19121));
  INVX1 G43201 (.I(W12549), .ZN(W19122));
  INVX1 G43202 (.I(W3120), .ZN(W19123));
  INVX1 G43203 (.I(W19974), .ZN(O5906));
  INVX1 G43204 (.I(I1557), .ZN(O1711));
  INVX1 G43205 (.I(W16593), .ZN(W19127));
  INVX1 G43206 (.I(W6321), .ZN(W19128));
  INVX1 G43207 (.I(W20680), .ZN(W31707));
  INVX1 G43208 (.I(W11139), .ZN(W19133));
  INVX1 G43209 (.I(W14361), .ZN(O5922));
  INVX1 G43210 (.I(W22112), .ZN(O5931));
  INVX1 G43211 (.I(W8958), .ZN(O1701));
  INVX1 G43212 (.I(W4376), .ZN(O5929));
  INVX1 G43213 (.I(W20437), .ZN(O5927));
  INVX1 G43214 (.I(W28994), .ZN(W31755));
  INVX1 G43215 (.I(W1674), .ZN(W19085));
  INVX1 G43216 (.I(W9016), .ZN(O1703));
  INVX1 G43217 (.I(W13043), .ZN(W31750));
  INVX1 G43218 (.I(I109), .ZN(O1706));
  INVX1 G43219 (.I(W1893), .ZN(O1713));
  INVX1 G43220 (.I(W15220), .ZN(W19095));
  INVX1 G43221 (.I(W29186), .ZN(W31742));
  INVX1 G43222 (.I(W15414), .ZN(W31741));
  INVX1 G43223 (.I(W16459), .ZN(W31740));
  INVX1 G43224 (.I(W551), .ZN(O1707));
  INVX1 G43225 (.I(W26265), .ZN(O5920));
  INVX1 G43226 (.I(W1054), .ZN(O5919));
  INVX1 G43227 (.I(W6632), .ZN(O5918));
  INVX1 G43228 (.I(I248), .ZN(W19102));
  INVX1 G43229 (.I(W19069), .ZN(O5880));
  INVX1 G43230 (.I(W23570), .ZN(O5889));
  INVX1 G43231 (.I(W8812), .ZN(W19171));
  INVX1 G43232 (.I(W2837), .ZN(W19176));
  INVX1 G43233 (.I(W31084), .ZN(O5883));
  INVX1 G43234 (.I(W12987), .ZN(W31663));
  INVX1 G43235 (.I(I496), .ZN(O5882));
  INVX1 G43236 (.I(W13983), .ZN(W19182));
  INVX1 G43237 (.I(I1378), .ZN(O5881));
  INVX1 G43238 (.I(W9939), .ZN(W19183));
  INVX1 G43239 (.I(W5800), .ZN(W31672));
  INVX1 G43240 (.I(W9903), .ZN(W19184));
  INVX1 G43241 (.I(W15506), .ZN(W19188));
  INVX1 G43242 (.I(W14852), .ZN(W19191));
  INVX1 G43243 (.I(W16499), .ZN(W19192));
  INVX1 G43244 (.I(W14719), .ZN(W31650));
  INVX1 G43245 (.I(W14481), .ZN(W19193));
  INVX1 G43246 (.I(W7256), .ZN(O5874));
  INVX1 G43247 (.I(W25410), .ZN(W31647));
  INVX1 G43248 (.I(I1838), .ZN(O5873));
  INVX1 G43249 (.I(W13304), .ZN(O1718));
  INVX1 G43250 (.I(W24734), .ZN(O5900));
  INVX1 G43251 (.I(W6069), .ZN(W19141));
  INVX1 G43252 (.I(W1749), .ZN(W31699));
  INVX1 G43253 (.I(W7434), .ZN(W19143));
  INVX1 G43254 (.I(W4690), .ZN(W31697));
  INVX1 G43255 (.I(W13986), .ZN(W31696));
  INVX1 G43256 (.I(W6297), .ZN(W19154));
  INVX1 G43257 (.I(W19497), .ZN(O5895));
  INVX1 G43258 (.I(W6231), .ZN(W19155));
  INVX1 G43259 (.I(I1958), .ZN(W21603));
  INVX1 G43260 (.I(W19130), .ZN(W19159));
  INVX1 G43261 (.I(W26068), .ZN(W31684));
  INVX1 G43262 (.I(W10534), .ZN(W19160));
  INVX1 G43263 (.I(W4116), .ZN(W19161));
  INVX1 G43264 (.I(W5882), .ZN(W19162));
  INVX1 G43265 (.I(W19726), .ZN(O5891));
  INVX1 G43266 (.I(W736), .ZN(W31678));
  INVX1 G43267 (.I(W17303), .ZN(W19167));
  INVX1 G43268 (.I(W5587), .ZN(W31675));
  INVX1 G43269 (.I(W18435), .ZN(W24128));
  INVX1 G43270 (.I(W23689), .ZN(W26624));
  INVX1 G43271 (.I(W21239), .ZN(W26623));
  INVX1 G43272 (.I(W12018), .ZN(O2977));
  INVX1 G43273 (.I(W24075), .ZN(W24117));
  INVX1 G43274 (.I(W22365), .ZN(O3811));
  INVX1 G43275 (.I(W1044), .ZN(W24118));
  INVX1 G43276 (.I(W21681), .ZN(W24122));
  INVX1 G43277 (.I(W1626), .ZN(W24125));
  INVX1 G43278 (.I(W19251), .ZN(O3808));
  INVX1 G43279 (.I(W5171), .ZN(W26613));
  INVX1 G43280 (.I(W17219), .ZN(W26625));
  INVX1 G43281 (.I(W15368), .ZN(O2979));
  INVX1 G43282 (.I(W16192), .ZN(W24133));
  INVX1 G43283 (.I(W24060), .ZN(W26603));
  INVX1 G43284 (.I(W21077), .ZN(W24140));
  INVX1 G43285 (.I(W309), .ZN(W26599));
  INVX1 G43286 (.I(W19276), .ZN(O2982));
  INVX1 G43287 (.I(W893), .ZN(O2987));
  INVX1 G43288 (.I(W6495), .ZN(W26593));
  INVX1 G43289 (.I(W17895), .ZN(O2988));
  INVX1 G43290 (.I(W8237), .ZN(W24096));
  INVX1 G43291 (.I(W2756), .ZN(W24081));
  INVX1 G43292 (.I(W23161), .ZN(W24082));
  INVX1 G43293 (.I(W25404), .ZN(O3822));
  INVX1 G43294 (.I(W10875), .ZN(W24085));
  INVX1 G43295 (.I(W8598), .ZN(O3820));
  INVX1 G43296 (.I(W25309), .ZN(O3819));
  INVX1 G43297 (.I(W16468), .ZN(W26649));
  INVX1 G43298 (.I(W8894), .ZN(W26646));
  INVX1 G43299 (.I(W14354), .ZN(O2968));
  INVX1 G43300 (.I(W13323), .ZN(W24156));
  INVX1 G43301 (.I(W19423), .ZN(W26640));
  INVX1 G43302 (.I(W22140), .ZN(W24098));
  INVX1 G43303 (.I(W1162), .ZN(W26638));
  INVX1 G43304 (.I(W8890), .ZN(W26635));
  INVX1 G43305 (.I(I1520), .ZN(O2972));
  INVX1 G43306 (.I(W16398), .ZN(O2974));
  INVX1 G43307 (.I(I915), .ZN(W26631));
  INVX1 G43308 (.I(W26356), .ZN(W26628));
  INVX1 G43309 (.I(W16514), .ZN(W26627));
  INVX1 G43310 (.I(W5191), .ZN(W26548));
  INVX1 G43311 (.I(W8855), .ZN(W26559));
  INVX1 G43312 (.I(W7704), .ZN(W24192));
  INVX1 G43313 (.I(I1642), .ZN(O3794));
  INVX1 G43314 (.I(I258), .ZN(W24199));
  INVX1 G43315 (.I(W6735), .ZN(W24200));
  INVX1 G43316 (.I(W14572), .ZN(O3793));
  INVX1 G43317 (.I(W18703), .ZN(W26553));
  INVX1 G43318 (.I(W11590), .ZN(W26552));
  INVX1 G43319 (.I(W6360), .ZN(W26551));
  INVX1 G43320 (.I(W11492), .ZN(W26560));
  INVX1 G43321 (.I(W1927), .ZN(W26547));
  INVX1 G43322 (.I(W12410), .ZN(W24203));
  INVX1 G43323 (.I(W8045), .ZN(W24204));
  INVX1 G43324 (.I(W12275), .ZN(W24206));
  INVX1 G43325 (.I(W21501), .ZN(O3790));
  INVX1 G43326 (.I(W17418), .ZN(O3789));
  INVX1 G43327 (.I(W4765), .ZN(W26540));
  INVX1 G43328 (.I(W687), .ZN(W26539));
  INVX1 G43329 (.I(W1388), .ZN(W26537));
  INVX1 G43330 (.I(W15523), .ZN(W26576));
  INVX1 G43331 (.I(W25212), .ZN(O3802));
  INVX1 G43332 (.I(W14864), .ZN(W26587));
  INVX1 G43333 (.I(W17801), .ZN(W26586));
  INVX1 G43334 (.I(W19691), .ZN(W24160));
  INVX1 G43335 (.I(W3177), .ZN(W24162));
  INVX1 G43336 (.I(W20338), .ZN(W24163));
  INVX1 G43337 (.I(W20307), .ZN(W24165));
  INVX1 G43338 (.I(W12297), .ZN(W24166));
  INVX1 G43339 (.I(W7147), .ZN(O3798));
  INVX1 G43340 (.I(I1003), .ZN(W26658));
  INVX1 G43341 (.I(W25876), .ZN(W26573));
  INVX1 G43342 (.I(W13948), .ZN(O2990));
  INVX1 G43343 (.I(W3147), .ZN(O2991));
  INVX1 G43344 (.I(W1025), .ZN(W26569));
  INVX1 G43345 (.I(W20610), .ZN(W24179));
  INVX1 G43346 (.I(W2956), .ZN(W26564));
  INVX1 G43347 (.I(W3180), .ZN(W24183));
  INVX1 G43348 (.I(W10449), .ZN(O2996));
  INVX1 G43349 (.I(W18662), .ZN(O2997));
  INVX1 G43350 (.I(W13817), .ZN(W23997));
  INVX1 G43351 (.I(W1766), .ZN(O2940));
  INVX1 G43352 (.I(W3279), .ZN(W23986));
  INVX1 G43353 (.I(W13085), .ZN(O3856));
  INVX1 G43354 (.I(I1764), .ZN(O2941));
  INVX1 G43355 (.I(W12116), .ZN(W23990));
  INVX1 G43356 (.I(W7987), .ZN(O2943));
  INVX1 G43357 (.I(W2971), .ZN(O3854));
  INVX1 G43358 (.I(W1431), .ZN(O3853));
  INVX1 G43359 (.I(I340), .ZN(W23994));
  INVX1 G43360 (.I(W2107), .ZN(W26734));
  INVX1 G43361 (.I(W14268), .ZN(W23983));
  INVX1 G43362 (.I(W19077), .ZN(W24004));
  INVX1 G43363 (.I(W5474), .ZN(W26726));
  INVX1 G43364 (.I(W22032), .ZN(W24007));
  INVX1 G43365 (.I(I580), .ZN(O3846));
  INVX1 G43366 (.I(W18872), .ZN(W24010));
  INVX1 G43367 (.I(W19405), .ZN(W24015));
  INVX1 G43368 (.I(W1470), .ZN(W26720));
  INVX1 G43369 (.I(I1280), .ZN(W24018));
  INVX1 G43370 (.I(W8909), .ZN(W24024));
  INVX1 G43371 (.I(W25255), .ZN(W26759));
  INVX1 G43372 (.I(W2170), .ZN(O2932));
  INVX1 G43373 (.I(W9157), .ZN(W23964));
  INVX1 G43374 (.I(W8641), .ZN(W26766));
  INVX1 G43375 (.I(W5276), .ZN(O3862));
  INVX1 G43376 (.I(W15217), .ZN(W23967));
  INVX1 G43377 (.I(W20077), .ZN(O2934));
  INVX1 G43378 (.I(W5481), .ZN(O3860));
  INVX1 G43379 (.I(W12459), .ZN(W23970));
  INVX1 G43380 (.I(W11337), .ZN(W26760));
  INVX1 G43381 (.I(I60), .ZN(W26714));
  INVX1 G43382 (.I(W8265), .ZN(W23972));
  INVX1 G43383 (.I(W23071), .ZN(W23974));
  INVX1 G43384 (.I(W3297), .ZN(W26756));
  INVX1 G43385 (.I(W14391), .ZN(W26755));
  INVX1 G43386 (.I(W8482), .ZN(W23976));
  INVX1 G43387 (.I(W17337), .ZN(W23978));
  INVX1 G43388 (.I(W11638), .ZN(O2938));
  INVX1 G43389 (.I(W21023), .ZN(O3858));
  INVX1 G43390 (.I(W26428), .ZN(W26748));
  INVX1 G43391 (.I(I662), .ZN(O2963));
  INVX1 G43392 (.I(W22160), .ZN(W24049));
  INVX1 G43393 (.I(W13302), .ZN(W24050));
  INVX1 G43394 (.I(W3125), .ZN(O3832));
  INVX1 G43395 (.I(W24172), .ZN(W26681));
  INVX1 G43396 (.I(W24513), .ZN(W26680));
  INVX1 G43397 (.I(W16773), .ZN(W24055));
  INVX1 G43398 (.I(W4523), .ZN(W24062));
  INVX1 G43399 (.I(W13235), .ZN(W24064));
  INVX1 G43400 (.I(W14352), .ZN(O3828));
  INVX1 G43401 (.I(W15846), .ZN(W26685));
  INVX1 G43402 (.I(W311), .ZN(W24069));
  INVX1 G43403 (.I(W8903), .ZN(W26668));
  INVX1 G43404 (.I(W10844), .ZN(O3825));
  INVX1 G43405 (.I(W4986), .ZN(W24073));
  INVX1 G43406 (.I(W9911), .ZN(W26663));
  INVX1 G43407 (.I(W9781), .ZN(W24076));
  INVX1 G43408 (.I(W12334), .ZN(W26661));
  INVX1 G43409 (.I(W17543), .ZN(W24077));
  INVX1 G43410 (.I(W1020), .ZN(O2966));
  INVX1 G43411 (.I(W23937), .ZN(O3839));
  INVX1 G43412 (.I(W20871), .ZN(W24025));
  INVX1 G43413 (.I(W23045), .ZN(W26712));
  INVX1 G43414 (.I(W4631), .ZN(O2952));
  INVX1 G43415 (.I(W2366), .ZN(O2953));
  INVX1 G43416 (.I(W18272), .ZN(O3841));
  INVX1 G43417 (.I(W11660), .ZN(W26706));
  INVX1 G43418 (.I(W14639), .ZN(W24030));
  INVX1 G43419 (.I(W5852), .ZN(W26704));
  INVX1 G43420 (.I(W18473), .ZN(O3840));
  INVX1 G43421 (.I(W22989), .ZN(O3000));
  INVX1 G43422 (.I(W11150), .ZN(O2955));
  INVX1 G43423 (.I(W16037), .ZN(W26698));
  INVX1 G43424 (.I(W19395), .ZN(W24036));
  INVX1 G43425 (.I(W3706), .ZN(W24040));
  INVX1 G43426 (.I(W21263), .ZN(O3837));
  INVX1 G43427 (.I(W6925), .ZN(W24042));
  INVX1 G43428 (.I(W7706), .ZN(W24044));
  INVX1 G43429 (.I(I1736), .ZN(O3836));
  INVX1 G43430 (.I(W3577), .ZN(O2959));
  INVX1 G43431 (.I(W3387), .ZN(W26370));
  INVX1 G43432 (.I(W19653), .ZN(W26383));
  INVX1 G43433 (.I(W11689), .ZN(O3737));
  INVX1 G43434 (.I(W4551), .ZN(O3736));
  INVX1 G43435 (.I(W19842), .ZN(W24366));
  INVX1 G43436 (.I(W8806), .ZN(O3735));
  INVX1 G43437 (.I(W23933), .ZN(O3059));
  INVX1 G43438 (.I(W1826), .ZN(O3060));
  INVX1 G43439 (.I(W23165), .ZN(O3061));
  INVX1 G43440 (.I(W25744), .ZN(W26374));
  INVX1 G43441 (.I(W9116), .ZN(O3063));
  INVX1 G43442 (.I(W23473), .ZN(W24363));
  INVX1 G43443 (.I(W10179), .ZN(O3065));
  INVX1 G43444 (.I(W12333), .ZN(O3731));
  INVX1 G43445 (.I(W7819), .ZN(O3066));
  INVX1 G43446 (.I(W6144), .ZN(W24381));
  INVX1 G43447 (.I(W13639), .ZN(W24388));
  INVX1 G43448 (.I(W11574), .ZN(W26361));
  INVX1 G43449 (.I(W17761), .ZN(W26360));
  INVX1 G43450 (.I(I1122), .ZN(O3069));
  INVX1 G43451 (.I(W999), .ZN(W26357));
  INVX1 G43452 (.I(W1184), .ZN(W26405));
  INVX1 G43453 (.I(I1946), .ZN(W26418));
  INVX1 G43454 (.I(W2544), .ZN(O3747));
  INVX1 G43455 (.I(W5703), .ZN(W24326));
  INVX1 G43456 (.I(W20004), .ZN(W26413));
  INVX1 G43457 (.I(W25128), .ZN(O3746));
  INVX1 G43458 (.I(W12972), .ZN(O3045));
  INVX1 G43459 (.I(W24051), .ZN(O3046));
  INVX1 G43460 (.I(W12056), .ZN(W24338));
  INVX1 G43461 (.I(W15948), .ZN(O3047));
  INVX1 G43462 (.I(W18294), .ZN(W26356));
  INVX1 G43463 (.I(W3657), .ZN(O3049));
  INVX1 G43464 (.I(W10976), .ZN(O3050));
  INVX1 G43465 (.I(W7694), .ZN(O3051));
  INVX1 G43466 (.I(W19310), .ZN(O3052));
  INVX1 G43467 (.I(W12284), .ZN(O3053));
  INVX1 G43468 (.I(W14918), .ZN(O3744));
  INVX1 G43469 (.I(W17665), .ZN(W26394));
  INVX1 G43470 (.I(W5238), .ZN(W24352));
  INVX1 G43471 (.I(W23621), .ZN(O3054));
  INVX1 G43472 (.I(W8435), .ZN(O3081));
  INVX1 G43473 (.I(I1508), .ZN(W24418));
  INVX1 G43474 (.I(I1478), .ZN(O3079));
  INVX1 G43475 (.I(W22793), .ZN(O3717));
  INVX1 G43476 (.I(W9400), .ZN(O3716));
  INVX1 G43477 (.I(I198), .ZN(W24421));
  INVX1 G43478 (.I(W12505), .ZN(O3713));
  INVX1 G43479 (.I(W2061), .ZN(W26318));
  INVX1 G43480 (.I(W1861), .ZN(W26315));
  INVX1 G43481 (.I(W2073), .ZN(W24427));
  INVX1 G43482 (.I(W6261), .ZN(O3077));
  INVX1 G43483 (.I(W19155), .ZN(W24431));
  INVX1 G43484 (.I(W9731), .ZN(W26308));
  INVX1 G43485 (.I(W4687), .ZN(W26307));
  INVX1 G43486 (.I(W13473), .ZN(W26306));
  INVX1 G43487 (.I(W11006), .ZN(W24433));
  INVX1 G43488 (.I(W6480), .ZN(O3709));
  INVX1 G43489 (.I(W22558), .ZN(W24447));
  INVX1 G43490 (.I(W3217), .ZN(W24448));
  INVX1 G43491 (.I(W20763), .ZN(O3086));
  INVX1 G43492 (.I(W7562), .ZN(W26344));
  INVX1 G43493 (.I(W17745), .ZN(W24393));
  INVX1 G43494 (.I(W12831), .ZN(W26353));
  INVX1 G43495 (.I(W15032), .ZN(O3072));
  INVX1 G43496 (.I(W21767), .ZN(W24399));
  INVX1 G43497 (.I(W22311), .ZN(W24401));
  INVX1 G43498 (.I(W22943), .ZN(W26348));
  INVX1 G43499 (.I(W12090), .ZN(O3073));
  INVX1 G43500 (.I(W1066), .ZN(O3074));
  INVX1 G43501 (.I(I1308), .ZN(W26345));
  INVX1 G43502 (.I(W20355), .ZN(W26419));
  INVX1 G43503 (.I(W13062), .ZN(W26340));
  INVX1 G43504 (.I(I926), .ZN(W26339));
  INVX1 G43505 (.I(W10377), .ZN(W26338));
  INVX1 G43506 (.I(W23725), .ZN(O3724));
  INVX1 G43507 (.I(W8012), .ZN(W26334));
  INVX1 G43508 (.I(W4853), .ZN(W24411));
  INVX1 G43509 (.I(W12530), .ZN(W24412));
  INVX1 G43510 (.I(W2849), .ZN(W26331));
  INVX1 G43511 (.I(W9939), .ZN(O3721));
  INVX1 G43512 (.I(I1908), .ZN(O3772));
  INVX1 G43513 (.I(W17759), .ZN(W24238));
  INVX1 G43514 (.I(W11551), .ZN(W26502));
  INVX1 G43515 (.I(W3227), .ZN(W24241));
  INVX1 G43516 (.I(W7910), .ZN(O3014));
  INVX1 G43517 (.I(W11869), .ZN(W24246));
  INVX1 G43518 (.I(W12905), .ZN(W26493));
  INVX1 G43519 (.I(W23256), .ZN(W26491));
  INVX1 G43520 (.I(W26385), .ZN(W26490));
  INVX1 G43521 (.I(W22099), .ZN(W24252));
  INVX1 G43522 (.I(W267), .ZN(W26505));
  INVX1 G43523 (.I(W421), .ZN(W26486));
  INVX1 G43524 (.I(W11066), .ZN(O3020));
  INVX1 G43525 (.I(W4374), .ZN(W26484));
  INVX1 G43526 (.I(W271), .ZN(W24258));
  INVX1 G43527 (.I(W18873), .ZN(W26482));
  INVX1 G43528 (.I(W25475), .ZN(O3771));
  INVX1 G43529 (.I(W8133), .ZN(O3770));
  INVX1 G43530 (.I(W15764), .ZN(O3768));
  INVX1 G43531 (.I(W22947), .ZN(W26476));
  INVX1 G43532 (.I(W1745), .ZN(O3781));
  INVX1 G43533 (.I(W14548), .ZN(O3787));
  INVX1 G43534 (.I(W21590), .ZN(O3002));
  INVX1 G43535 (.I(W3792), .ZN(O3786));
  INVX1 G43536 (.I(W9588), .ZN(O3004));
  INVX1 G43537 (.I(I1958), .ZN(O3005));
  INVX1 G43538 (.I(W3450), .ZN(O3783));
  INVX1 G43539 (.I(W9865), .ZN(W24220));
  INVX1 G43540 (.I(W23684), .ZN(W26523));
  INVX1 G43541 (.I(W12561), .ZN(W24221));
  INVX1 G43542 (.I(W21713), .ZN(W26475));
  INVX1 G43543 (.I(W14211), .ZN(W26518));
  INVX1 G43544 (.I(W2143), .ZN(O3007));
  INVX1 G43545 (.I(W1888), .ZN(W26515));
  INVX1 G43546 (.I(W10927), .ZN(W24226));
  INVX1 G43547 (.I(W16069), .ZN(W26513));
  INVX1 G43548 (.I(W2913), .ZN(W26512));
  INVX1 G43549 (.I(W6875), .ZN(W24231));
  INVX1 G43550 (.I(W12981), .ZN(W24232));
  INVX1 G43551 (.I(W10604), .ZN(W26507));
  INVX1 G43552 (.I(W4301), .ZN(W24307));
  INVX1 G43553 (.I(W6965), .ZN(W26448));
  INVX1 G43554 (.I(W13513), .ZN(O3036));
  INVX1 G43555 (.I(W4405), .ZN(W26445));
  INVX1 G43556 (.I(W26344), .ZN(W26444));
  INVX1 G43557 (.I(W13355), .ZN(W26442));
  INVX1 G43558 (.I(W1899), .ZN(O3038));
  INVX1 G43559 (.I(W10033), .ZN(W26440));
  INVX1 G43560 (.I(W13702), .ZN(W26439));
  INVX1 G43561 (.I(W25565), .ZN(O3756));
  INVX1 G43562 (.I(W10652), .ZN(W24295));
  INVX1 G43563 (.I(W22), .ZN(W26435));
  INVX1 G43564 (.I(W15916), .ZN(W26433));
  INVX1 G43565 (.I(W15803), .ZN(W24311));
  INVX1 G43566 (.I(W12560), .ZN(O3042));
  INVX1 G43567 (.I(I814), .ZN(W24313));
  INVX1 G43568 (.I(W16268), .ZN(W24314));
  INVX1 G43569 (.I(W15039), .ZN(O3751));
  INVX1 G43570 (.I(W6284), .ZN(W24320));
  INVX1 G43571 (.I(W18799), .ZN(W24322));
  INVX1 G43572 (.I(W8879), .ZN(W26462));
  INVX1 G43573 (.I(W18843), .ZN(W26474));
  INVX1 G43574 (.I(W23807), .ZN(W24261));
  INVX1 G43575 (.I(W21031), .ZN(W26470));
  INVX1 G43576 (.I(W19413), .ZN(W24268));
  INVX1 G43577 (.I(W12341), .ZN(O3024));
  INVX1 G43578 (.I(W9174), .ZN(O3026));
  INVX1 G43579 (.I(W23390), .ZN(O3027));
  INVX1 G43580 (.I(W11293), .ZN(O3028));
  INVX1 G43581 (.I(W9011), .ZN(W24282));
  INVX1 G43582 (.I(W5050), .ZN(W23959));
  INVX1 G43583 (.I(W12876), .ZN(W24285));
  INVX1 G43584 (.I(W23210), .ZN(W26459));
  INVX1 G43585 (.I(W1013), .ZN(W26458));
  INVX1 G43586 (.I(W7798), .ZN(O3760));
  INVX1 G43587 (.I(W20465), .ZN(O3033));
  INVX1 G43588 (.I(I1438), .ZN(O3034));
  INVX1 G43589 (.I(W14646), .ZN(W24293));
  INVX1 G43590 (.I(W9302), .ZN(O3759));
  INVX1 G43591 (.I(W2066), .ZN(O3035));
  INVX1 G43592 (.I(W582), .ZN(W27105));
  INVX1 G43593 (.I(W26383), .ZN(W27121));
  INVX1 G43594 (.I(W17431), .ZN(O3992));
  INVX1 G43595 (.I(W14616), .ZN(W27118));
  INVX1 G43596 (.I(W11852), .ZN(W23609));
  INVX1 G43597 (.I(W12265), .ZN(W23611));
  INVX1 G43598 (.I(W11893), .ZN(W23614));
  INVX1 G43599 (.I(W16906), .ZN(O3988));
  INVX1 G43600 (.I(W2449), .ZN(W27111));
  INVX1 G43601 (.I(W21803), .ZN(O2831));
  INVX1 G43602 (.I(W12641), .ZN(O3984));
  INVX1 G43603 (.I(W15859), .ZN(W23602));
  INVX1 G43604 (.I(W16182), .ZN(O2832));
  INVX1 G43605 (.I(W5956), .ZN(W23625));
  INVX1 G43606 (.I(W14972), .ZN(W27100));
  INVX1 G43607 (.I(W7515), .ZN(O3982));
  INVX1 G43608 (.I(W7811), .ZN(O3981));
  INVX1 G43609 (.I(W20282), .ZN(W23636));
  INVX1 G43610 (.I(W19582), .ZN(W27095));
  INVX1 G43611 (.I(W12071), .ZN(W23638));
  INVX1 G43612 (.I(W7551), .ZN(W27091));
  INVX1 G43613 (.I(W18644), .ZN(W23589));
  INVX1 G43614 (.I(W9528), .ZN(W23579));
  INVX1 G43615 (.I(W20365), .ZN(O4000));
  INVX1 G43616 (.I(W4751), .ZN(O3999));
  INVX1 G43617 (.I(W7109), .ZN(O3997));
  INVX1 G43618 (.I(I457), .ZN(W23581));
  INVX1 G43619 (.I(W14691), .ZN(O2819));
  INVX1 G43620 (.I(W3334), .ZN(W23583));
  INVX1 G43621 (.I(W20569), .ZN(W23586));
  INVX1 G43622 (.I(W781), .ZN(O2821));
  INVX1 G43623 (.I(W4016), .ZN(O2839));
  INVX1 G43624 (.I(I1626), .ZN(W23590));
  INVX1 G43625 (.I(W3579), .ZN(W23591));
  INVX1 G43626 (.I(W11318), .ZN(W27134));
  INVX1 G43627 (.I(W22902), .ZN(O2823));
  INVX1 G43628 (.I(W5573), .ZN(W27131));
  INVX1 G43629 (.I(W8407), .ZN(W23597));
  INVX1 G43630 (.I(W20511), .ZN(W27128));
  INVX1 G43631 (.I(W14214), .ZN(W27126));
  INVX1 G43632 (.I(W23304), .ZN(O2825));
  INVX1 G43633 (.I(W22757), .ZN(W23684));
  INVX1 G43634 (.I(W16458), .ZN(W23677));
  INVX1 G43635 (.I(I704), .ZN(W27046));
  INVX1 G43636 (.I(W12307), .ZN(W23679));
  INVX1 G43637 (.I(W15825), .ZN(W27044));
  INVX1 G43638 (.I(W16810), .ZN(O3967));
  INVX1 G43639 (.I(W20683), .ZN(O3965));
  INVX1 G43640 (.I(W6810), .ZN(W27039));
  INVX1 G43641 (.I(W411), .ZN(W23682));
  INVX1 G43642 (.I(W5044), .ZN(W23683));
  INVX1 G43643 (.I(W836), .ZN(O2848));
  INVX1 G43644 (.I(W10736), .ZN(O2850));
  INVX1 G43645 (.I(W19568), .ZN(W27032));
  INVX1 G43646 (.I(W5232), .ZN(O3964));
  INVX1 G43647 (.I(W2550), .ZN(W23691));
  INVX1 G43648 (.I(W7974), .ZN(W27028));
  INVX1 G43649 (.I(W7180), .ZN(W23693));
  INVX1 G43650 (.I(W14367), .ZN(W27025));
  INVX1 G43651 (.I(W11552), .ZN(O2852));
  INVX1 G43652 (.I(W7328), .ZN(O2854));
  INVX1 G43653 (.I(W23359), .ZN(W27065));
  INVX1 G43654 (.I(W11622), .ZN(W27083));
  INVX1 G43655 (.I(W12100), .ZN(O3979));
  INVX1 G43656 (.I(W26739), .ZN(W27081));
  INVX1 G43657 (.I(W12395), .ZN(O3976));
  INVX1 G43658 (.I(W4487), .ZN(W27074));
  INVX1 G43659 (.I(W19102), .ZN(O3975));
  INVX1 G43660 (.I(W10696), .ZN(W23657));
  INVX1 G43661 (.I(W1022), .ZN(W27071));
  INVX1 G43662 (.I(W11514), .ZN(W23658));
  INVX1 G43663 (.I(W272), .ZN(W27149));
  INVX1 G43664 (.I(W8818), .ZN(W27064));
  INVX1 G43665 (.I(W15905), .ZN(W27063));
  INVX1 G43666 (.I(W21144), .ZN(W23665));
  INVX1 G43667 (.I(W11447), .ZN(W23667));
  INVX1 G43668 (.I(W602), .ZN(W27057));
  INVX1 G43669 (.I(W1515), .ZN(W23669));
  INVX1 G43670 (.I(W26074), .ZN(W27055));
  INVX1 G43671 (.I(W10021), .ZN(O2846));
  INVX1 G43672 (.I(W10821), .ZN(W23675));
  INVX1 G43673 (.I(W26892), .ZN(O4029));
  INVX1 G43674 (.I(W21719), .ZN(O2797));
  INVX1 G43675 (.I(W16973), .ZN(W23498));
  INVX1 G43676 (.I(W6764), .ZN(O2798));
  INVX1 G43677 (.I(W14270), .ZN(W23503));
  INVX1 G43678 (.I(W13422), .ZN(W27238));
  INVX1 G43679 (.I(W3944), .ZN(O4030));
  INVX1 G43680 (.I(W24016), .ZN(W27235));
  INVX1 G43681 (.I(W18392), .ZN(O2800));
  INVX1 G43682 (.I(W10754), .ZN(W23506));
  INVX1 G43683 (.I(W25833), .ZN(W27247));
  INVX1 G43684 (.I(W468), .ZN(W27229));
  INVX1 G43685 (.I(W21229), .ZN(O2801));
  INVX1 G43686 (.I(W7651), .ZN(W27224));
  INVX1 G43687 (.I(I1968), .ZN(W23516));
  INVX1 G43688 (.I(W21534), .ZN(W27220));
  INVX1 G43689 (.I(W13721), .ZN(O2805));
  INVX1 G43690 (.I(W26524), .ZN(O4026));
  INVX1 G43691 (.I(I661), .ZN(W27213));
  INVX1 G43692 (.I(W7645), .ZN(W23526));
  INVX1 G43693 (.I(W3597), .ZN(O2787));
  INVX1 G43694 (.I(W6039), .ZN(O4047));
  INVX1 G43695 (.I(W8123), .ZN(W23468));
  INVX1 G43696 (.I(W16021), .ZN(W23469));
  INVX1 G43697 (.I(W6242), .ZN(W27269));
  INVX1 G43698 (.I(W4930), .ZN(W27267));
  INVX1 G43699 (.I(W17777), .ZN(W23472));
  INVX1 G43700 (.I(W51), .ZN(W23473));
  INVX1 G43701 (.I(W9897), .ZN(O2786));
  INVX1 G43702 (.I(W6411), .ZN(W27261));
  INVX1 G43703 (.I(W24299), .ZN(W27210));
  INVX1 G43704 (.I(W11699), .ZN(O4040));
  INVX1 G43705 (.I(W21161), .ZN(O2788));
  INVX1 G43706 (.I(W6501), .ZN(O2791));
  INVX1 G43707 (.I(W22074), .ZN(O4039));
  INVX1 G43708 (.I(W15712), .ZN(W23484));
  INVX1 G43709 (.I(W4837), .ZN(W23486));
  INVX1 G43710 (.I(W7126), .ZN(O2793));
  INVX1 G43711 (.I(W18916), .ZN(O4037));
  INVX1 G43712 (.I(W11043), .ZN(W27248));
  INVX1 G43713 (.I(W21654), .ZN(W23568));
  INVX1 G43714 (.I(W23294), .ZN(W27173));
  INVX1 G43715 (.I(W9214), .ZN(O2814));
  INVX1 G43716 (.I(W13644), .ZN(W23563));
  INVX1 G43717 (.I(W20018), .ZN(O4008));
  INVX1 G43718 (.I(W18805), .ZN(W27168));
  INVX1 G43719 (.I(I81), .ZN(W23565));
  INVX1 G43720 (.I(W14967), .ZN(W27164));
  INVX1 G43721 (.I(W13251), .ZN(O4007));
  INVX1 G43722 (.I(W25666), .ZN(W27162));
  INVX1 G43723 (.I(W14667), .ZN(W23558));
  INVX1 G43724 (.I(W15204), .ZN(W27160));
  INVX1 G43725 (.I(W25853), .ZN(O4006));
  INVX1 G43726 (.I(W1781), .ZN(W23571));
  INVX1 G43727 (.I(W21524), .ZN(W27156));
  INVX1 G43728 (.I(W5036), .ZN(W23572));
  INVX1 G43729 (.I(W4372), .ZN(O4003));
  INVX1 G43730 (.I(W12385), .ZN(W23573));
  INVX1 G43731 (.I(W15270), .ZN(W23576));
  INVX1 G43732 (.I(W15560), .ZN(W23578));
  INVX1 G43733 (.I(W13548), .ZN(W23537));
  INVX1 G43734 (.I(W24468), .ZN(O4023));
  INVX1 G43735 (.I(W936), .ZN(W27205));
  INVX1 G43736 (.I(I285), .ZN(W27204));
  INVX1 G43737 (.I(W9299), .ZN(W23531));
  INVX1 G43738 (.I(W18176), .ZN(O4022));
  INVX1 G43739 (.I(W11110), .ZN(W27199));
  INVX1 G43740 (.I(W19381), .ZN(W27198));
  INVX1 G43741 (.I(W22028), .ZN(W23533));
  INVX1 G43742 (.I(W11464), .ZN(W27193));
  INVX1 G43743 (.I(W14313), .ZN(O2855));
  INVX1 G43744 (.I(W21354), .ZN(O4016));
  INVX1 G43745 (.I(W1506), .ZN(O2811));
  INVX1 G43746 (.I(W12143), .ZN(W27186));
  INVX1 G43747 (.I(W21920), .ZN(W23545));
  INVX1 G43748 (.I(W26731), .ZN(W27183));
  INVX1 G43749 (.I(W20652), .ZN(O2812));
  INVX1 G43750 (.I(W15753), .ZN(W23554));
  INVX1 G43751 (.I(W3486), .ZN(W23556));
  INVX1 G43752 (.I(I618), .ZN(W23557));
  INVX1 G43753 (.I(W9428), .ZN(O2906));
  INVX1 G43754 (.I(W7311), .ZN(W23840));
  INVX1 G43755 (.I(W24779), .ZN(W26875));
  INVX1 G43756 (.I(W20298), .ZN(W23843));
  INVX1 G43757 (.I(W17739), .ZN(W26872));
  INVX1 G43758 (.I(W1844), .ZN(W26871));
  INVX1 G43759 (.I(W14318), .ZN(W23848));
  INVX1 G43760 (.I(I51), .ZN(W26865));
  INVX1 G43761 (.I(W6051), .ZN(O2901));
  INVX1 G43762 (.I(W2746), .ZN(O2905));
  INVX1 G43763 (.I(W17968), .ZN(O3895));
  INVX1 G43764 (.I(W23095), .ZN(W23839));
  INVX1 G43765 (.I(W957), .ZN(W26856));
  INVX1 G43766 (.I(W16157), .ZN(W26855));
  INVX1 G43767 (.I(W3196), .ZN(W23862));
  INVX1 G43768 (.I(W2133), .ZN(W23864));
  INVX1 G43769 (.I(W21921), .ZN(W26851));
  INVX1 G43770 (.I(W21907), .ZN(O3892));
  INVX1 G43771 (.I(W7034), .ZN(W23865));
  INVX1 G43772 (.I(I1875), .ZN(O2908));
  INVX1 G43773 (.I(W22287), .ZN(W26846));
  INVX1 G43774 (.I(W9629), .ZN(W26896));
  INVX1 G43775 (.I(W936), .ZN(O3916));
  INVX1 G43776 (.I(W15153), .ZN(W23804));
  INVX1 G43777 (.I(W17348), .ZN(W23807));
  INVX1 G43778 (.I(W7293), .ZN(W26905));
  INVX1 G43779 (.I(W10820), .ZN(W23809));
  INVX1 G43780 (.I(W7151), .ZN(O2887));
  INVX1 G43781 (.I(W20365), .ZN(W23820));
  INVX1 G43782 (.I(W1412), .ZN(O2890));
  INVX1 G43783 (.I(W21313), .ZN(W26897));
  INVX1 G43784 (.I(W13827), .ZN(O3891));
  INVX1 G43785 (.I(W4407), .ZN(O3911));
  INVX1 G43786 (.I(W2920), .ZN(W26892));
  INVX1 G43787 (.I(W12635), .ZN(W26889));
  INVX1 G43788 (.I(W114), .ZN(O3908));
  INVX1 G43789 (.I(W24526), .ZN(O3905));
  INVX1 G43790 (.I(W17516), .ZN(O2893));
  INVX1 G43791 (.I(W21748), .ZN(W23832));
  INVX1 G43792 (.I(W9823), .ZN(O3902));
  INVX1 G43793 (.I(W11320), .ZN(W26880));
  INVX1 G43794 (.I(W19508), .ZN(W23934));
  INVX1 G43795 (.I(W2387), .ZN(W23913));
  INVX1 G43796 (.I(W17994), .ZN(O2919));
  INVX1 G43797 (.I(W17919), .ZN(W23916));
  INVX1 G43798 (.I(W12100), .ZN(W23919));
  INVX1 G43799 (.I(W14373), .ZN(O2923));
  INVX1 G43800 (.I(W22175), .ZN(O3875));
  INVX1 G43801 (.I(W2292), .ZN(O3874));
  INVX1 G43802 (.I(W13524), .ZN(W23925));
  INVX1 G43803 (.I(W19662), .ZN(W23929));
  INVX1 G43804 (.I(W9123), .ZN(W23912));
  INVX1 G43805 (.I(W3359), .ZN(W26791));
  INVX1 G43806 (.I(I978), .ZN(W26790));
  INVX1 G43807 (.I(W14523), .ZN(W26789));
  INVX1 G43808 (.I(W8511), .ZN(O2926));
  INVX1 G43809 (.I(W3200), .ZN(O3868));
  INVX1 G43810 (.I(W14915), .ZN(W23947));
  INVX1 G43811 (.I(W12990), .ZN(O2930));
  INVX1 G43812 (.I(W4966), .ZN(W26773));
  INVX1 G43813 (.I(W7769), .ZN(W23957));
  INVX1 G43814 (.I(W80), .ZN(O2914));
  INVX1 G43815 (.I(W5232), .ZN(O2910));
  INVX1 G43816 (.I(W5280), .ZN(W26843));
  INVX1 G43817 (.I(W1962), .ZN(W26842));
  INVX1 G43818 (.I(I1418), .ZN(O2911));
  INVX1 G43819 (.I(W16974), .ZN(W23871));
  INVX1 G43820 (.I(W12804), .ZN(O2913));
  INVX1 G43821 (.I(W17986), .ZN(W23879));
  INVX1 G43822 (.I(W17594), .ZN(O3888));
  INVX1 G43823 (.I(W18379), .ZN(W23882));
  INVX1 G43824 (.I(W383), .ZN(W23803));
  INVX1 G43825 (.I(W19159), .ZN(O2916));
  INVX1 G43826 (.I(W19626), .ZN(W26826));
  INVX1 G43827 (.I(W3840), .ZN(W23891));
  INVX1 G43828 (.I(W21099), .ZN(W23892));
  INVX1 G43829 (.I(W20450), .ZN(W23896));
  INVX1 G43830 (.I(I797), .ZN(W23901));
  INVX1 G43831 (.I(W23341), .ZN(W23905));
  INVX1 G43832 (.I(W17904), .ZN(W23908));
  INVX1 G43833 (.I(W6777), .ZN(W23911));
  INVX1 G43834 (.I(W2463), .ZN(W26982));
  INVX1 G43835 (.I(I601), .ZN(O2861));
  INVX1 G43836 (.I(W14579), .ZN(O2862));
  INVX1 G43837 (.I(W17059), .ZN(O2863));
  INVX1 G43838 (.I(W22711), .ZN(W23737));
  INVX1 G43839 (.I(W19924), .ZN(O3952));
  INVX1 G43840 (.I(W23061), .ZN(W26988));
  INVX1 G43841 (.I(W5630), .ZN(O3951));
  INVX1 G43842 (.I(W5224), .ZN(W26985));
  INVX1 G43843 (.I(W11780), .ZN(W23740));
  INVX1 G43844 (.I(W1548), .ZN(W23730));
  INVX1 G43845 (.I(W13795), .ZN(W26981));
  INVX1 G43846 (.I(W11689), .ZN(W23743));
  INVX1 G43847 (.I(W21742), .ZN(W26979));
  INVX1 G43848 (.I(W17548), .ZN(W23744));
  INVX1 G43849 (.I(W3490), .ZN(W26976));
  INVX1 G43850 (.I(W17979), .ZN(O3949));
  INVX1 G43851 (.I(W6069), .ZN(W23749));
  INVX1 G43852 (.I(W16589), .ZN(W23751));
  INVX1 G43853 (.I(W10454), .ZN(W23753));
  INVX1 G43854 (.I(W5671), .ZN(W23714));
  INVX1 G43855 (.I(W22853), .ZN(W27017));
  INVX1 G43856 (.I(W7224), .ZN(W23706));
  INVX1 G43857 (.I(W20620), .ZN(W27015));
  INVX1 G43858 (.I(W9033), .ZN(W23708));
  INVX1 G43859 (.I(W24997), .ZN(W27011));
  INVX1 G43860 (.I(W21811), .ZN(O2857));
  INVX1 G43861 (.I(W16540), .ZN(W27009));
  INVX1 G43862 (.I(W11674), .ZN(W27008));
  INVX1 G43863 (.I(W6010), .ZN(W23713));
  INVX1 G43864 (.I(W6526), .ZN(O3946));
  INVX1 G43865 (.I(W13158), .ZN(W23715));
  INVX1 G43866 (.I(W6392), .ZN(W27003));
  INVX1 G43867 (.I(I1824), .ZN(W27002));
  INVX1 G43868 (.I(W8154), .ZN(O3957));
  INVX1 G43869 (.I(W20527), .ZN(O2859));
  INVX1 G43870 (.I(W9376), .ZN(W26998));
  INVX1 G43871 (.I(W15760), .ZN(W23725));
  INVX1 G43872 (.I(W21923), .ZN(O3954));
  INVX1 G43873 (.I(W6769), .ZN(W23728));
  INVX1 G43874 (.I(W7033), .ZN(O2880));
  INVX1 G43875 (.I(W4193), .ZN(W23782));
  INVX1 G43876 (.I(W12448), .ZN(O3929));
  INVX1 G43877 (.I(W23724), .ZN(O3928));
  INVX1 G43878 (.I(W8535), .ZN(W23784));
  INVX1 G43879 (.I(W10422), .ZN(W26933));
  INVX1 G43880 (.I(W3825), .ZN(O2878));
  INVX1 G43881 (.I(W7944), .ZN(O2879));
  INVX1 G43882 (.I(W16287), .ZN(W23788));
  INVX1 G43883 (.I(W10893), .ZN(O3925));
  INVX1 G43884 (.I(W17962), .ZN(W23781));
  INVX1 G43885 (.I(W15233), .ZN(W26926));
  INVX1 G43886 (.I(W12896), .ZN(O3923));
  INVX1 G43887 (.I(W24726), .ZN(W26924));
  INVX1 G43888 (.I(W22946), .ZN(W26923));
  INVX1 G43889 (.I(W16220), .ZN(W23791));
  INVX1 G43890 (.I(W6481), .ZN(W26919));
  INVX1 G43891 (.I(W21915), .ZN(W23794));
  INVX1 G43892 (.I(W1704), .ZN(O3918));
  INVX1 G43893 (.I(W20013), .ZN(W23801));
  INVX1 G43894 (.I(I1419), .ZN(O2871));
  INVX1 G43895 (.I(W18454), .ZN(W23754));
  INVX1 G43896 (.I(W22369), .ZN(W26965));
  INVX1 G43897 (.I(W1787), .ZN(O3944));
  INVX1 G43898 (.I(W4603), .ZN(O2869));
  INVX1 G43899 (.I(W25), .ZN(O3943));
  INVX1 G43900 (.I(W26238), .ZN(W26958));
  INVX1 G43901 (.I(W9176), .ZN(W26957));
  INVX1 G43902 (.I(W10886), .ZN(W23763));
  INVX1 G43903 (.I(W17000), .ZN(W23764));
  INVX1 G43904 (.I(W18150), .ZN(O3087));
  INVX1 G43905 (.I(W20486), .ZN(W23766));
  INVX1 G43906 (.I(W19029), .ZN(W23769));
  INVX1 G43907 (.I(W15393), .ZN(W23770));
  INVX1 G43908 (.I(W26401), .ZN(O3936));
  INVX1 G43909 (.I(W21467), .ZN(W26946));
  INVX1 G43910 (.I(W18051), .ZN(W23772));
  INVX1 G43911 (.I(W16937), .ZN(O2874));
  INVX1 G43912 (.I(W9792), .ZN(O3934));
  INVX1 G43913 (.I(W9942), .ZN(W23776));
  INVX1 G43914 (.I(W18569), .ZN(W25673));
  INVX1 G43915 (.I(W2668), .ZN(W25011));
  INVX1 G43916 (.I(W3797), .ZN(W25682));
  INVX1 G43917 (.I(W4159), .ZN(W25013));
  INVX1 G43918 (.I(W15002), .ZN(W25680));
  INVX1 G43919 (.I(W8472), .ZN(W25679));
  INVX1 G43920 (.I(W9505), .ZN(W25678));
  INVX1 G43921 (.I(W4265), .ZN(W25677));
  INVX1 G43922 (.I(W8968), .ZN(W25676));
  INVX1 G43923 (.I(W20148), .ZN(O3267));
  INVX1 G43924 (.I(W4458), .ZN(W25674));
  INVX1 G43925 (.I(W20290), .ZN(W25685));
  INVX1 G43926 (.I(W13552), .ZN(O3269));
  INVX1 G43927 (.I(W10889), .ZN(W25021));
  INVX1 G43928 (.I(W16723), .ZN(W25023));
  INVX1 G43929 (.I(W19428), .ZN(W25666));
  INVX1 G43930 (.I(W11478), .ZN(O3488));
  INVX1 G43931 (.I(W11111), .ZN(O3271));
  INVX1 G43932 (.I(W19966), .ZN(O3486));
  INVX1 G43933 (.I(W10558), .ZN(W25032));
  INVX1 G43934 (.I(W7538), .ZN(O3484));
  INVX1 G43935 (.I(W6235), .ZN(O3497));
  INVX1 G43936 (.I(W4450), .ZN(O3502));
  INVX1 G43937 (.I(W6872), .ZN(W24985));
  INVX1 G43938 (.I(W10034), .ZN(W24988));
  INVX1 G43939 (.I(W24158), .ZN(W25708));
  INVX1 G43940 (.I(W16101), .ZN(W24989));
  INVX1 G43941 (.I(I1217), .ZN(W24990));
  INVX1 G43942 (.I(W3187), .ZN(W24994));
  INVX1 G43943 (.I(W25630), .ZN(O3498));
  INVX1 G43944 (.I(W10988), .ZN(W25702));
  INVX1 G43945 (.I(W24256), .ZN(W25654));
  INVX1 G43946 (.I(W23955), .ZN(W24995));
  INVX1 G43947 (.I(W2633), .ZN(W25695));
  INVX1 G43948 (.I(W10068), .ZN(W25004));
  INVX1 G43949 (.I(W22510), .ZN(W25692));
  INVX1 G43950 (.I(W5792), .ZN(O3494));
  INVX1 G43951 (.I(W15641), .ZN(W25689));
  INVX1 G43952 (.I(W23276), .ZN(W25688));
  INVX1 G43953 (.I(W15396), .ZN(W25008));
  INVX1 G43954 (.I(W8223), .ZN(O3493));
  INVX1 G43955 (.I(W9168), .ZN(W25610));
  INVX1 G43956 (.I(W18158), .ZN(W25066));
  INVX1 G43957 (.I(W24889), .ZN(W25070));
  INVX1 G43958 (.I(W13284), .ZN(W25618));
  INVX1 G43959 (.I(W4577), .ZN(W25617));
  INVX1 G43960 (.I(W19761), .ZN(O3286));
  INVX1 G43961 (.I(W18297), .ZN(O3471));
  INVX1 G43962 (.I(W18630), .ZN(W25073));
  INVX1 G43963 (.I(W5931), .ZN(W25074));
  INVX1 G43964 (.I(W3273), .ZN(W25078));
  INVX1 G43965 (.I(W10292), .ZN(W25623));
  INVX1 G43966 (.I(W16911), .ZN(O3289));
  INVX1 G43967 (.I(W8337), .ZN(W25608));
  INVX1 G43968 (.I(W7222), .ZN(W25081));
  INVX1 G43969 (.I(W23802), .ZN(O3467));
  INVX1 G43970 (.I(W6363), .ZN(O3291));
  INVX1 G43971 (.I(W11733), .ZN(W25602));
  INVX1 G43972 (.I(W1152), .ZN(W25086));
  INVX1 G43973 (.I(W8266), .ZN(O3292));
  INVX1 G43974 (.I(W8961), .ZN(O3293));
  INVX1 G43975 (.I(W7350), .ZN(W25639));
  INVX1 G43976 (.I(W24116), .ZN(W25653));
  INVX1 G43977 (.I(W16173), .ZN(W25652));
  INVX1 G43978 (.I(W23293), .ZN(W25651));
  INVX1 G43979 (.I(W3362), .ZN(O3274));
  INVX1 G43980 (.I(W21708), .ZN(O3483));
  INVX1 G43981 (.I(W10376), .ZN(W25646));
  INVX1 G43982 (.I(W8430), .ZN(O3481));
  INVX1 G43983 (.I(W13273), .ZN(O3277));
  INVX1 G43984 (.I(W24550), .ZN(W25049));
  INVX1 G43985 (.I(W16990), .ZN(W25715));
  INVX1 G43986 (.I(W25608), .ZN(W25638));
  INVX1 G43987 (.I(W24766), .ZN(W25052));
  INVX1 G43988 (.I(W5796), .ZN(O3477));
  INVX1 G43989 (.I(W11992), .ZN(W25055));
  INVX1 G43990 (.I(W24231), .ZN(O3280));
  INVX1 G43991 (.I(W18519), .ZN(O3282));
  INVX1 G43992 (.I(W23533), .ZN(W25060));
  INVX1 G43993 (.I(W7719), .ZN(O3474));
  INVX1 G43994 (.I(W23491), .ZN(W25624));
  INVX1 G43995 (.I(W12211), .ZN(O3240));
  INVX1 G43996 (.I(W4952), .ZN(W24900));
  INVX1 G43997 (.I(I567), .ZN(O3533));
  INVX1 G43998 (.I(W15882), .ZN(W25795));
  INVX1 G43999 (.I(W17735), .ZN(O3532));
  INVX1 G44000 (.I(W24786), .ZN(W25793));
  INVX1 G44001 (.I(W15842), .ZN(W25792));
  INVX1 G44002 (.I(W22708), .ZN(O3531));
  INVX1 G44003 (.I(W20516), .ZN(O3238));
  INVX1 G44004 (.I(W10848), .ZN(W24912));
  INVX1 G44005 (.I(W11101), .ZN(O3534));
  INVX1 G44006 (.I(W9652), .ZN(W24916));
  INVX1 G44007 (.I(W16131), .ZN(O3241));
  INVX1 G44008 (.I(W6494), .ZN(O3526));
  INVX1 G44009 (.I(W14769), .ZN(W25779));
  INVX1 G44010 (.I(W14055), .ZN(W24921));
  INVX1 G44011 (.I(W7957), .ZN(W25776));
  INVX1 G44012 (.I(W13343), .ZN(W24924));
  INVX1 G44013 (.I(W20366), .ZN(W25774));
  INVX1 G44014 (.I(W24024), .ZN(W24926));
  INVX1 G44015 (.I(W20189), .ZN(W24875));
  INVX1 G44016 (.I(W19146), .ZN(O3544));
  INVX1 G44017 (.I(W20698), .ZN(W25831));
  INVX1 G44018 (.I(W2159), .ZN(W25829));
  INVX1 G44019 (.I(W18308), .ZN(W24870));
  INVX1 G44020 (.I(W20942), .ZN(W24872));
  INVX1 G44021 (.I(W7011), .ZN(W25826));
  INVX1 G44022 (.I(W9295), .ZN(O3542));
  INVX1 G44023 (.I(W8844), .ZN(W24873));
  INVX1 G44024 (.I(W2956), .ZN(O3224));
  INVX1 G44025 (.I(W23994), .ZN(O3244));
  INVX1 G44026 (.I(W2027), .ZN(O3226));
  INVX1 G44027 (.I(W24308), .ZN(W25818));
  INVX1 G44028 (.I(W16644), .ZN(O3538));
  INVX1 G44029 (.I(W9652), .ZN(W24883));
  INVX1 G44030 (.I(W24047), .ZN(O3537));
  INVX1 G44031 (.I(W17576), .ZN(O3229));
  INVX1 G44032 (.I(W9272), .ZN(W25806));
  INVX1 G44033 (.I(W2249), .ZN(O3233));
  INVX1 G44034 (.I(W14989), .ZN(W25800));
  INVX1 G44035 (.I(W5932), .ZN(O3508));
  INVX1 G44036 (.I(W4320), .ZN(O3512));
  INVX1 G44037 (.I(W14417), .ZN(O3255));
  INVX1 G44038 (.I(W19608), .ZN(W25740));
  INVX1 G44039 (.I(W19214), .ZN(W25739));
  INVX1 G44040 (.I(W1301), .ZN(W24960));
  INVX1 G44041 (.I(W5446), .ZN(O3510));
  INVX1 G44042 (.I(W14803), .ZN(W24963));
  INVX1 G44043 (.I(W4115), .ZN(O3258));
  INVX1 G44044 (.I(W18711), .ZN(W25730));
  INVX1 G44045 (.I(W22250), .ZN(W24952));
  INVX1 G44046 (.I(W12255), .ZN(W25727));
  INVX1 G44047 (.I(W18461), .ZN(O3259));
  INVX1 G44048 (.I(W13451), .ZN(W25723));
  INVX1 G44049 (.I(W15179), .ZN(O3506));
  INVX1 G44050 (.I(W18608), .ZN(W24975));
  INVX1 G44051 (.I(W8848), .ZN(O3504));
  INVX1 G44052 (.I(W3263), .ZN(W25718));
  INVX1 G44053 (.I(W7268), .ZN(W25717));
  INVX1 G44054 (.I(W13349), .ZN(O3503));
  INVX1 G44055 (.I(W23352), .ZN(O3517));
  INVX1 G44056 (.I(W19782), .ZN(W24930));
  INVX1 G44057 (.I(W20150), .ZN(W24932));
  INVX1 G44058 (.I(W9275), .ZN(W24934));
  INVX1 G44059 (.I(W15907), .ZN(O3246));
  INVX1 G44060 (.I(W23179), .ZN(W24937));
  INVX1 G44061 (.I(W25218), .ZN(O3522));
  INVX1 G44062 (.I(W99), .ZN(O3248));
  INVX1 G44063 (.I(W9120), .ZN(O3520));
  INVX1 G44064 (.I(W12363), .ZN(O3519));
  INVX1 G44065 (.I(W21044), .ZN(W25598));
  INVX1 G44066 (.I(W21009), .ZN(O3516));
  INVX1 G44067 (.I(W18055), .ZN(W24941));
  INVX1 G44068 (.I(W16546), .ZN(W25754));
  INVX1 G44069 (.I(W10439), .ZN(W24943));
  INVX1 G44070 (.I(W13199), .ZN(O3250));
  INVX1 G44071 (.I(W20248), .ZN(W25749));
  INVX1 G44072 (.I(W12607), .ZN(O3515));
  INVX1 G44073 (.I(W24496), .ZN(W24950));
  INVX1 G44074 (.I(W19944), .ZN(W25745));
  INVX1 G44075 (.I(W21684), .ZN(W25420));
  INVX1 G44076 (.I(W1762), .ZN(O3419));
  INVX1 G44077 (.I(W4853), .ZN(O3344));
  INVX1 G44078 (.I(W16193), .ZN(W25431));
  INVX1 G44079 (.I(W18821), .ZN(W25430));
  INVX1 G44080 (.I(W17693), .ZN(W25428));
  INVX1 G44081 (.I(W7005), .ZN(O3416));
  INVX1 G44082 (.I(W25314), .ZN(O3415));
  INVX1 G44083 (.I(W24267), .ZN(W25260));
  INVX1 G44084 (.I(W21640), .ZN(W25261));
  INVX1 G44085 (.I(W24632), .ZN(W25262));
  INVX1 G44086 (.I(W21438), .ZN(W25435));
  INVX1 G44087 (.I(W2405), .ZN(W25263));
  INVX1 G44088 (.I(W20941), .ZN(W25418));
  INVX1 G44089 (.I(W9573), .ZN(O3414));
  INVX1 G44090 (.I(W8340), .ZN(O3348));
  INVX1 G44091 (.I(W3406), .ZN(O3349));
  INVX1 G44092 (.I(W21158), .ZN(W25268));
  INVX1 G44093 (.I(W21046), .ZN(O3351));
  INVX1 G44094 (.I(W15327), .ZN(W25409));
  INVX1 G44095 (.I(W24243), .ZN(O3411));
  INVX1 G44096 (.I(W5129), .ZN(W25452));
  INVX1 G44097 (.I(W13257), .ZN(W25228));
  INVX1 G44098 (.I(I1495), .ZN(W25466));
  INVX1 G44099 (.I(W21278), .ZN(O3338));
  INVX1 G44100 (.I(W15709), .ZN(W25462));
  INVX1 G44101 (.I(W9827), .ZN(W25461));
  INVX1 G44102 (.I(W14550), .ZN(O3339));
  INVX1 G44103 (.I(W22175), .ZN(W25458));
  INVX1 G44104 (.I(W723), .ZN(W25455));
  INVX1 G44105 (.I(W6829), .ZN(W25454));
  INVX1 G44106 (.I(W8635), .ZN(O3352));
  INVX1 G44107 (.I(W17423), .ZN(O3426));
  INVX1 G44108 (.I(W24494), .ZN(W25449));
  INVX1 G44109 (.I(I873), .ZN(W25448));
  INVX1 G44110 (.I(W23596), .ZN(W25446));
  INVX1 G44111 (.I(W17737), .ZN(W25245));
  INVX1 G44112 (.I(W10376), .ZN(W25246));
  INVX1 G44113 (.I(W23431), .ZN(W25249));
  INVX1 G44114 (.I(W20104), .ZN(O3421));
  INVX1 G44115 (.I(W12441), .ZN(W25437));
  INVX1 G44116 (.I(W25283), .ZN(O3377));
  INVX1 G44117 (.I(W3611), .ZN(O3372));
  INVX1 G44118 (.I(W20655), .ZN(W25319));
  INVX1 G44119 (.I(W6734), .ZN(O3375));
  INVX1 G44120 (.I(W4529), .ZN(W25364));
  INVX1 G44121 (.I(W10176), .ZN(O3390));
  INVX1 G44122 (.I(W24795), .ZN(O3389));
  INVX1 G44123 (.I(W24131), .ZN(O3376));
  INVX1 G44124 (.I(W19887), .ZN(W25359));
  INVX1 G44125 (.I(W15631), .ZN(W25331));
  INVX1 G44126 (.I(W7044), .ZN(O3369));
  INVX1 G44127 (.I(W18883), .ZN(W25355));
  INVX1 G44128 (.I(W908), .ZN(W25334));
  INVX1 G44129 (.I(W21429), .ZN(O3379));
  INVX1 G44130 (.I(W16597), .ZN(O3385));
  INVX1 G44131 (.I(W16104), .ZN(W25349));
  INVX1 G44132 (.I(W1707), .ZN(O3383));
  INVX1 G44133 (.I(W5619), .ZN(W25341));
  INVX1 G44134 (.I(W2809), .ZN(W25345));
  INVX1 G44135 (.I(W9017), .ZN(W25344));
  INVX1 G44136 (.I(W17112), .ZN(W25286));
  INVX1 G44137 (.I(W19833), .ZN(O3354));
  INVX1 G44138 (.I(W3037), .ZN(O3355));
  INVX1 G44139 (.I(W16948), .ZN(W25403));
  INVX1 G44140 (.I(W24060), .ZN(W25277));
  INVX1 G44141 (.I(W24960), .ZN(W25281));
  INVX1 G44142 (.I(W1852), .ZN(O3409));
  INVX1 G44143 (.I(W11153), .ZN(O3408));
  INVX1 G44144 (.I(W4466), .ZN(O3407));
  INVX1 G44145 (.I(W709), .ZN(O3358));
  INVX1 G44146 (.I(W12470), .ZN(W25225));
  INVX1 G44147 (.I(W7546), .ZN(W25292));
  INVX1 G44148 (.I(W15561), .ZN(W25294));
  INVX1 G44149 (.I(W9667), .ZN(W25388));
  INVX1 G44150 (.I(W12474), .ZN(W25385));
  INVX1 G44151 (.I(W2176), .ZN(O3400));
  INVX1 G44152 (.I(W7474), .ZN(O3399));
  INVX1 G44153 (.I(W22125), .ZN(O3398));
  INVX1 G44154 (.I(W11239), .ZN(W25304));
  INVX1 G44155 (.I(W11020), .ZN(W25375));
  INVX1 G44156 (.I(W2103), .ZN(W25134));
  INVX1 G44157 (.I(W22430), .ZN(O3457));
  INVX1 G44158 (.I(W13623), .ZN(W25127));
  INVX1 G44159 (.I(W16389), .ZN(W25130));
  INVX1 G44160 (.I(W20764), .ZN(W25131));
  INVX1 G44161 (.I(W21019), .ZN(W25557));
  INVX1 G44162 (.I(W21236), .ZN(W25556));
  INVX1 G44163 (.I(W1631), .ZN(W25555));
  INVX1 G44164 (.I(W24844), .ZN(W25554));
  INVX1 G44165 (.I(W22136), .ZN(O3454));
  INVX1 G44166 (.I(W17808), .ZN(W25119));
  INVX1 G44167 (.I(W16045), .ZN(W25136));
  INVX1 G44168 (.I(W17744), .ZN(W25137));
  INVX1 G44169 (.I(W2365), .ZN(W25139));
  INVX1 G44170 (.I(W9172), .ZN(W25142));
  INVX1 G44171 (.I(W3350), .ZN(W25543));
  INVX1 G44172 (.I(W6609), .ZN(W25542));
  INVX1 G44173 (.I(I1476), .ZN(W25146));
  INVX1 G44174 (.I(W19427), .ZN(O3313));
  INVX1 G44175 (.I(W10134), .ZN(W25539));
  INVX1 G44176 (.I(W10996), .ZN(W25583));
  INVX1 G44177 (.I(W2280), .ZN(W25090));
  INVX1 G44178 (.I(W19245), .ZN(W25596));
  INVX1 G44179 (.I(W10744), .ZN(O3295));
  INVX1 G44180 (.I(W2038), .ZN(W25092));
  INVX1 G44181 (.I(W3783), .ZN(W25592));
  INVX1 G44182 (.I(W14365), .ZN(W25590));
  INVX1 G44183 (.I(W12309), .ZN(W25589));
  INVX1 G44184 (.I(W17186), .ZN(W25588));
  INVX1 G44185 (.I(W16325), .ZN(O3298));
  INVX1 G44186 (.I(W14233), .ZN(O3314));
  INVX1 G44187 (.I(W625), .ZN(O3299));
  INVX1 G44188 (.I(W17390), .ZN(W25579));
  INVX1 G44189 (.I(W1421), .ZN(W25577));
  INVX1 G44190 (.I(W12941), .ZN(O3461));
  INVX1 G44191 (.I(W1268), .ZN(O3303));
  INVX1 G44192 (.I(W16866), .ZN(W25108));
  INVX1 G44193 (.I(W12431), .ZN(W25110));
  INVX1 G44194 (.I(W9068), .ZN(W25111));
  INVX1 G44195 (.I(W17007), .ZN(W25116));
  INVX1 G44196 (.I(W9360), .ZN(O3329));
  INVX1 G44197 (.I(W1543), .ZN(W25497));
  INVX1 G44198 (.I(W12166), .ZN(W25199));
  INVX1 G44199 (.I(W21320), .ZN(W25494));
  INVX1 G44200 (.I(W17462), .ZN(W25492));
  INVX1 G44201 (.I(W9091), .ZN(W25202));
  INVX1 G44202 (.I(W7838), .ZN(W25489));
  INVX1 G44203 (.I(W12290), .ZN(W25205));
  INVX1 G44204 (.I(W25420), .ZN(O3434));
  INVX1 G44205 (.I(W5830), .ZN(W25208));
  INVX1 G44206 (.I(W21881), .ZN(O3439));
  INVX1 G44207 (.I(W3924), .ZN(W25482));
  INVX1 G44208 (.I(W1552), .ZN(W25480));
  INVX1 G44209 (.I(W16297), .ZN(W25212));
  INVX1 G44210 (.I(W11321), .ZN(W25213));
  INVX1 G44211 (.I(W11533), .ZN(W25476));
  INVX1 G44212 (.I(W14235), .ZN(W25475));
  INVX1 G44213 (.I(W18392), .ZN(W25473));
  INVX1 G44214 (.I(W19055), .ZN(W25219));
  INVX1 G44215 (.I(W22468), .ZN(O3332));
  INVX1 G44216 (.I(W24680), .ZN(O3446));
  INVX1 G44217 (.I(W2440), .ZN(W25151));
  INVX1 G44218 (.I(W18954), .ZN(W25158));
  INVX1 G44219 (.I(W13031), .ZN(W25531));
  INVX1 G44220 (.I(W8958), .ZN(W25160));
  INVX1 G44221 (.I(W11400), .ZN(O3318));
  INVX1 G44222 (.I(W13894), .ZN(W25168));
  INVX1 G44223 (.I(W8873), .ZN(O3447));
  INVX1 G44224 (.I(W24577), .ZN(W25170));
  INVX1 G44225 (.I(W13169), .ZN(W25523));
  INVX1 G44226 (.I(W178), .ZN(W24864));
  INVX1 G44227 (.I(W4937), .ZN(O3445));
  INVX1 G44228 (.I(W20137), .ZN(W25520));
  INVX1 G44229 (.I(W17493), .ZN(W25517));
  INVX1 G44230 (.I(I1709), .ZN(O3443));
  INVX1 G44231 (.I(I1445), .ZN(O3322));
  INVX1 G44232 (.I(W3691), .ZN(W25179));
  INVX1 G44233 (.I(W3597), .ZN(O3323));
  INVX1 G44234 (.I(W23769), .ZN(O3440));
  INVX1 G44235 (.I(W14338), .ZN(W25182));
  INVX1 G44236 (.I(W11677), .ZN(O3647));
  INVX1 G44237 (.I(W10725), .ZN(W24571));
  INVX1 G44238 (.I(W4251), .ZN(O3653));
  INVX1 G44239 (.I(W22130), .ZN(O3651));
  INVX1 G44240 (.I(W19852), .ZN(O3126));
  INVX1 G44241 (.I(W19565), .ZN(O3127));
  INVX1 G44242 (.I(W4228), .ZN(W24582));
  INVX1 G44243 (.I(W2083), .ZN(O3649));
  INVX1 G44244 (.I(I1977), .ZN(W24583));
  INVX1 G44245 (.I(W1690), .ZN(O3648));
  INVX1 G44246 (.I(I687), .ZN(O3128));
  INVX1 G44247 (.I(W8238), .ZN(W26154));
  INVX1 G44248 (.I(W2651), .ZN(O3129));
  INVX1 G44249 (.I(W17534), .ZN(W24594));
  INVX1 G44250 (.I(W4195), .ZN(O3132));
  INVX1 G44251 (.I(W18533), .ZN(W26131));
  INVX1 G44252 (.I(W4882), .ZN(W24598));
  INVX1 G44253 (.I(W11389), .ZN(W26129));
  INVX1 G44254 (.I(W19263), .ZN(O3134));
  INVX1 G44255 (.I(W6358), .ZN(W26127));
  INVX1 G44256 (.I(W10618), .ZN(W26126));
  INVX1 G44257 (.I(W14167), .ZN(O3116));
  INVX1 G44258 (.I(W19740), .ZN(W26180));
  INVX1 G44259 (.I(W17702), .ZN(W26179));
  INVX1 G44260 (.I(W3689), .ZN(W26178));
  INVX1 G44261 (.I(W12068), .ZN(W24549));
  INVX1 G44262 (.I(W10391), .ZN(W26175));
  INVX1 G44263 (.I(W602), .ZN(W24553));
  INVX1 G44264 (.I(W10783), .ZN(W24558));
  INVX1 G44265 (.I(W17890), .ZN(W24559));
  INVX1 G44266 (.I(W17640), .ZN(W24560));
  INVX1 G44267 (.I(W11220), .ZN(O3135));
  INVX1 G44268 (.I(W21727), .ZN(W26166));
  INVX1 G44269 (.I(W19266), .ZN(W26164));
  INVX1 G44270 (.I(W23201), .ZN(O3660));
  INVX1 G44271 (.I(W16775), .ZN(O3659));
  INVX1 G44272 (.I(W7609), .ZN(O3657));
  INVX1 G44273 (.I(W1747), .ZN(O3120));
  INVX1 G44274 (.I(W2344), .ZN(O3121));
  INVX1 G44275 (.I(W2730), .ZN(O3122));
  INVX1 G44276 (.I(W7447), .ZN(W24570));
  INVX1 G44277 (.I(W5491), .ZN(W24648));
  INVX1 G44278 (.I(W15775), .ZN(W26095));
  INVX1 G44279 (.I(W26034), .ZN(W26094));
  INVX1 G44280 (.I(W21057), .ZN(W24634));
  INVX1 G44281 (.I(W11678), .ZN(W24636));
  INVX1 G44282 (.I(W16699), .ZN(W24641));
  INVX1 G44283 (.I(W12064), .ZN(W24642));
  INVX1 G44284 (.I(W2581), .ZN(W24643));
  INVX1 G44285 (.I(W11515), .ZN(W24644));
  INVX1 G44286 (.I(W26008), .ZN(W26084));
  INVX1 G44287 (.I(W23336), .ZN(O3629));
  INVX1 G44288 (.I(W14856), .ZN(W24650));
  INVX1 G44289 (.I(W11035), .ZN(W24654));
  INVX1 G44290 (.I(W45), .ZN(W24655));
  INVX1 G44291 (.I(W25745), .ZN(O3620));
  INVX1 G44292 (.I(W10686), .ZN(W26074));
  INVX1 G44293 (.I(W4967), .ZN(W24660));
  INVX1 G44294 (.I(W3345), .ZN(W24662));
  INVX1 G44295 (.I(W23954), .ZN(W24664));
  INVX1 G44296 (.I(W4449), .ZN(W24668));
  INVX1 G44297 (.I(W22954), .ZN(W26112));
  INVX1 G44298 (.I(W20231), .ZN(O3136));
  INVX1 G44299 (.I(W9257), .ZN(O3641));
  INVX1 G44300 (.I(W3838), .ZN(W26122));
  INVX1 G44301 (.I(W11068), .ZN(W24605));
  INVX1 G44302 (.I(I687), .ZN(O3138));
  INVX1 G44303 (.I(W12480), .ZN(W26118));
  INVX1 G44304 (.I(W5427), .ZN(W24609));
  INVX1 G44305 (.I(W25935), .ZN(W26116));
  INVX1 G44306 (.I(W8024), .ZN(O3139));
  INVX1 G44307 (.I(W25350), .ZN(O3665));
  INVX1 G44308 (.I(W585), .ZN(W24626));
  INVX1 G44309 (.I(W16514), .ZN(O3147));
  INVX1 G44310 (.I(W14120), .ZN(W26105));
  INVX1 G44311 (.I(W9539), .ZN(W24629));
  INVX1 G44312 (.I(W8610), .ZN(O3148));
  INVX1 G44313 (.I(W19700), .ZN(W24632));
  INVX1 G44314 (.I(W13216), .ZN(O3631));
  INVX1 G44315 (.I(W5223), .ZN(O3630));
  INVX1 G44316 (.I(W1454), .ZN(W26097));
  INVX1 G44317 (.I(W20662), .ZN(W24487));
  INVX1 G44318 (.I(W25752), .ZN(O3697));
  INVX1 G44319 (.I(W3644), .ZN(W24478));
  INVX1 G44320 (.I(W3858), .ZN(W26260));
  INVX1 G44321 (.I(W12822), .ZN(W24480));
  INVX1 G44322 (.I(W22117), .ZN(W24482));
  INVX1 G44323 (.I(W20285), .ZN(W26256));
  INVX1 G44324 (.I(W15072), .ZN(W24484));
  INVX1 G44325 (.I(W21602), .ZN(W24485));
  INVX1 G44326 (.I(W25203), .ZN(W26253));
  INVX1 G44327 (.I(W4167), .ZN(W24473));
  INVX1 G44328 (.I(W4676), .ZN(W26251));
  INVX1 G44329 (.I(W3394), .ZN(O3097));
  INVX1 G44330 (.I(W20030), .ZN(O3694));
  INVX1 G44331 (.I(W26100), .ZN(W26247));
  INVX1 G44332 (.I(W5591), .ZN(W24492));
  INVX1 G44333 (.I(I262), .ZN(O3692));
  INVX1 G44334 (.I(W22284), .ZN(W26243));
  INVX1 G44335 (.I(W18700), .ZN(O3691));
  INVX1 G44336 (.I(W6662), .ZN(O3690));
  INVX1 G44337 (.I(I1772), .ZN(W26281));
  INVX1 G44338 (.I(W16813), .ZN(W24452));
  INVX1 G44339 (.I(W8917), .ZN(O3088));
  INVX1 G44340 (.I(W15362), .ZN(W26292));
  INVX1 G44341 (.I(W18526), .ZN(O3705));
  INVX1 G44342 (.I(W21413), .ZN(W26290));
  INVX1 G44343 (.I(W21839), .ZN(W26288));
  INVX1 G44344 (.I(W5412), .ZN(W24458));
  INVX1 G44345 (.I(W3502), .ZN(O3704));
  INVX1 G44346 (.I(W6939), .ZN(W24461));
  INVX1 G44347 (.I(W4364), .ZN(W26239));
  INVX1 G44348 (.I(W13280), .ZN(W24466));
  INVX1 G44349 (.I(W15188), .ZN(W26278));
  INVX1 G44350 (.I(W15371), .ZN(W26277));
  INVX1 G44351 (.I(W3572), .ZN(W26276));
  INVX1 G44352 (.I(W7805), .ZN(W24469));
  INVX1 G44353 (.I(W561), .ZN(W26272));
  INVX1 G44354 (.I(W17808), .ZN(W26270));
  INVX1 G44355 (.I(I964), .ZN(W26269));
  INVX1 G44356 (.I(W22573), .ZN(O3698));
  INVX1 G44357 (.I(W4607), .ZN(W24530));
  INVX1 G44358 (.I(W287), .ZN(W24523));
  INVX1 G44359 (.I(W24352), .ZN(W24524));
  INVX1 G44360 (.I(W20721), .ZN(W26206));
  INVX1 G44361 (.I(W4817), .ZN(O3108));
  INVX1 G44362 (.I(W5764), .ZN(W26204));
  INVX1 G44363 (.I(W99), .ZN(W24526));
  INVX1 G44364 (.I(W23850), .ZN(W26200));
  INVX1 G44365 (.I(W23106), .ZN(W24529));
  INVX1 G44366 (.I(W11992), .ZN(W26198));
  INVX1 G44367 (.I(W4216), .ZN(W26211));
  INVX1 G44368 (.I(W1115), .ZN(W24531));
  INVX1 G44369 (.I(W11968), .ZN(W24532));
  INVX1 G44370 (.I(W9419), .ZN(W24534));
  INVX1 G44371 (.I(W14862), .ZN(O3673));
  INVX1 G44372 (.I(W3784), .ZN(W24540));
  INVX1 G44373 (.I(W7152), .ZN(O3668));
  INVX1 G44374 (.I(W10416), .ZN(W24546));
  INVX1 G44375 (.I(W12702), .ZN(W26183));
  INVX1 G44376 (.I(W788), .ZN(O3113));
  INVX1 G44377 (.I(W5272), .ZN(O3106));
  INVX1 G44378 (.I(W2080), .ZN(W24496));
  INVX1 G44379 (.I(W15072), .ZN(W24497));
  INVX1 G44380 (.I(W22908), .ZN(O3102));
  INVX1 G44381 (.I(W12860), .ZN(W26232));
  INVX1 G44382 (.I(W19348), .ZN(O3103));
  INVX1 G44383 (.I(W9142), .ZN(W26228));
  INVX1 G44384 (.I(W1068), .ZN(W26227));
  INVX1 G44385 (.I(W14307), .ZN(W24509));
  INVX1 G44386 (.I(W11583), .ZN(W24510));
  INVX1 G44387 (.I(W7638), .ZN(W24670));
  INVX1 G44388 (.I(W2250), .ZN(W26221));
  INVX1 G44389 (.I(W5735), .ZN(W24513));
  INVX1 G44390 (.I(W22330), .ZN(W26219));
  INVX1 G44391 (.I(W1145), .ZN(O3682));
  INVX1 G44392 (.I(W6252), .ZN(W26216));
  INVX1 G44393 (.I(W21420), .ZN(O3681));
  INVX1 G44394 (.I(W14741), .ZN(W24515));
  INVX1 G44395 (.I(W10541), .ZN(W24517));
  INVX1 G44396 (.I(W5756), .ZN(O3679));
  INVX1 G44397 (.I(W873), .ZN(O3196));
  INVX1 G44398 (.I(W12321), .ZN(W25930));
  INVX1 G44399 (.I(W15801), .ZN(W24782));
  INVX1 G44400 (.I(W9687), .ZN(W24784));
  INVX1 G44401 (.I(W5908), .ZN(W24786));
  INVX1 G44402 (.I(W25811), .ZN(O3579));
  INVX1 G44403 (.I(W10683), .ZN(W25923));
  INVX1 G44404 (.I(W15074), .ZN(W25921));
  INVX1 G44405 (.I(W23059), .ZN(W25919));
  INVX1 G44406 (.I(W5195), .ZN(O3577));
  INVX1 G44407 (.I(W5237), .ZN(O3575));
  INVX1 G44408 (.I(I100), .ZN(W24781));
  INVX1 G44409 (.I(W291), .ZN(O3197));
  INVX1 G44410 (.I(W10141), .ZN(W24799));
  INVX1 G44411 (.I(W22372), .ZN(W25906));
  INVX1 G44412 (.I(W1017), .ZN(W24801));
  INVX1 G44413 (.I(W24460), .ZN(W24802));
  INVX1 G44414 (.I(W20245), .ZN(W25902));
  INVX1 G44415 (.I(W21696), .ZN(O3198));
  INVX1 G44416 (.I(W15458), .ZN(W25898));
  INVX1 G44417 (.I(W2909), .ZN(O3566));
  INVX1 G44418 (.I(W23899), .ZN(W24770));
  INVX1 G44419 (.I(W24517), .ZN(O3186));
  INVX1 G44420 (.I(W174), .ZN(W24759));
  INVX1 G44421 (.I(W24127), .ZN(W24760));
  INVX1 G44422 (.I(W15845), .ZN(W25954));
  INVX1 G44423 (.I(W6836), .ZN(O3586));
  INVX1 G44424 (.I(W12322), .ZN(W25951));
  INVX1 G44425 (.I(W12039), .ZN(W24764));
  INVX1 G44426 (.I(W22510), .ZN(W24765));
  INVX1 G44427 (.I(W3390), .ZN(O3189));
  INVX1 G44428 (.I(W800), .ZN(W25894));
  INVX1 G44429 (.I(W18229), .ZN(W25944));
  INVX1 G44430 (.I(W16174), .ZN(W25943));
  INVX1 G44431 (.I(W15681), .ZN(W24771));
  INVX1 G44432 (.I(W14561), .ZN(W24773));
  INVX1 G44433 (.I(W799), .ZN(O3584));
  INVX1 G44434 (.I(W14543), .ZN(W24774));
  INVX1 G44435 (.I(W21119), .ZN(W25936));
  INVX1 G44436 (.I(W21448), .ZN(O3583));
  INVX1 G44437 (.I(W906), .ZN(W25932));
  INVX1 G44438 (.I(W9524), .ZN(W24850));
  INVX1 G44439 (.I(W5893), .ZN(W24842));
  INVX1 G44440 (.I(W22260), .ZN(W24846));
  INVX1 G44441 (.I(W24094), .ZN(W25859));
  INVX1 G44442 (.I(W24585), .ZN(O3553));
  INVX1 G44443 (.I(W22888), .ZN(O3552));
  INVX1 G44444 (.I(W24207), .ZN(O3551));
  INVX1 G44445 (.I(W18106), .ZN(W25855));
  INVX1 G44446 (.I(W15383), .ZN(W25854));
  INVX1 G44447 (.I(W17202), .ZN(W25851));
  INVX1 G44448 (.I(W17153), .ZN(O3556));
  INVX1 G44449 (.I(W7914), .ZN(W25849));
  INVX1 G44450 (.I(W9852), .ZN(O3216));
  INVX1 G44451 (.I(W12932), .ZN(W25847));
  INVX1 G44452 (.I(W8227), .ZN(W24857));
  INVX1 G44453 (.I(W10459), .ZN(W24861));
  INVX1 G44454 (.I(W17180), .ZN(W25842));
  INVX1 G44455 (.I(W24518), .ZN(W25841));
  INVX1 G44456 (.I(W9636), .ZN(W25838));
  INVX1 G44457 (.I(W9949), .ZN(W25837));
  INVX1 G44458 (.I(W22070), .ZN(O3203));
  INVX1 G44459 (.I(W1734), .ZN(W25891));
  INVX1 G44460 (.I(W11561), .ZN(O3199));
  INVX1 G44461 (.I(W16300), .ZN(W25888));
  INVX1 G44462 (.I(W7948), .ZN(O3565));
  INVX1 G44463 (.I(W8819), .ZN(W25886));
  INVX1 G44464 (.I(W13499), .ZN(W25885));
  INVX1 G44465 (.I(W5128), .ZN(O3564));
  INVX1 G44466 (.I(W14695), .ZN(O3200));
  INVX1 G44467 (.I(I10), .ZN(W24821));
  INVX1 G44468 (.I(W14055), .ZN(O3185));
  INVX1 G44469 (.I(W4855), .ZN(O3205));
  INVX1 G44470 (.I(W2621), .ZN(W24830));
  INVX1 G44471 (.I(W20069), .ZN(W24833));
  INVX1 G44472 (.I(I1807), .ZN(W24834));
  INVX1 G44473 (.I(W20310), .ZN(O3560));
  INVX1 G44474 (.I(W22184), .ZN(W25870));
  INVX1 G44475 (.I(W1984), .ZN(W25869));
  INVX1 G44476 (.I(W20163), .ZN(W25868));
  INVX1 G44477 (.I(W18959), .ZN(O3558));
  INVX1 G44478 (.I(W12777), .ZN(O3167));
  INVX1 G44479 (.I(W8337), .ZN(O3609));
  INVX1 G44480 (.I(W16393), .ZN(W26039));
  INVX1 G44481 (.I(W19845), .ZN(W26038));
  INVX1 G44482 (.I(W16233), .ZN(W26037));
  INVX1 G44483 (.I(W18995), .ZN(W26034));
  INVX1 G44484 (.I(W19461), .ZN(O3166));
  INVX1 G44485 (.I(W22527), .ZN(W24694));
  INVX1 G44486 (.I(W15926), .ZN(W24695));
  INVX1 G44487 (.I(W5207), .ZN(W24696));
  INVX1 G44488 (.I(W19179), .ZN(O3162));
  INVX1 G44489 (.I(W9214), .ZN(W26026));
  INVX1 G44490 (.I(W13694), .ZN(W24702));
  INVX1 G44491 (.I(W214), .ZN(W26024));
  INVX1 G44492 (.I(W15844), .ZN(W24703));
  INVX1 G44493 (.I(W14447), .ZN(W26022));
  INVX1 G44494 (.I(W23628), .ZN(W24704));
  INVX1 G44495 (.I(W2720), .ZN(W26019));
  INVX1 G44496 (.I(I1902), .ZN(O3169));
  INVX1 G44497 (.I(W8158), .ZN(W26017));
  INVX1 G44498 (.I(W17526), .ZN(W26056));
  INVX1 G44499 (.I(W16592), .ZN(W26066));
  INVX1 G44500 (.I(I1872), .ZN(W24671));
  INVX1 G44501 (.I(W23177), .ZN(W24672));
  INVX1 G44502 (.I(W16262), .ZN(W24673));
  INVX1 G44503 (.I(W9312), .ZN(W26062));
  INVX1 G44504 (.I(W1981), .ZN(O3159));
  INVX1 G44505 (.I(W15715), .ZN(W26059));
  INVX1 G44506 (.I(W24770), .ZN(O3616));
  INVX1 G44507 (.I(W9203), .ZN(O3615));
  INVX1 G44508 (.I(W22754), .ZN(W24710));
  INVX1 G44509 (.I(W10344), .ZN(W24678));
  INVX1 G44510 (.I(W11876), .ZN(O3613));
  INVX1 G44511 (.I(W6999), .ZN(W24680));
  INVX1 G44512 (.I(W21325), .ZN(W26050));
  INVX1 G44513 (.I(W12875), .ZN(O3161));
  INVX1 G44514 (.I(W24981), .ZN(W26048));
  INVX1 G44515 (.I(W23287), .ZN(W26047));
  INVX1 G44516 (.I(W18515), .ZN(O3610));
  INVX1 G44517 (.I(W921), .ZN(W26045));
  INVX1 G44518 (.I(W17982), .ZN(W24751));
  INVX1 G44519 (.I(W21521), .ZN(W25981));
  INVX1 G44520 (.I(W1409), .ZN(W24739));
  INVX1 G44521 (.I(W957), .ZN(W24740));
  INVX1 G44522 (.I(W6137), .ZN(W25978));
  INVX1 G44523 (.I(W12560), .ZN(W25976));
  INVX1 G44524 (.I(W16864), .ZN(W25975));
  INVX1 G44525 (.I(W497), .ZN(W24742));
  INVX1 G44526 (.I(W8168), .ZN(W24744));
  INVX1 G44527 (.I(W17549), .ZN(O3182));
  INVX1 G44528 (.I(W18545), .ZN(W24735));
  INVX1 G44529 (.I(W22541), .ZN(W24752));
  INVX1 G44530 (.I(W18430), .ZN(W24755));
  INVX1 G44531 (.I(W7416), .ZN(O3588));
  INVX1 G44532 (.I(W24913), .ZN(W25964));
  INVX1 G44533 (.I(W3546), .ZN(O3587));
  INVX1 G44534 (.I(W23152), .ZN(O3184));
  INVX1 G44535 (.I(I1318), .ZN(W25961));
  INVX1 G44536 (.I(W9091), .ZN(W25960));
  INVX1 G44537 (.I(W3097), .ZN(W25959));
  INVX1 G44538 (.I(W15240), .ZN(W24724));
  INVX1 G44539 (.I(I1040), .ZN(W24711));
  INVX1 G44540 (.I(W8955), .ZN(W26013));
  INVX1 G44541 (.I(W16931), .ZN(W26012));
  INVX1 G44542 (.I(W9011), .ZN(W24712));
  INVX1 G44543 (.I(W10244), .ZN(W24717));
  INVX1 G44544 (.I(W1469), .ZN(O3172));
  INVX1 G44545 (.I(W65), .ZN(W26004));
  INVX1 G44546 (.I(W17748), .ZN(W26003));
  INVX1 G44547 (.I(W12101), .ZN(O3599));
  INVX1 G44548 (.I(W10021), .ZN(O2785));
  INVX1 G44549 (.I(W21729), .ZN(W24726));
  INVX1 G44550 (.I(W10471), .ZN(W25995));
  INVX1 G44551 (.I(W19448), .ZN(W24728));
  INVX1 G44552 (.I(W10046), .ZN(W25992));
  INVX1 G44553 (.I(W18615), .ZN(O3593));
  INVX1 G44554 (.I(W14965), .ZN(W25989));
  INVX1 G44555 (.I(W21881), .ZN(W25988));
  INVX1 G44556 (.I(W9391), .ZN(W25985));
  INVX1 G44557 (.I(W22102), .ZN(W25984));
  INVX1 G44558 (.I(W3334), .ZN(W22243));
  INVX1 G44559 (.I(W23905), .ZN(O4533));
  INVX1 G44560 (.I(W12388), .ZN(W22225));
  INVX1 G44561 (.I(W43), .ZN(O4531));
  INVX1 G44562 (.I(W28435), .ZN(W28530));
  INVX1 G44563 (.I(W14119), .ZN(O2455));
  INVX1 G44564 (.I(W7950), .ZN(W28526));
  INVX1 G44565 (.I(W7833), .ZN(W28525));
  INVX1 G44566 (.I(W14242), .ZN(W22233));
  INVX1 G44567 (.I(W4030), .ZN(W22235));
  INVX1 G44568 (.I(W7760), .ZN(W28521));
  INVX1 G44569 (.I(W19144), .ZN(O2452));
  INVX1 G44570 (.I(W19363), .ZN(O4526));
  INVX1 G44571 (.I(W15721), .ZN(O2459));
  INVX1 G44572 (.I(W12323), .ZN(O4524));
  INVX1 G44573 (.I(W5352), .ZN(W22250));
  INVX1 G44574 (.I(W19552), .ZN(W22253));
  INVX1 G44575 (.I(W7106), .ZN(W22256));
  INVX1 G44576 (.I(W4282), .ZN(W28506));
  INVX1 G44577 (.I(W322), .ZN(O2460));
  INVX1 G44578 (.I(W13390), .ZN(W28504));
  INVX1 G44579 (.I(W6374), .ZN(W22212));
  INVX1 G44580 (.I(W12135), .ZN(W22198));
  INVX1 G44581 (.I(W2574), .ZN(O2445));
  INVX1 G44582 (.I(W6916), .ZN(W22203));
  INVX1 G44583 (.I(W22143), .ZN(W22204));
  INVX1 G44584 (.I(I1945), .ZN(W22206));
  INVX1 G44585 (.I(W6523), .ZN(W28555));
  INVX1 G44586 (.I(W23434), .ZN(W28554));
  INVX1 G44587 (.I(W14074), .ZN(W28553));
  INVX1 G44588 (.I(W8891), .ZN(W28551));
  INVX1 G44589 (.I(W7543), .ZN(W22260));
  INVX1 G44590 (.I(W25550), .ZN(O4536));
  INVX1 G44591 (.I(W1352), .ZN(W22213));
  INVX1 G44592 (.I(W12442), .ZN(W22214));
  INVX1 G44593 (.I(W5441), .ZN(W28544));
  INVX1 G44594 (.I(W14640), .ZN(W28543));
  INVX1 G44595 (.I(W12285), .ZN(W22218));
  INVX1 G44596 (.I(W25739), .ZN(W28541));
  INVX1 G44597 (.I(W22023), .ZN(W28539));
  INVX1 G44598 (.I(W16809), .ZN(W22220));
  INVX1 G44599 (.I(W12357), .ZN(O4510));
  INVX1 G44600 (.I(W6982), .ZN(W22292));
  INVX1 G44601 (.I(W19562), .ZN(W22293));
  INVX1 G44602 (.I(W19680), .ZN(W22294));
  INVX1 G44603 (.I(W25978), .ZN(W28466));
  INVX1 G44604 (.I(W6548), .ZN(W22297));
  INVX1 G44605 (.I(W10316), .ZN(O2470));
  INVX1 G44606 (.I(W16953), .ZN(W28463));
  INVX1 G44607 (.I(W20665), .ZN(W28462));
  INVX1 G44608 (.I(W3436), .ZN(W28461));
  INVX1 G44609 (.I(W12994), .ZN(O2468));
  INVX1 G44610 (.I(W14078), .ZN(W22302));
  INVX1 G44611 (.I(W3838), .ZN(O2475));
  INVX1 G44612 (.I(W12396), .ZN(O4507));
  INVX1 G44613 (.I(W11941), .ZN(W22307));
  INVX1 G44614 (.I(W19846), .ZN(O2476));
  INVX1 G44615 (.I(W14294), .ZN(W22311));
  INVX1 G44616 (.I(W7597), .ZN(W28447));
  INVX1 G44617 (.I(W19308), .ZN(O4503));
  INVX1 G44618 (.I(W2864), .ZN(W28445));
  INVX1 G44619 (.I(W7865), .ZN(W22276));
  INVX1 G44620 (.I(W28453), .ZN(W28501));
  INVX1 G44621 (.I(W20248), .ZN(W22261));
  INVX1 G44622 (.I(W5850), .ZN(W28497));
  INVX1 G44623 (.I(W14032), .ZN(W22265));
  INVX1 G44624 (.I(W5450), .ZN(W22269));
  INVX1 G44625 (.I(I786), .ZN(W28494));
  INVX1 G44626 (.I(W13633), .ZN(O2463));
  INVX1 G44627 (.I(W13776), .ZN(O4519));
  INVX1 G44628 (.I(W12251), .ZN(W28488));
  INVX1 G44629 (.I(W7467), .ZN(W22197));
  INVX1 G44630 (.I(W3902), .ZN(O2464));
  INVX1 G44631 (.I(W10893), .ZN(W22279));
  INVX1 G44632 (.I(W3977), .ZN(W22282));
  INVX1 G44633 (.I(W6673), .ZN(W28481));
  INVX1 G44634 (.I(W2641), .ZN(W22284));
  INVX1 G44635 (.I(W15555), .ZN(O2466));
  INVX1 G44636 (.I(W19604), .ZN(O2467));
  INVX1 G44637 (.I(W7149), .ZN(W22287));
  INVX1 G44638 (.I(W19948), .ZN(W28475));
  INVX1 G44639 (.I(W3781), .ZN(W28634));
  INVX1 G44640 (.I(W12373), .ZN(W22126));
  INVX1 G44641 (.I(W14879), .ZN(W28647));
  INVX1 G44642 (.I(W5567), .ZN(W28644));
  INVX1 G44643 (.I(W8881), .ZN(O4568));
  INVX1 G44644 (.I(W16435), .ZN(W22132));
  INVX1 G44645 (.I(W6534), .ZN(O4565));
  INVX1 G44646 (.I(W2121), .ZN(W22134));
  INVX1 G44647 (.I(W14820), .ZN(W28637));
  INVX1 G44648 (.I(W19800), .ZN(O4564));
  INVX1 G44649 (.I(W15226), .ZN(W22135));
  INVX1 G44650 (.I(W19908), .ZN(W28650));
  INVX1 G44651 (.I(W25009), .ZN(O4562));
  INVX1 G44652 (.I(W14817), .ZN(O4561));
  INVX1 G44653 (.I(W10102), .ZN(O2434));
  INVX1 G44654 (.I(W21681), .ZN(W22154));
  INVX1 G44655 (.I(W21826), .ZN(W22155));
  INVX1 G44656 (.I(W20967), .ZN(W22156));
  INVX1 G44657 (.I(W15551), .ZN(W22157));
  INVX1 G44658 (.I(W14465), .ZN(W22158));
  INVX1 G44659 (.I(W20089), .ZN(W28615));
  INVX1 G44660 (.I(W20214), .ZN(O4575));
  INVX1 G44661 (.I(W10157), .ZN(W28683));
  INVX1 G44662 (.I(W18301), .ZN(W22093));
  INVX1 G44663 (.I(W1298), .ZN(O2423));
  INVX1 G44664 (.I(W13872), .ZN(W28671));
  INVX1 G44665 (.I(W18814), .ZN(O4577));
  INVX1 G44666 (.I(W6487), .ZN(W22103));
  INVX1 G44667 (.I(W21799), .ZN(O2425));
  INVX1 G44668 (.I(W11255), .ZN(W28666));
  INVX1 G44669 (.I(W21769), .ZN(W22107));
  INVX1 G44670 (.I(W11652), .ZN(W22160));
  INVX1 G44671 (.I(W13436), .ZN(W22108));
  INVX1 G44672 (.I(W6058), .ZN(W22109));
  INVX1 G44673 (.I(W287), .ZN(O2427));
  INVX1 G44674 (.I(W3360), .ZN(W22113));
  INVX1 G44675 (.I(W6392), .ZN(W22114));
  INVX1 G44676 (.I(W11811), .ZN(W28655));
  INVX1 G44677 (.I(I712), .ZN(W22116));
  INVX1 G44678 (.I(W14378), .ZN(W28653));
  INVX1 G44679 (.I(I1572), .ZN(W22123));
  INVX1 G44680 (.I(W10314), .ZN(W28573));
  INVX1 G44681 (.I(W14960), .ZN(O2442));
  INVX1 G44682 (.I(W5260), .ZN(W28583));
  INVX1 G44683 (.I(W11838), .ZN(W22186));
  INVX1 G44684 (.I(W1052), .ZN(W22187));
  INVX1 G44685 (.I(W3803), .ZN(W22188));
  INVX1 G44686 (.I(W16546), .ZN(W28578));
  INVX1 G44687 (.I(W6416), .ZN(W28577));
  INVX1 G44688 (.I(W12420), .ZN(W22190));
  INVX1 G44689 (.I(W20428), .ZN(W28574));
  INVX1 G44690 (.I(W19613), .ZN(W28585));
  INVX1 G44691 (.I(W2691), .ZN(W22192));
  INVX1 G44692 (.I(I780), .ZN(W22193));
  INVX1 G44693 (.I(W22583), .ZN(O4545));
  INVX1 G44694 (.I(W3530), .ZN(W22194));
  INVX1 G44695 (.I(W20292), .ZN(W28568));
  INVX1 G44696 (.I(W18737), .ZN(W28567));
  INVX1 G44697 (.I(W22548), .ZN(O4544));
  INVX1 G44698 (.I(I1386), .ZN(W22195));
  INVX1 G44699 (.I(W11559), .ZN(W28563));
  INVX1 G44700 (.I(W13817), .ZN(O2436));
  INVX1 G44701 (.I(I1782), .ZN(W28613));
  INVX1 G44702 (.I(W21792), .ZN(W28612));
  INVX1 G44703 (.I(W24290), .ZN(W28611));
  INVX1 G44704 (.I(W12949), .ZN(O4559));
  INVX1 G44705 (.I(W4691), .ZN(O4558));
  INVX1 G44706 (.I(W577), .ZN(W28608));
  INVX1 G44707 (.I(W25435), .ZN(W28607));
  INVX1 G44708 (.I(W2015), .ZN(W22163));
  INVX1 G44709 (.I(I188), .ZN(W28604));
  INVX1 G44710 (.I(W11433), .ZN(W22315));
  INVX1 G44711 (.I(W10717), .ZN(O2437));
  INVX1 G44712 (.I(W3511), .ZN(W22172));
  INVX1 G44713 (.I(W5884), .ZN(W22174));
  INVX1 G44714 (.I(W15698), .ZN(W22175));
  INVX1 G44715 (.I(W7561), .ZN(W28596));
  INVX1 G44716 (.I(W11201), .ZN(O4552));
  INVX1 G44717 (.I(W22070), .ZN(W22180));
  INVX1 G44718 (.I(W12653), .ZN(O4550));
  INVX1 G44719 (.I(W3653), .ZN(O2441));
  INVX1 G44720 (.I(W11015), .ZN(W28278));
  INVX1 G44721 (.I(W28257), .ZN(O4431));
  INVX1 G44722 (.I(W8559), .ZN(O4430));
  INVX1 G44723 (.I(W3726), .ZN(W22439));
  INVX1 G44724 (.I(W2332), .ZN(W28285));
  INVX1 G44725 (.I(W14477), .ZN(W28284));
  INVX1 G44726 (.I(W2057), .ZN(O4429));
  INVX1 G44727 (.I(W22166), .ZN(O4428));
  INVX1 G44728 (.I(W18015), .ZN(W22442));
  INVX1 G44729 (.I(W5853), .ZN(W28280));
  INVX1 G44730 (.I(W2119), .ZN(W22445));
  INVX1 G44731 (.I(W8190), .ZN(W28289));
  INVX1 G44732 (.I(W10816), .ZN(W22449));
  INVX1 G44733 (.I(W3131), .ZN(W22452));
  INVX1 G44734 (.I(W8745), .ZN(W22454));
  INVX1 G44735 (.I(W14241), .ZN(O4423));
  INVX1 G44736 (.I(W13552), .ZN(O2518));
  INVX1 G44737 (.I(W4064), .ZN(W22457));
  INVX1 G44738 (.I(W9129), .ZN(O2522));
  INVX1 G44739 (.I(W22188), .ZN(W22468));
  INVX1 G44740 (.I(W3746), .ZN(W28261));
  INVX1 G44741 (.I(W3369), .ZN(O4436));
  INVX1 G44742 (.I(W2268), .ZN(O2504));
  INVX1 G44743 (.I(W27269), .ZN(W28319));
  INVX1 G44744 (.I(I1304), .ZN(O2506));
  INVX1 G44745 (.I(W10361), .ZN(W22417));
  INVX1 G44746 (.I(W2545), .ZN(O4442));
  INVX1 G44747 (.I(W27897), .ZN(O4441));
  INVX1 G44748 (.I(W19043), .ZN(W22424));
  INVX1 G44749 (.I(W12854), .ZN(O2510));
  INVX1 G44750 (.I(W27023), .ZN(O4437));
  INVX1 G44751 (.I(I1426), .ZN(W22478));
  INVX1 G44752 (.I(W10487), .ZN(W28300));
  INVX1 G44753 (.I(W4702), .ZN(W28299));
  INVX1 G44754 (.I(W3005), .ZN(W28298));
  INVX1 G44755 (.I(W17908), .ZN(W22433));
  INVX1 G44756 (.I(W15653), .ZN(W28296));
  INVX1 G44757 (.I(I1983), .ZN(O2513));
  INVX1 G44758 (.I(I991), .ZN(O4433));
  INVX1 G44759 (.I(W18874), .ZN(W28291));
  INVX1 G44760 (.I(I1618), .ZN(O2514));
  INVX1 G44761 (.I(W12919), .ZN(W28220));
  INVX1 G44762 (.I(W10604), .ZN(W28234));
  INVX1 G44763 (.I(I1293), .ZN(W22505));
  INVX1 G44764 (.I(W5521), .ZN(O2538));
  INVX1 G44765 (.I(W16570), .ZN(O4409));
  INVX1 G44766 (.I(W21386), .ZN(W28228));
  INVX1 G44767 (.I(W4074), .ZN(O2539));
  INVX1 G44768 (.I(W3620), .ZN(W22515));
  INVX1 G44769 (.I(W1616), .ZN(W22516));
  INVX1 G44770 (.I(I1868), .ZN(W22519));
  INVX1 G44771 (.I(I467), .ZN(W28235));
  INVX1 G44772 (.I(W398), .ZN(W22525));
  INVX1 G44773 (.I(W20070), .ZN(W28217));
  INVX1 G44774 (.I(W22045), .ZN(W28215));
  INVX1 G44775 (.I(W2980), .ZN(W22532));
  INVX1 G44776 (.I(W10348), .ZN(O2544));
  INVX1 G44777 (.I(W2645), .ZN(W22538));
  INVX1 G44778 (.I(W17903), .ZN(W22539));
  INVX1 G44779 (.I(W16403), .ZN(W28206));
  INVX1 G44780 (.I(W20108), .ZN(O4398));
  INVX1 G44781 (.I(W20633), .ZN(W28248));
  INVX1 G44782 (.I(W5957), .ZN(O4420));
  INVX1 G44783 (.I(W5933), .ZN(W28257));
  INVX1 G44784 (.I(W13289), .ZN(W28256));
  INVX1 G44785 (.I(W11683), .ZN(W22482));
  INVX1 G44786 (.I(W11062), .ZN(W22483));
  INVX1 G44787 (.I(W16837), .ZN(W28252));
  INVX1 G44788 (.I(W11709), .ZN(O2530));
  INVX1 G44789 (.I(I683), .ZN(W28250));
  INVX1 G44790 (.I(W11421), .ZN(O4419));
  INVX1 G44791 (.I(W15568), .ZN(O2503));
  INVX1 G44792 (.I(W7449), .ZN(W28247));
  INVX1 G44793 (.I(W9681), .ZN(O4418));
  INVX1 G44794 (.I(W22453), .ZN(W22487));
  INVX1 G44795 (.I(I698), .ZN(W22488));
  INVX1 G44796 (.I(W9082), .ZN(W22493));
  INVX1 G44797 (.I(W23241), .ZN(O4414));
  INVX1 G44798 (.I(W19823), .ZN(W22496));
  INVX1 G44799 (.I(W6655), .ZN(O2534));
  INVX1 G44800 (.I(W2813), .ZN(W28236));
  INVX1 G44801 (.I(W4187), .ZN(O4478));
  INVX1 G44802 (.I(W10547), .ZN(W28400));
  INVX1 G44803 (.I(W2295), .ZN(W22355));
  INVX1 G44804 (.I(W23882), .ZN(W28398));
  INVX1 G44805 (.I(W16784), .ZN(W22356));
  INVX1 G44806 (.I(W19648), .ZN(W28395));
  INVX1 G44807 (.I(W9873), .ZN(W28393));
  INVX1 G44808 (.I(W5712), .ZN(O2488));
  INVX1 G44809 (.I(W8213), .ZN(W28391));
  INVX1 G44810 (.I(W9313), .ZN(W22364));
  INVX1 G44811 (.I(W3290), .ZN(O4482));
  INVX1 G44812 (.I(W18428), .ZN(O2490));
  INVX1 G44813 (.I(W4056), .ZN(W28386));
  INVX1 G44814 (.I(W17593), .ZN(O4477));
  INVX1 G44815 (.I(W21676), .ZN(O4476));
  INVX1 G44816 (.I(W25779), .ZN(W28382));
  INVX1 G44817 (.I(W6307), .ZN(W22372));
  INVX1 G44818 (.I(W16116), .ZN(O4472));
  INVX1 G44819 (.I(W14750), .ZN(O4471));
  INVX1 G44820 (.I(W5685), .ZN(W28377));
  INVX1 G44821 (.I(W25608), .ZN(W28420));
  INVX1 G44822 (.I(W14481), .ZN(W28441));
  INVX1 G44823 (.I(W18476), .ZN(W28438));
  INVX1 G44824 (.I(W18754), .ZN(O4500));
  INVX1 G44825 (.I(W16613), .ZN(O4499));
  INVX1 G44826 (.I(I1806), .ZN(O2480));
  INVX1 G44827 (.I(I358), .ZN(W22321));
  INVX1 G44828 (.I(W25656), .ZN(W28429));
  INVX1 G44829 (.I(W17984), .ZN(W22329));
  INVX1 G44830 (.I(I804), .ZN(W22332));
  INVX1 G44831 (.I(W21762), .ZN(W22374));
  INVX1 G44832 (.I(W11143), .ZN(W28419));
  INVX1 G44833 (.I(W14475), .ZN(W28416));
  INVX1 G44834 (.I(W4773), .ZN(W22341));
  INVX1 G44835 (.I(W4718), .ZN(W28413));
  INVX1 G44836 (.I(I263), .ZN(W22342));
  INVX1 G44837 (.I(W10679), .ZN(W22346));
  INVX1 G44838 (.I(W20980), .ZN(W22347));
  INVX1 G44839 (.I(W21012), .ZN(O4484));
  INVX1 G44840 (.I(W11490), .ZN(W22352));
  INVX1 G44841 (.I(W13679), .ZN(O4452));
  INVX1 G44842 (.I(W22637), .ZN(O4460));
  INVX1 G44843 (.I(W6411), .ZN(W22396));
  INVX1 G44844 (.I(W20480), .ZN(O4458));
  INVX1 G44845 (.I(W6342), .ZN(O4457));
  INVX1 G44846 (.I(W2568), .ZN(W28342));
  INVX1 G44847 (.I(W9559), .ZN(W22397));
  INVX1 G44848 (.I(W6887), .ZN(W28339));
  INVX1 G44849 (.I(W4190), .ZN(W22399));
  INVX1 G44850 (.I(W16577), .ZN(W22400));
  INVX1 G44851 (.I(W18892), .ZN(O2498));
  INVX1 G44852 (.I(W15757), .ZN(O4451));
  INVX1 G44853 (.I(W5056), .ZN(O4450));
  INVX1 G44854 (.I(W480), .ZN(W28330));
  INVX1 G44855 (.I(W18623), .ZN(O2501));
  INVX1 G44856 (.I(W13417), .ZN(W22407));
  INVX1 G44857 (.I(W10392), .ZN(O2502));
  INVX1 G44858 (.I(W19293), .ZN(O4448));
  INVX1 G44859 (.I(I288), .ZN(W28324));
  INVX1 G44860 (.I(W2652), .ZN(O4447));
  INVX1 G44861 (.I(I1330), .ZN(W22383));
  INVX1 G44862 (.I(W12824), .ZN(W28374));
  INVX1 G44863 (.I(W8149), .ZN(O2491));
  INVX1 G44864 (.I(W6983), .ZN(W22376));
  INVX1 G44865 (.I(W14819), .ZN(W22377));
  INVX1 G44866 (.I(W17149), .ZN(O2493));
  INVX1 G44867 (.I(W968), .ZN(W22381));
  INVX1 G44868 (.I(W26817), .ZN(W28365));
  INVX1 G44869 (.I(W1133), .ZN(O4468));
  INVX1 G44870 (.I(W19980), .ZN(W28363));
  INVX1 G44871 (.I(W4663), .ZN(W22088));
  INVX1 G44872 (.I(W7063), .ZN(W28361));
  INVX1 G44873 (.I(I82), .ZN(W22384));
  INVX1 G44874 (.I(W18274), .ZN(W22386));
  INVX1 G44875 (.I(W9461), .ZN(W22387));
  INVX1 G44876 (.I(W2003), .ZN(O4466));
  INVX1 G44877 (.I(W23527), .ZN(O4465));
  INVX1 G44878 (.I(W3782), .ZN(W28355));
  INVX1 G44879 (.I(W12342), .ZN(W28354));
  INVX1 G44880 (.I(W25823), .ZN(O4461));
  INVX1 G44881 (.I(W8391), .ZN(O2333));
  INVX1 G44882 (.I(W2936), .ZN(W21775));
  INVX1 G44883 (.I(W10692), .ZN(W21776));
  INVX1 G44884 (.I(W239), .ZN(O2329));
  INVX1 G44885 (.I(W16308), .ZN(W21778));
  INVX1 G44886 (.I(W8957), .ZN(W21780));
  INVX1 G44887 (.I(I1580), .ZN(O2330));
  INVX1 G44888 (.I(W21741), .ZN(O4702));
  INVX1 G44889 (.I(W26310), .ZN(W29012));
  INVX1 G44890 (.I(W6815), .ZN(O4701));
  INVX1 G44891 (.I(W16687), .ZN(O2332));
  INVX1 G44892 (.I(W5903), .ZN(O4707));
  INVX1 G44893 (.I(W15813), .ZN(W21788));
  INVX1 G44894 (.I(W3986), .ZN(W29005));
  INVX1 G44895 (.I(W1846), .ZN(W21791));
  INVX1 G44896 (.I(W28099), .ZN(W29001));
  INVX1 G44897 (.I(W20483), .ZN(W29000));
  INVX1 G44898 (.I(W17117), .ZN(W28997));
  INVX1 G44899 (.I(W1110), .ZN(W21795));
  INVX1 G44900 (.I(W17500), .ZN(W28995));
  INVX1 G44901 (.I(W10625), .ZN(O2336));
  INVX1 G44902 (.I(W13712), .ZN(W21764));
  INVX1 G44903 (.I(W17553), .ZN(O2326));
  INVX1 G44904 (.I(W6690), .ZN(O4719));
  INVX1 G44905 (.I(W12157), .ZN(W29045));
  INVX1 G44906 (.I(W8275), .ZN(W21758));
  INVX1 G44907 (.I(W9013), .ZN(W29043));
  INVX1 G44908 (.I(W971), .ZN(W29042));
  INVX1 G44909 (.I(W12490), .ZN(W29040));
  INVX1 G44910 (.I(W23749), .ZN(W29039));
  INVX1 G44911 (.I(W4777), .ZN(O4717));
  INVX1 G44912 (.I(W8728), .ZN(W21800));
  INVX1 G44913 (.I(W1475), .ZN(W21765));
  INVX1 G44914 (.I(W7706), .ZN(O4714));
  INVX1 G44915 (.I(W645), .ZN(W21766));
  INVX1 G44916 (.I(W12368), .ZN(O4713));
  INVX1 G44917 (.I(W16457), .ZN(O4711));
  INVX1 G44918 (.I(W27111), .ZN(W29027));
  INVX1 G44919 (.I(W13220), .ZN(W21770));
  INVX1 G44920 (.I(W4732), .ZN(W21771));
  INVX1 G44921 (.I(W9695), .ZN(W21773));
  INVX1 G44922 (.I(W11645), .ZN(O2350));
  INVX1 G44923 (.I(W18697), .ZN(W28961));
  INVX1 G44924 (.I(W28559), .ZN(W28960));
  INVX1 G44925 (.I(W5380), .ZN(W21833));
  INVX1 G44926 (.I(W7919), .ZN(W21835));
  INVX1 G44927 (.I(I1898), .ZN(W21838));
  INVX1 G44928 (.I(W24248), .ZN(O4678));
  INVX1 G44929 (.I(W13253), .ZN(W21840));
  INVX1 G44930 (.I(W6746), .ZN(O4677));
  INVX1 G44931 (.I(W5593), .ZN(O2349));
  INVX1 G44932 (.I(W6194), .ZN(O4682));
  INVX1 G44933 (.I(W20564), .ZN(W21845));
  INVX1 G44934 (.I(W26311), .ZN(W28945));
  INVX1 G44935 (.I(W7993), .ZN(W28944));
  INVX1 G44936 (.I(W25223), .ZN(O4674));
  INVX1 G44937 (.I(W7061), .ZN(O4673));
  INVX1 G44938 (.I(W9028), .ZN(O4672));
  INVX1 G44939 (.I(W1898), .ZN(W28938));
  INVX1 G44940 (.I(W4749), .ZN(O4671));
  INVX1 G44941 (.I(W4291), .ZN(W21853));
  INVX1 G44942 (.I(W27636), .ZN(O4690));
  INVX1 G44943 (.I(I1682), .ZN(W28989));
  INVX1 G44944 (.I(W9553), .ZN(W21801));
  INVX1 G44945 (.I(W9056), .ZN(W21802));
  INVX1 G44946 (.I(W21559), .ZN(O2337));
  INVX1 G44947 (.I(W12741), .ZN(W21805));
  INVX1 G44948 (.I(W17772), .ZN(W21810));
  INVX1 G44949 (.I(W16755), .ZN(W21811));
  INVX1 G44950 (.I(I1368), .ZN(O2339));
  INVX1 G44951 (.I(W18241), .ZN(O2340));
  INVX1 G44952 (.I(W9633), .ZN(W21754));
  INVX1 G44953 (.I(W14074), .ZN(O4689));
  INVX1 G44954 (.I(W22790), .ZN(O4688));
  INVX1 G44955 (.I(W7523), .ZN(O2341));
  INVX1 G44956 (.I(W23149), .ZN(W28974));
  INVX1 G44957 (.I(W295), .ZN(O4684));
  INVX1 G44958 (.I(W265), .ZN(W21827));
  INVX1 G44959 (.I(W15044), .ZN(O2346));
  INVX1 G44960 (.I(W12346), .ZN(W28965));
  INVX1 G44961 (.I(W12181), .ZN(W28964));
  INVX1 G44962 (.I(W9765), .ZN(W21652));
  INVX1 G44963 (.I(W1546), .ZN(O2302));
  INVX1 G44964 (.I(I936), .ZN(W21645));
  INVX1 G44965 (.I(W11133), .ZN(W29147));
  INVX1 G44966 (.I(W20782), .ZN(W29146));
  INVX1 G44967 (.I(W20654), .ZN(W21646));
  INVX1 G44968 (.I(I812), .ZN(W29144));
  INVX1 G44969 (.I(W14658), .ZN(W21648));
  INVX1 G44970 (.I(W23165), .ZN(O4765));
  INVX1 G44971 (.I(W4472), .ZN(O2303));
  INVX1 G44972 (.I(W13318), .ZN(W29151));
  INVX1 G44973 (.I(W27411), .ZN(W29138));
  INVX1 G44974 (.I(W12399), .ZN(W21656));
  INVX1 G44975 (.I(W18906), .ZN(W21657));
  INVX1 G44976 (.I(W23706), .ZN(W29134));
  INVX1 G44977 (.I(W12979), .ZN(W21658));
  INVX1 G44978 (.I(W12974), .ZN(W29131));
  INVX1 G44979 (.I(W18579), .ZN(W21664));
  INVX1 G44980 (.I(W14555), .ZN(O4759));
  INVX1 G44981 (.I(W10783), .ZN(W21666));
  INVX1 G44982 (.I(I271), .ZN(W21627));
  INVX1 G44983 (.I(W16831), .ZN(W21606));
  INVX1 G44984 (.I(W1031), .ZN(W21608));
  INVX1 G44985 (.I(W6415), .ZN(O2293));
  INVX1 G44986 (.I(I64), .ZN(W29175));
  INVX1 G44987 (.I(W15220), .ZN(W29173));
  INVX1 G44988 (.I(W3237), .ZN(W21614));
  INVX1 G44989 (.I(W20221), .ZN(W29171));
  INVX1 G44990 (.I(W16587), .ZN(W21620));
  INVX1 G44991 (.I(W7999), .ZN(O2298));
  INVX1 G44992 (.I(W19464), .ZN(W21668));
  INVX1 G44993 (.I(W1718), .ZN(W21628));
  INVX1 G44994 (.I(W11535), .ZN(W21630));
  INVX1 G44995 (.I(W25018), .ZN(W29162));
  INVX1 G44996 (.I(W5292), .ZN(O2300));
  INVX1 G44997 (.I(W1479), .ZN(W29158));
  INVX1 G44998 (.I(W19836), .ZN(W21635));
  INVX1 G44999 (.I(W16314), .ZN(W29156));
  INVX1 G45000 (.I(W24692), .ZN(O4768));
  INVX1 G45001 (.I(W16432), .ZN(W21640));
  INVX1 G45002 (.I(W403), .ZN(W21737));
  INVX1 G45003 (.I(W6561), .ZN(W21717));
  INVX1 G45004 (.I(W21831), .ZN(O4735));
  INVX1 G45005 (.I(W26264), .ZN(W29082));
  INVX1 G45006 (.I(W3910), .ZN(O4733));
  INVX1 G45007 (.I(W2768), .ZN(W21720));
  INVX1 G45008 (.I(W16386), .ZN(W21721));
  INVX1 G45009 (.I(W209), .ZN(W21724));
  INVX1 G45010 (.I(W7767), .ZN(O4728));
  INVX1 G45011 (.I(W24685), .ZN(O4726));
  INVX1 G45012 (.I(W7467), .ZN(W21716));
  INVX1 G45013 (.I(W6403), .ZN(O2320));
  INVX1 G45014 (.I(W15332), .ZN(W21741));
  INVX1 G45015 (.I(W18929), .ZN(O2324));
  INVX1 G45016 (.I(W12530), .ZN(W21745));
  INVX1 G45017 (.I(W13329), .ZN(W29056));
  INVX1 G45018 (.I(I1742), .ZN(W21747));
  INVX1 G45019 (.I(W28554), .ZN(W29053));
  INVX1 G45020 (.I(W12973), .ZN(W29052));
  INVX1 G45021 (.I(W21976), .ZN(W29050));
  INVX1 G45022 (.I(W17133), .ZN(W21698));
  INVX1 G45023 (.I(W3615), .ZN(W21674));
  INVX1 G45024 (.I(W2213), .ZN(W21682));
  INVX1 G45025 (.I(W4351), .ZN(W21688));
  INVX1 G45026 (.I(W8530), .ZN(O4750));
  INVX1 G45027 (.I(W6338), .ZN(W29110));
  INVX1 G45028 (.I(W10176), .ZN(O4749));
  INVX1 G45029 (.I(W1361), .ZN(W29107));
  INVX1 G45030 (.I(I904), .ZN(O4747));
  INVX1 G45031 (.I(W13905), .ZN(O4745));
  INVX1 G45032 (.I(W16972), .ZN(W28935));
  INVX1 G45033 (.I(W14336), .ZN(O2313));
  INVX1 G45034 (.I(W8252), .ZN(O2314));
  INVX1 G45035 (.I(W7201), .ZN(W29098));
  INVX1 G45036 (.I(W1229), .ZN(O4742));
  INVX1 G45037 (.I(W4792), .ZN(W21710));
  INVX1 G45038 (.I(W11343), .ZN(W29090));
  INVX1 G45039 (.I(W2777), .ZN(W21715));
  INVX1 G45040 (.I(W23776), .ZN(W29087));
  INVX1 G45041 (.I(W6968), .ZN(O4737));
  INVX1 G45042 (.I(W7008), .ZN(W22019));
  INVX1 G45043 (.I(W1626), .ZN(W28776));
  INVX1 G45044 (.I(W12317), .ZN(O4614));
  INVX1 G45045 (.I(W14615), .ZN(O2397));
  INVX1 G45046 (.I(W4848), .ZN(O4613));
  INVX1 G45047 (.I(W18959), .ZN(W22014));
  INVX1 G45048 (.I(W17870), .ZN(W28769));
  INVX1 G45049 (.I(W23503), .ZN(O4610));
  INVX1 G45050 (.I(W5780), .ZN(O4609));
  INVX1 G45051 (.I(W13888), .ZN(O4608));
  INVX1 G45052 (.I(I1939), .ZN(W22018));
  INVX1 G45053 (.I(W16680), .ZN(W22006));
  INVX1 G45054 (.I(W19356), .ZN(O4606));
  INVX1 G45055 (.I(W2391), .ZN(O2406));
  INVX1 G45056 (.I(W21896), .ZN(W28752));
  INVX1 G45057 (.I(W7543), .ZN(W22029));
  INVX1 G45058 (.I(W5572), .ZN(W28749));
  INVX1 G45059 (.I(I426), .ZN(W22035));
  INVX1 G45060 (.I(W12321), .ZN(W22039));
  INVX1 G45061 (.I(W5050), .ZN(W22041));
  INVX1 G45062 (.I(W17501), .ZN(O4602));
  INVX1 G45063 (.I(I1013), .ZN(W28795));
  INVX1 G45064 (.I(W2337), .ZN(W21968));
  INVX1 G45065 (.I(W6346), .ZN(W28811));
  INVX1 G45066 (.I(W2648), .ZN(W28807));
  INVX1 G45067 (.I(W28429), .ZN(W28806));
  INVX1 G45068 (.I(W28142), .ZN(W28803));
  INVX1 G45069 (.I(I1267), .ZN(W21983));
  INVX1 G45070 (.I(W5749), .ZN(O4623));
  INVX1 G45071 (.I(I1123), .ZN(W21987));
  INVX1 G45072 (.I(I1754), .ZN(W21988));
  INVX1 G45073 (.I(W26255), .ZN(W28743));
  INVX1 G45074 (.I(W594), .ZN(W21993));
  INVX1 G45075 (.I(W12055), .ZN(W28792));
  INVX1 G45076 (.I(W4040), .ZN(O4618));
  INVX1 G45077 (.I(W22571), .ZN(O4616));
  INVX1 G45078 (.I(W5610), .ZN(W22002));
  INVX1 G45079 (.I(W15458), .ZN(W28784));
  INVX1 G45080 (.I(W8156), .ZN(W22003));
  INVX1 G45081 (.I(W27621), .ZN(O4615));
  INVX1 G45082 (.I(W6473), .ZN(W28781));
  INVX1 G45083 (.I(W18442), .ZN(O2419));
  INVX1 G45084 (.I(W8590), .ZN(W28712));
  INVX1 G45085 (.I(W4822), .ZN(W28711));
  INVX1 G45086 (.I(W3283), .ZN(W22063));
  INVX1 G45087 (.I(W398), .ZN(W28709));
  INVX1 G45088 (.I(W21118), .ZN(O2417));
  INVX1 G45089 (.I(W10996), .ZN(W22074));
  INVX1 G45090 (.I(W8063), .ZN(O4583));
  INVX1 G45091 (.I(W15557), .ZN(W28700));
  INVX1 G45092 (.I(W28351), .ZN(W28699));
  INVX1 G45093 (.I(W21690), .ZN(O2415));
  INVX1 G45094 (.I(W15478), .ZN(W28697));
  INVX1 G45095 (.I(W28618), .ZN(W28695));
  INVX1 G45096 (.I(W19700), .ZN(W28694));
  INVX1 G45097 (.I(W3386), .ZN(W22078));
  INVX1 G45098 (.I(W11966), .ZN(W22079));
  INVX1 G45099 (.I(W1823), .ZN(O2420));
  INVX1 G45100 (.I(W17634), .ZN(O4582));
  INVX1 G45101 (.I(W13835), .ZN(O4581));
  INVX1 G45102 (.I(W16151), .ZN(W28685));
  INVX1 G45103 (.I(W26166), .ZN(W28730));
  INVX1 G45104 (.I(W6230), .ZN(W22043));
  INVX1 G45105 (.I(W5019), .ZN(O4600));
  INVX1 G45106 (.I(W12620), .ZN(W22044));
  INVX1 G45107 (.I(W12855), .ZN(O4598));
  INVX1 G45108 (.I(W9824), .ZN(W28738));
  INVX1 G45109 (.I(W27471), .ZN(O4597));
  INVX1 G45110 (.I(W18916), .ZN(O4596));
  INVX1 G45111 (.I(I507), .ZN(W28734));
  INVX1 G45112 (.I(W2317), .ZN(O4594));
  INVX1 G45113 (.I(W9214), .ZN(W28814));
  INVX1 G45114 (.I(W7328), .ZN(O4593));
  INVX1 G45115 (.I(W21492), .ZN(W28727));
  INVX1 G45116 (.I(W12721), .ZN(W28725));
  INVX1 G45117 (.I(W14079), .ZN(O4592));
  INVX1 G45118 (.I(W27188), .ZN(W28723));
  INVX1 G45119 (.I(W11618), .ZN(O4591));
  INVX1 G45120 (.I(W11537), .ZN(W28721));
  INVX1 G45121 (.I(W7355), .ZN(W22053));
  INVX1 G45122 (.I(W951), .ZN(W28718));
  INVX1 G45123 (.I(W1955), .ZN(O2368));
  INVX1 G45124 (.I(W13166), .ZN(O2362));
  INVX1 G45125 (.I(W15640), .ZN(W21880));
  INVX1 G45126 (.I(W13606), .ZN(W28905));
  INVX1 G45127 (.I(W3316), .ZN(O4662));
  INVX1 G45128 (.I(W19526), .ZN(O4661));
  INVX1 G45129 (.I(W10757), .ZN(W21884));
  INVX1 G45130 (.I(W8882), .ZN(O4657));
  INVX1 G45131 (.I(W8482), .ZN(W28896));
  INVX1 G45132 (.I(W28656), .ZN(O4654));
  INVX1 G45133 (.I(W6517), .ZN(W28909));
  INVX1 G45134 (.I(I895), .ZN(W21893));
  INVX1 G45135 (.I(W17702), .ZN(W28889));
  INVX1 G45136 (.I(W15854), .ZN(W28888));
  INVX1 G45137 (.I(I834), .ZN(W28884));
  INVX1 G45138 (.I(W9491), .ZN(W21903));
  INVX1 G45139 (.I(W20703), .ZN(W21904));
  INVX1 G45140 (.I(W19119), .ZN(W28879));
  INVX1 G45141 (.I(W2640), .ZN(W21905));
  INVX1 G45142 (.I(W17463), .ZN(O4648));
  INVX1 G45143 (.I(I1286), .ZN(W21862));
  INVX1 G45144 (.I(W8998), .ZN(W28934));
  INVX1 G45145 (.I(W15775), .ZN(W28933));
  INVX1 G45146 (.I(W24641), .ZN(O4670));
  INVX1 G45147 (.I(W5046), .ZN(W21854));
  INVX1 G45148 (.I(W15704), .ZN(W28930));
  INVX1 G45149 (.I(W8972), .ZN(W21855));
  INVX1 G45150 (.I(W18601), .ZN(W21856));
  INVX1 G45151 (.I(W6799), .ZN(O4668));
  INVX1 G45152 (.I(W23039), .ZN(O4667));
  INVX1 G45153 (.I(W15802), .ZN(W21907));
  INVX1 G45154 (.I(W17573), .ZN(O2355));
  INVX1 G45155 (.I(I1523), .ZN(W28921));
  INVX1 G45156 (.I(W16461), .ZN(W28920));
  INVX1 G45157 (.I(W8362), .ZN(W21866));
  INVX1 G45158 (.I(W13002), .ZN(O2356));
  INVX1 G45159 (.I(W8859), .ZN(O2358));
  INVX1 G45160 (.I(W16124), .ZN(W21871));
  INVX1 G45161 (.I(W13718), .ZN(W21873));
  INVX1 G45162 (.I(W5071), .ZN(O2360));
  INVX1 G45163 (.I(W25802), .ZN(W28828));
  INVX1 G45164 (.I(W10471), .ZN(O4634));
  INVX1 G45165 (.I(W5016), .ZN(W28841));
  INVX1 G45166 (.I(W20492), .ZN(W21940));
  INVX1 G45167 (.I(W7258), .ZN(W28837));
  INVX1 G45168 (.I(I1535), .ZN(O2381));
  INVX1 G45169 (.I(W6585), .ZN(O2382));
  INVX1 G45170 (.I(W13089), .ZN(W21945));
  INVX1 G45171 (.I(W11954), .ZN(W21948));
  INVX1 G45172 (.I(I755), .ZN(W21950));
  INVX1 G45173 (.I(W1318), .ZN(W28846));
  INVX1 G45174 (.I(W17184), .ZN(W28827));
  INVX1 G45175 (.I(I1477), .ZN(W21954));
  INVX1 G45176 (.I(W17555), .ZN(W21955));
  INVX1 G45177 (.I(W9391), .ZN(O2385));
  INVX1 G45178 (.I(W18407), .ZN(O2386));
  INVX1 G45179 (.I(W8118), .ZN(O2387));
  INVX1 G45180 (.I(W26447), .ZN(W28818));
  INVX1 G45181 (.I(W4994), .ZN(W21967));
  INVX1 G45182 (.I(W15417), .ZN(W28815));
  INVX1 G45183 (.I(W9058), .ZN(W28862));
  INVX1 G45184 (.I(W5569), .ZN(W28874));
  INVX1 G45185 (.I(W24814), .ZN(W28873));
  INVX1 G45186 (.I(W26511), .ZN(W28872));
  INVX1 G45187 (.I(W18344), .ZN(W21910));
  INVX1 G45188 (.I(W26393), .ZN(O4646));
  INVX1 G45189 (.I(W17999), .ZN(W28869));
  INVX1 G45190 (.I(W10820), .ZN(W21911));
  INVX1 G45191 (.I(W12836), .ZN(O2374));
  INVX1 G45192 (.I(W8956), .ZN(W21915));
  INVX1 G45193 (.I(W6085), .ZN(W22544));
  INVX1 G45194 (.I(W16863), .ZN(O2375));
  INVX1 G45195 (.I(W736), .ZN(W21918));
  INVX1 G45196 (.I(W19095), .ZN(W21919));
  INVX1 G45197 (.I(W4004), .ZN(O4640));
  INVX1 G45198 (.I(W5300), .ZN(W21924));
  INVX1 G45199 (.I(W15827), .ZN(W21927));
  INVX1 G45200 (.I(W5698), .ZN(W21928));
  INVX1 G45201 (.I(W10390), .ZN(W28849));
  INVX1 G45202 (.I(W17232), .ZN(W21930));
  INVX1 G45203 (.I(W15152), .ZN(W23160));
  INVX1 G45204 (.I(W6953), .ZN(O2690));
  INVX1 G45205 (.I(W3343), .ZN(W23145));
  INVX1 G45206 (.I(W13924), .ZN(O2693));
  INVX1 G45207 (.I(W25084), .ZN(W27585));
  INVX1 G45208 (.I(W21134), .ZN(O4154));
  INVX1 G45209 (.I(I1209), .ZN(W23157));
  INVX1 G45210 (.I(W14766), .ZN(O4153));
  INVX1 G45211 (.I(W10113), .ZN(W23158));
  INVX1 G45212 (.I(W19279), .ZN(W23159));
  INVX1 G45213 (.I(W17988), .ZN(W27577));
  INVX1 G45214 (.I(I970), .ZN(O4159));
  INVX1 G45215 (.I(W15970), .ZN(W23163));
  INVX1 G45216 (.I(W11533), .ZN(W27573));
  INVX1 G45217 (.I(W21044), .ZN(W27572));
  INVX1 G45218 (.I(W1635), .ZN(W27570));
  INVX1 G45219 (.I(W2477), .ZN(O2695));
  INVX1 G45220 (.I(W1143), .ZN(O4150));
  INVX1 G45221 (.I(W9598), .ZN(W27567));
  INVX1 G45222 (.I(W16466), .ZN(W27566));
  INVX1 G45223 (.I(W609), .ZN(W23167));
  INVX1 G45224 (.I(W14169), .ZN(W23112));
  INVX1 G45225 (.I(W17173), .ZN(W27629));
  INVX1 G45226 (.I(W22598), .ZN(W27628));
  INVX1 G45227 (.I(W16870), .ZN(W23104));
  INVX1 G45228 (.I(W5266), .ZN(W27626));
  INVX1 G45229 (.I(W3565), .ZN(W23106));
  INVX1 G45230 (.I(W19000), .ZN(W27624));
  INVX1 G45231 (.I(W17430), .ZN(W23108));
  INVX1 G45232 (.I(I1287), .ZN(W23109));
  INVX1 G45233 (.I(W529), .ZN(W27618));
  INVX1 G45234 (.I(W463), .ZN(W27563));
  INVX1 G45235 (.I(W7056), .ZN(W27613));
  INVX1 G45236 (.I(W23013), .ZN(O4166));
  INVX1 G45237 (.I(W369), .ZN(W27610));
  INVX1 G45238 (.I(W16406), .ZN(W27609));
  INVX1 G45239 (.I(I781), .ZN(O4164));
  INVX1 G45240 (.I(W13608), .ZN(O2682));
  INVX1 G45241 (.I(W11636), .ZN(W27599));
  INVX1 G45242 (.I(W27433), .ZN(W27595));
  INVX1 G45243 (.I(W3051), .ZN(W27594));
  INVX1 G45244 (.I(W13449), .ZN(W23223));
  INVX1 G45245 (.I(W6032), .ZN(O4139));
  INVX1 G45246 (.I(W12130), .ZN(W27531));
  INVX1 G45247 (.I(W16726), .ZN(O4138));
  INVX1 G45248 (.I(W3327), .ZN(W23206));
  INVX1 G45249 (.I(W2045), .ZN(W27526));
  INVX1 G45250 (.I(W23050), .ZN(O2710));
  INVX1 G45251 (.I(W11731), .ZN(W23214));
  INVX1 G45252 (.I(W21145), .ZN(W23216));
  INVX1 G45253 (.I(W7954), .ZN(W23222));
  INVX1 G45254 (.I(W6093), .ZN(O2707));
  INVX1 G45255 (.I(W15938), .ZN(O2714));
  INVX1 G45256 (.I(W8649), .ZN(W23229));
  INVX1 G45257 (.I(W18718), .ZN(W27514));
  INVX1 G45258 (.I(W16557), .ZN(W27512));
  INVX1 G45259 (.I(W1334), .ZN(W23232));
  INVX1 G45260 (.I(W20583), .ZN(W23233));
  INVX1 G45261 (.I(W13574), .ZN(O2717));
  INVX1 G45262 (.I(W13386), .ZN(O4129));
  INVX1 G45263 (.I(I1468), .ZN(O2718));
  INVX1 G45264 (.I(I1738), .ZN(O4145));
  INVX1 G45265 (.I(W14545), .ZN(W23170));
  INVX1 G45266 (.I(W450), .ZN(O4148));
  INVX1 G45267 (.I(W3433), .ZN(O4147));
  INVX1 G45268 (.I(W3843), .ZN(O2696));
  INVX1 G45269 (.I(W10495), .ZN(W23173));
  INVX1 G45270 (.I(W13754), .ZN(W27557));
  INVX1 G45271 (.I(W11093), .ZN(W27556));
  INVX1 G45272 (.I(W9092), .ZN(W27555));
  INVX1 G45273 (.I(I1153), .ZN(O2697));
  INVX1 G45274 (.I(W15999), .ZN(W27630));
  INVX1 G45275 (.I(W9572), .ZN(W23178));
  INVX1 G45276 (.I(W20345), .ZN(W23179));
  INVX1 G45277 (.I(W8721), .ZN(O2699));
  INVX1 G45278 (.I(W9852), .ZN(W27546));
  INVX1 G45279 (.I(W16351), .ZN(O2700));
  INVX1 G45280 (.I(I32), .ZN(W27543));
  INVX1 G45281 (.I(W14362), .ZN(W23188));
  INVX1 G45282 (.I(I335), .ZN(W23192));
  INVX1 G45283 (.I(W5745), .ZN(W27535));
  INVX1 G45284 (.I(W23356), .ZN(W27703));
  INVX1 G45285 (.I(W10615), .ZN(O2664));
  INVX1 G45286 (.I(W26792), .ZN(W27715));
  INVX1 G45287 (.I(W2983), .ZN(W27714));
  INVX1 G45288 (.I(W8405), .ZN(W27712));
  INVX1 G45289 (.I(W10869), .ZN(W23028));
  INVX1 G45290 (.I(W10262), .ZN(O4204));
  INVX1 G45291 (.I(W12724), .ZN(O4203));
  INVX1 G45292 (.I(W15465), .ZN(O4202));
  INVX1 G45293 (.I(W27337), .ZN(W27704));
  INVX1 G45294 (.I(W8732), .ZN(W27719));
  INVX1 G45295 (.I(W19734), .ZN(W23039));
  INVX1 G45296 (.I(W5139), .ZN(W23040));
  INVX1 G45297 (.I(W14467), .ZN(W23041));
  INVX1 G45298 (.I(W1833), .ZN(O2668));
  INVX1 G45299 (.I(W11233), .ZN(O4197));
  INVX1 G45300 (.I(W4713), .ZN(W27692));
  INVX1 G45301 (.I(W751), .ZN(O4193));
  INVX1 G45302 (.I(W8326), .ZN(W23052));
  INVX1 G45303 (.I(I1727), .ZN(W23054));
  INVX1 G45304 (.I(W12008), .ZN(W27732));
  INVX1 G45305 (.I(W7339), .ZN(O2655));
  INVX1 G45306 (.I(W18992), .ZN(W23000));
  INVX1 G45307 (.I(W16863), .ZN(W23001));
  INVX1 G45308 (.I(W8806), .ZN(W27741));
  INVX1 G45309 (.I(W10044), .ZN(W27738));
  INVX1 G45310 (.I(W26826), .ZN(W27737));
  INVX1 G45311 (.I(W8525), .ZN(W23009));
  INVX1 G45312 (.I(W22738), .ZN(W23012));
  INVX1 G45313 (.I(W4779), .ZN(O2659));
  INVX1 G45314 (.I(W24246), .ZN(W27684));
  INVX1 G45315 (.I(W16554), .ZN(W23016));
  INVX1 G45316 (.I(W5168), .ZN(W27729));
  INVX1 G45317 (.I(W17329), .ZN(W23018));
  INVX1 G45318 (.I(W5334), .ZN(W27727));
  INVX1 G45319 (.I(W7078), .ZN(O2660));
  INVX1 G45320 (.I(W14349), .ZN(W23020));
  INVX1 G45321 (.I(W23291), .ZN(W27723));
  INVX1 G45322 (.I(W18098), .ZN(O2662));
  INVX1 G45323 (.I(W15634), .ZN(O4210));
  INVX1 G45324 (.I(W6212), .ZN(O4174));
  INVX1 G45325 (.I(W12358), .ZN(W23075));
  INVX1 G45326 (.I(W15906), .ZN(W23076));
  INVX1 G45327 (.I(W985), .ZN(W27657));
  INVX1 G45328 (.I(W8685), .ZN(W23077));
  INVX1 G45329 (.I(W26985), .ZN(O4178));
  INVX1 G45330 (.I(I626), .ZN(W23080));
  INVX1 G45331 (.I(W6915), .ZN(O4176));
  INVX1 G45332 (.I(W20130), .ZN(W27649));
  INVX1 G45333 (.I(W18077), .ZN(W23082));
  INVX1 G45334 (.I(W7585), .ZN(W23074));
  INVX1 G45335 (.I(W5509), .ZN(W23086));
  INVX1 G45336 (.I(W14999), .ZN(W23090));
  INVX1 G45337 (.I(W14348), .ZN(W23095));
  INVX1 G45338 (.I(I300), .ZN(O2676));
  INVX1 G45339 (.I(W22412), .ZN(W23097));
  INVX1 G45340 (.I(W13141), .ZN(W23099));
  INVX1 G45341 (.I(W27585), .ZN(O4170));
  INVX1 G45342 (.I(W5612), .ZN(W27632));
  INVX1 G45343 (.I(W11802), .ZN(W23103));
  INVX1 G45344 (.I(W2445), .ZN(O4186));
  INVX1 G45345 (.I(W9935), .ZN(W27682));
  INVX1 G45346 (.I(W17191), .ZN(O2670));
  INVX1 G45347 (.I(W27455), .ZN(O4191));
  INVX1 G45348 (.I(W14300), .ZN(O4190));
  INVX1 G45349 (.I(W2448), .ZN(O4189));
  INVX1 G45350 (.I(W20266), .ZN(W23059));
  INVX1 G45351 (.I(W8331), .ZN(O4188));
  INVX1 G45352 (.I(W10891), .ZN(W23061));
  INVX1 G45353 (.I(W20946), .ZN(W23062));
  INVX1 G45354 (.I(W26646), .ZN(W27505));
  INVX1 G45355 (.I(W19693), .ZN(W23064));
  INVX1 G45356 (.I(W14371), .ZN(W27669));
  INVX1 G45357 (.I(W15465), .ZN(W23066));
  INVX1 G45358 (.I(W2640), .ZN(W27667));
  INVX1 G45359 (.I(W23933), .ZN(O4183));
  INVX1 G45360 (.I(W20819), .ZN(O2673));
  INVX1 G45361 (.I(W683), .ZN(W27663));
  INVX1 G45362 (.I(W10019), .ZN(W23070));
  INVX1 G45363 (.I(W18100), .ZN(W23072));
  INVX1 G45364 (.I(W16925), .ZN(O2765));
  INVX1 G45365 (.I(W4789), .ZN(O4078));
  INVX1 G45366 (.I(W7922), .ZN(W23388));
  INVX1 G45367 (.I(W23300), .ZN(O4077));
  INVX1 G45368 (.I(W18730), .ZN(W23390));
  INVX1 G45369 (.I(W11430), .ZN(O2762));
  INVX1 G45370 (.I(W7620), .ZN(W23394));
  INVX1 G45371 (.I(W4440), .ZN(W23396));
  INVX1 G45372 (.I(W4113), .ZN(W23397));
  INVX1 G45373 (.I(W6327), .ZN(O2763));
  INVX1 G45374 (.I(W15866), .ZN(W27349));
  INVX1 G45375 (.I(W24526), .ZN(W27363));
  INVX1 G45376 (.I(W22689), .ZN(W23403));
  INVX1 G45377 (.I(W4232), .ZN(W23406));
  INVX1 G45378 (.I(W2219), .ZN(W23408));
  INVX1 G45379 (.I(W23813), .ZN(O4070));
  INVX1 G45380 (.I(W96), .ZN(O2766));
  INVX1 G45381 (.I(W15440), .ZN(W27339));
  INVX1 G45382 (.I(W142), .ZN(W27337));
  INVX1 G45383 (.I(W8073), .ZN(W27336));
  INVX1 G45384 (.I(W25487), .ZN(W27334));
  INVX1 G45385 (.I(W4276), .ZN(O4084));
  INVX1 G45386 (.I(W7197), .ZN(W23349));
  INVX1 G45387 (.I(I634), .ZN(W27390));
  INVX1 G45388 (.I(W9545), .ZN(O2749));
  INVX1 G45389 (.I(I1954), .ZN(W27388));
  INVX1 G45390 (.I(W17035), .ZN(O4087));
  INVX1 G45391 (.I(W11405), .ZN(O4086));
  INVX1 G45392 (.I(W18456), .ZN(W23362));
  INVX1 G45393 (.I(W17422), .ZN(O2751));
  INVX1 G45394 (.I(W14679), .ZN(W27380));
  INVX1 G45395 (.I(W6354), .ZN(W27333));
  INVX1 G45396 (.I(W26846), .ZN(O4083));
  INVX1 G45397 (.I(W17852), .ZN(W27376));
  INVX1 G45398 (.I(W4660), .ZN(W27375));
  INVX1 G45399 (.I(W7612), .ZN(W23370));
  INVX1 G45400 (.I(W14419), .ZN(W27371));
  INVX1 G45401 (.I(W21299), .ZN(W27369));
  INVX1 G45402 (.I(W11284), .ZN(W23375));
  INVX1 G45403 (.I(W8911), .ZN(O2756));
  INVX1 G45404 (.I(W10258), .ZN(W23385));
  INVX1 G45405 (.I(W26331), .ZN(W27286));
  INVX1 G45406 (.I(I61), .ZN(O2775));
  INVX1 G45407 (.I(I459), .ZN(W23446));
  INVX1 G45408 (.I(W20095), .ZN(O2777));
  INVX1 G45409 (.I(W22680), .ZN(W27295));
  INVX1 G45410 (.I(I17), .ZN(O2779));
  INVX1 G45411 (.I(W13568), .ZN(W23451));
  INVX1 G45412 (.I(W18004), .ZN(W23452));
  INVX1 G45413 (.I(W21093), .ZN(W23453));
  INVX1 G45414 (.I(W967), .ZN(W23454));
  INVX1 G45415 (.I(W11137), .ZN(O4057));
  INVX1 G45416 (.I(W15349), .ZN(O2783));
  INVX1 G45417 (.I(W13883), .ZN(O4052));
  INVX1 G45418 (.I(W13343), .ZN(W23460));
  INVX1 G45419 (.I(W16704), .ZN(W23461));
  INVX1 G45420 (.I(W2729), .ZN(W23464));
  INVX1 G45421 (.I(W20747), .ZN(W27278));
  INVX1 G45422 (.I(W3148), .ZN(W27277));
  INVX1 G45423 (.I(I874), .ZN(O4049));
  INVX1 G45424 (.I(W11259), .ZN(W27275));
  INVX1 G45425 (.I(W26810), .ZN(W27321));
  INVX1 G45426 (.I(W13251), .ZN(W23413));
  INVX1 G45427 (.I(W8171), .ZN(W27331));
  INVX1 G45428 (.I(W24981), .ZN(O4067));
  INVX1 G45429 (.I(W340), .ZN(W23414));
  INVX1 G45430 (.I(W13183), .ZN(W23416));
  INVX1 G45431 (.I(W24135), .ZN(O4065));
  INVX1 G45432 (.I(W7278), .ZN(W23417));
  INVX1 G45433 (.I(W1546), .ZN(W27324));
  INVX1 G45434 (.I(W15887), .ZN(W27323));
  INVX1 G45435 (.I(W11219), .ZN(W23345));
  INVX1 G45436 (.I(I1981), .ZN(W27319));
  INVX1 G45437 (.I(W3878), .ZN(O4064));
  INVX1 G45438 (.I(W4384), .ZN(O4063));
  INVX1 G45439 (.I(W10742), .ZN(W23426));
  INVX1 G45440 (.I(W10534), .ZN(W27313));
  INVX1 G45441 (.I(W6178), .ZN(W27311));
  INVX1 G45442 (.I(W1151), .ZN(O2772));
  INVX1 G45443 (.I(W7254), .ZN(W23440));
  INVX1 G45444 (.I(W7387), .ZN(O2774));
  INVX1 G45445 (.I(W7578), .ZN(O4115));
  INVX1 G45446 (.I(W4176), .ZN(W27479));
  INVX1 G45447 (.I(W22582), .ZN(O4118));
  INVX1 G45448 (.I(W14476), .ZN(O2728));
  INVX1 G45449 (.I(W4736), .ZN(W23265));
  INVX1 G45450 (.I(I240), .ZN(O4117));
  INVX1 G45451 (.I(W18381), .ZN(W23266));
  INVX1 G45452 (.I(I893), .ZN(O4116));
  INVX1 G45453 (.I(W17499), .ZN(W23269));
  INVX1 G45454 (.I(W8104), .ZN(W27465));
  INVX1 G45455 (.I(W6845), .ZN(O2726));
  INVX1 G45456 (.I(W22585), .ZN(O4114));
  INVX1 G45457 (.I(W9036), .ZN(W27462));
  INVX1 G45458 (.I(W940), .ZN(O4113));
  INVX1 G45459 (.I(W5827), .ZN(W27460));
  INVX1 G45460 (.I(W131), .ZN(O4112));
  INVX1 G45461 (.I(W271), .ZN(W23272));
  INVX1 G45462 (.I(I255), .ZN(O4111));
  INVX1 G45463 (.I(W20040), .ZN(W27455));
  INVX1 G45464 (.I(W20826), .ZN(O2733));
  INVX1 G45465 (.I(I896), .ZN(W27492));
  INVX1 G45466 (.I(W7448), .ZN(W27504));
  INVX1 G45467 (.I(I172), .ZN(W27501));
  INVX1 G45468 (.I(W18469), .ZN(O2721));
  INVX1 G45469 (.I(W1707), .ZN(W27499));
  INVX1 G45470 (.I(W14332), .ZN(W27497));
  INVX1 G45471 (.I(W19007), .ZN(W23246));
  INVX1 G45472 (.I(W3445), .ZN(W23248));
  INVX1 G45473 (.I(I1265), .ZN(W27494));
  INVX1 G45474 (.I(W7524), .ZN(O2722));
  INVX1 G45475 (.I(W8993), .ZN(O4109));
  INVX1 G45476 (.I(W6822), .ZN(O4122));
  INVX1 G45477 (.I(W9900), .ZN(W23250));
  INVX1 G45478 (.I(W16132), .ZN(W27489));
  INVX1 G45479 (.I(W6984), .ZN(W27488));
  INVX1 G45480 (.I(W4154), .ZN(W27487));
  INVX1 G45481 (.I(W19988), .ZN(W23251));
  INVX1 G45482 (.I(W22037), .ZN(W27484));
  INVX1 G45483 (.I(W17704), .ZN(O2724));
  INVX1 G45484 (.I(W7843), .ZN(W23255));
  INVX1 G45485 (.I(W8737), .ZN(W27410));
  INVX1 G45486 (.I(W984), .ZN(W27424));
  INVX1 G45487 (.I(W9469), .ZN(W23315));
  INVX1 G45488 (.I(W20526), .ZN(O4098));
  INVX1 G45489 (.I(W16352), .ZN(W23318));
  INVX1 G45490 (.I(W10488), .ZN(W23319));
  INVX1 G45491 (.I(W600), .ZN(O2742));
  INVX1 G45492 (.I(W6462), .ZN(W23327));
  INVX1 G45493 (.I(W5150), .ZN(O4096));
  INVX1 G45494 (.I(W576), .ZN(W27411));
  INVX1 G45495 (.I(W6966), .ZN(W27425));
  INVX1 G45496 (.I(W5889), .ZN(W27408));
  INVX1 G45497 (.I(W7584), .ZN(O4093));
  INVX1 G45498 (.I(W16185), .ZN(W27405));
  INVX1 G45499 (.I(W15422), .ZN(O4091));
  INVX1 G45500 (.I(W8281), .ZN(O4090));
  INVX1 G45501 (.I(W21942), .ZN(W27398));
  INVX1 G45502 (.I(W10104), .ZN(W23341));
  INVX1 G45503 (.I(W11616), .ZN(W23342));
  INVX1 G45504 (.I(W7981), .ZN(W23343));
  INVX1 G45505 (.I(W11091), .ZN(W27441));
  INVX1 G45506 (.I(W12779), .ZN(W23277));
  INVX1 G45507 (.I(W11150), .ZN(W27450));
  INVX1 G45508 (.I(W17537), .ZN(O4107));
  INVX1 G45509 (.I(W8106), .ZN(W27448));
  INVX1 G45510 (.I(W10411), .ZN(O2734));
  INVX1 G45511 (.I(W18985), .ZN(W23283));
  INVX1 G45512 (.I(W16198), .ZN(W23284));
  INVX1 G45513 (.I(I1310), .ZN(W23287));
  INVX1 G45514 (.I(W3805), .ZN(O4105));
  INVX1 G45515 (.I(W7262), .ZN(W22995));
  INVX1 G45516 (.I(W2704), .ZN(W23290));
  INVX1 G45517 (.I(W21748), .ZN(W27439));
  INVX1 G45518 (.I(W7999), .ZN(O2736));
  INVX1 G45519 (.I(W17797), .ZN(W23302));
  INVX1 G45520 (.I(W10179), .ZN(W23304));
  INVX1 G45521 (.I(W14333), .ZN(O2738));
  INVX1 G45522 (.I(W3453), .ZN(W23307));
  INVX1 G45523 (.I(W17148), .ZN(O2739));
  INVX1 G45524 (.I(W20583), .ZN(W23310));
  INVX1 G45525 (.I(W2371), .ZN(O4327));
  INVX1 G45526 (.I(W12667), .ZN(W22681));
  INVX1 G45527 (.I(W10591), .ZN(W22682));
  INVX1 G45528 (.I(W11752), .ZN(W28060));
  INVX1 G45529 (.I(W15367), .ZN(W28059));
  INVX1 G45530 (.I(W676), .ZN(W22683));
  INVX1 G45531 (.I(W286), .ZN(W22684));
  INVX1 G45532 (.I(W8470), .ZN(O4331));
  INVX1 G45533 (.I(W20156), .ZN(O4330));
  INVX1 G45534 (.I(W24478), .ZN(O4329));
  INVX1 G45535 (.I(W16465), .ZN(O2584));
  INVX1 G45536 (.I(W8786), .ZN(W22678));
  INVX1 G45537 (.I(W21106), .ZN(W22697));
  INVX1 G45538 (.I(W14017), .ZN(O2587));
  INVX1 G45539 (.I(W13012), .ZN(W22701));
  INVX1 G45540 (.I(W27087), .ZN(W28043));
  INVX1 G45541 (.I(W731), .ZN(W28042));
  INVX1 G45542 (.I(W5399), .ZN(W28040));
  INVX1 G45543 (.I(W15385), .ZN(O4323));
  INVX1 G45544 (.I(W16164), .ZN(W22707));
  INVX1 G45545 (.I(W25636), .ZN(W28035));
  INVX1 G45546 (.I(W6238), .ZN(W22664));
  INVX1 G45547 (.I(W13929), .ZN(O2566));
  INVX1 G45548 (.I(W8394), .ZN(W28087));
  INVX1 G45549 (.I(W14557), .ZN(O2568));
  INVX1 G45550 (.I(W23785), .ZN(O4342));
  INVX1 G45551 (.I(I1839), .ZN(W22656));
  INVX1 G45552 (.I(W17496), .ZN(W22657));
  INVX1 G45553 (.I(W2986), .ZN(O2572));
  INVX1 G45554 (.I(W9950), .ZN(W28079));
  INVX1 G45555 (.I(W10836), .ZN(O2573));
  INVX1 G45556 (.I(W1480), .ZN(W22719));
  INVX1 G45557 (.I(W4781), .ZN(O4338));
  INVX1 G45558 (.I(W21805), .ZN(W28074));
  INVX1 G45559 (.I(W3541), .ZN(O2576));
  INVX1 G45560 (.I(W4279), .ZN(O2578));
  INVX1 G45561 (.I(W70), .ZN(W28070));
  INVX1 G45562 (.I(W21895), .ZN(W22674));
  INVX1 G45563 (.I(W23563), .ZN(O4336));
  INVX1 G45564 (.I(W8066), .ZN(W28066));
  INVX1 G45565 (.I(W4360), .ZN(O2581));
  INVX1 G45566 (.I(W21357), .ZN(O2603));
  INVX1 G45567 (.I(W11816), .ZN(W22750));
  INVX1 G45568 (.I(W8104), .ZN(W22754));
  INVX1 G45569 (.I(W13390), .ZN(W27993));
  INVX1 G45570 (.I(W14550), .ZN(O2602));
  INVX1 G45571 (.I(W21184), .ZN(W27991));
  INVX1 G45572 (.I(W10536), .ZN(W27990));
  INVX1 G45573 (.I(W8811), .ZN(W22758));
  INVX1 G45574 (.I(W23624), .ZN(W27988));
  INVX1 G45575 (.I(W19698), .ZN(W27986));
  INVX1 G45576 (.I(W2594), .ZN(O4309));
  INVX1 G45577 (.I(W13625), .ZN(W27984));
  INVX1 G45578 (.I(I1874), .ZN(W22762));
  INVX1 G45579 (.I(W16848), .ZN(O4306));
  INVX1 G45580 (.I(W15875), .ZN(O2605));
  INVX1 G45581 (.I(W5661), .ZN(W22765));
  INVX1 G45582 (.I(W1385), .ZN(W27978));
  INVX1 G45583 (.I(W18091), .ZN(W22768));
  INVX1 G45584 (.I(W2260), .ZN(O4301));
  INVX1 G45585 (.I(W1303), .ZN(O2608));
  INVX1 G45586 (.I(W10093), .ZN(O4312));
  INVX1 G45587 (.I(I1544), .ZN(W28029));
  INVX1 G45588 (.I(W17450), .ZN(W28027));
  INVX1 G45589 (.I(W7999), .ZN(W22725));
  INVX1 G45590 (.I(W23295), .ZN(O4315));
  INVX1 G45591 (.I(W3672), .ZN(O4314));
  INVX1 G45592 (.I(W11779), .ZN(W28019));
  INVX1 G45593 (.I(W19248), .ZN(W22731));
  INVX1 G45594 (.I(W11716), .ZN(W22733));
  INVX1 G45595 (.I(W14705), .ZN(O2595));
  INVX1 G45596 (.I(W15894), .ZN(O2565));
  INVX1 G45597 (.I(W436), .ZN(W28013));
  INVX1 G45598 (.I(W9918), .ZN(O2598));
  INVX1 G45599 (.I(W19794), .ZN(O2599));
  INVX1 G45600 (.I(W17450), .ZN(W28008));
  INVX1 G45601 (.I(W3831), .ZN(W22741));
  INVX1 G45602 (.I(W12719), .ZN(W22742));
  INVX1 G45603 (.I(W11314), .ZN(O4310));
  INVX1 G45604 (.I(W13814), .ZN(W28004));
  INVX1 G45605 (.I(W13334), .ZN(W22746));
  INVX1 G45606 (.I(W15173), .ZN(W28161));
  INVX1 G45607 (.I(W7455), .ZN(W22575));
  INVX1 G45608 (.I(W12412), .ZN(W22576));
  INVX1 G45609 (.I(W19751), .ZN(W28171));
  INVX1 G45610 (.I(W17835), .ZN(W22577));
  INVX1 G45611 (.I(I1074), .ZN(W22578));
  INVX1 G45612 (.I(W6946), .ZN(W22579));
  INVX1 G45613 (.I(W13709), .ZN(W22584));
  INVX1 G45614 (.I(W12057), .ZN(O4379));
  INVX1 G45615 (.I(W5808), .ZN(W22586));
  INVX1 G45616 (.I(W20931), .ZN(W22566));
  INVX1 G45617 (.I(W26193), .ZN(W28157));
  INVX1 G45618 (.I(W13662), .ZN(W22594));
  INVX1 G45619 (.I(I1594), .ZN(O4377));
  INVX1 G45620 (.I(W1479), .ZN(W28154));
  INVX1 G45621 (.I(W17913), .ZN(W22598));
  INVX1 G45622 (.I(W14632), .ZN(O4376));
  INVX1 G45623 (.I(W22893), .ZN(W28149));
  INVX1 G45624 (.I(W1415), .ZN(W22601));
  INVX1 G45625 (.I(I1306), .ZN(W28147));
  INVX1 G45626 (.I(W14566), .ZN(W28189));
  INVX1 G45627 (.I(W26901), .ZN(W28202));
  INVX1 G45628 (.I(W20508), .ZN(W22547));
  INVX1 G45629 (.I(W10307), .ZN(W22548));
  INVX1 G45630 (.I(W15694), .ZN(W28198));
  INVX1 G45631 (.I(W2103), .ZN(O4396));
  INVX1 G45632 (.I(W3742), .ZN(W28196));
  INVX1 G45633 (.I(W8475), .ZN(W22550));
  INVX1 G45634 (.I(W21632), .ZN(W22553));
  INVX1 G45635 (.I(W6944), .ZN(W22554));
  INVX1 G45636 (.I(W701), .ZN(O4374));
  INVX1 G45637 (.I(W5711), .ZN(O4390));
  INVX1 G45638 (.I(W8666), .ZN(W28186));
  INVX1 G45639 (.I(W8231), .ZN(O4389));
  INVX1 G45640 (.I(W4231), .ZN(W22559));
  INVX1 G45641 (.I(I1095), .ZN(W28182));
  INVX1 G45642 (.I(W4853), .ZN(W22560));
  INVX1 G45643 (.I(W1653), .ZN(W22564));
  INVX1 G45644 (.I(W1597), .ZN(O4385));
  INVX1 G45645 (.I(I1577), .ZN(W22565));
  INVX1 G45646 (.I(I108), .ZN(W22634));
  INVX1 G45647 (.I(W7342), .ZN(W22624));
  INVX1 G45648 (.I(W21846), .ZN(W28113));
  INVX1 G45649 (.I(W4956), .ZN(W28112));
  INVX1 G45650 (.I(W13273), .ZN(O4353));
  INVX1 G45651 (.I(I1541), .ZN(O4352));
  INVX1 G45652 (.I(W15064), .ZN(W22625));
  INVX1 G45653 (.I(W11415), .ZN(W22628));
  INVX1 G45654 (.I(W361), .ZN(W22630));
  INVX1 G45655 (.I(W13648), .ZN(W22632));
  INVX1 G45656 (.I(W15101), .ZN(O2560));
  INVX1 G45657 (.I(W1276), .ZN(W22635));
  INVX1 G45658 (.I(W20521), .ZN(O4348));
  INVX1 G45659 (.I(W19402), .ZN(W28098));
  INVX1 G45660 (.I(W24492), .ZN(O4347));
  INVX1 G45661 (.I(W15097), .ZN(W22639));
  INVX1 G45662 (.I(W4144), .ZN(W22640));
  INVX1 G45663 (.I(W10909), .ZN(O4344));
  INVX1 G45664 (.I(I1592), .ZN(W22642));
  INVX1 G45665 (.I(W17507), .ZN(O2563));
  INVX1 G45666 (.I(W22563), .ZN(W22610));
  INVX1 G45667 (.I(W7404), .ZN(O4373));
  INVX1 G45668 (.I(W40), .ZN(O4372));
  INVX1 G45669 (.I(W18920), .ZN(W22603));
  INVX1 G45670 (.I(W3179), .ZN(O4371));
  INVX1 G45671 (.I(W20139), .ZN(W28139));
  INVX1 G45672 (.I(W7831), .ZN(O4370));
  INVX1 G45673 (.I(W18526), .ZN(O2556));
  INVX1 G45674 (.I(W17034), .ZN(W22607));
  INVX1 G45675 (.I(W19157), .ZN(W28133));
  INVX1 G45676 (.I(W2494), .ZN(O2609));
  INVX1 G45677 (.I(W13022), .ZN(W22612));
  INVX1 G45678 (.I(W26069), .ZN(W28129));
  INVX1 G45679 (.I(W7908), .ZN(O4363));
  INVX1 G45680 (.I(W9118), .ZN(W28126));
  INVX1 G45681 (.I(W17081), .ZN(W22616));
  INVX1 G45682 (.I(W7245), .ZN(W28122));
  INVX1 G45683 (.I(W6877), .ZN(O4360));
  INVX1 G45684 (.I(W1307), .ZN(O4358));
  INVX1 G45685 (.I(W9235), .ZN(W22622));
  INVX1 G45686 (.I(W18873), .ZN(W22920));
  INVX1 G45687 (.I(W4958), .ZN(W27830));
  INVX1 G45688 (.I(W19220), .ZN(W22906));
  INVX1 G45689 (.I(W17561), .ZN(W22907));
  INVX1 G45690 (.I(W24699), .ZN(O4243));
  INVX1 G45691 (.I(W4427), .ZN(W22913));
  INVX1 G45692 (.I(W2244), .ZN(W22914));
  INVX1 G45693 (.I(I602), .ZN(O2636));
  INVX1 G45694 (.I(W13432), .ZN(W27819));
  INVX1 G45695 (.I(W12488), .ZN(W27818));
  INVX1 G45696 (.I(I208), .ZN(W22919));
  INVX1 G45697 (.I(W21027), .ZN(W27832));
  INVX1 G45698 (.I(W8743), .ZN(W22923));
  INVX1 G45699 (.I(W2072), .ZN(W22924));
  INVX1 G45700 (.I(W12310), .ZN(W22926));
  INVX1 G45701 (.I(W6927), .ZN(W27809));
  INVX1 G45702 (.I(W2134), .ZN(O4239));
  INVX1 G45703 (.I(W9929), .ZN(O2640));
  INVX1 G45704 (.I(W10782), .ZN(W27804));
  INVX1 G45705 (.I(W5540), .ZN(W22933));
  INVX1 G45706 (.I(W15570), .ZN(W27802));
  INVX1 G45707 (.I(W11760), .ZN(W27847));
  INVX1 G45708 (.I(W651), .ZN(W22877));
  INVX1 G45709 (.I(W9841), .ZN(W22882));
  INVX1 G45710 (.I(W24385), .ZN(O4255));
  INVX1 G45711 (.I(W19500), .ZN(W22883));
  INVX1 G45712 (.I(W2089), .ZN(O2627));
  INVX1 G45713 (.I(W13670), .ZN(W22889));
  INVX1 G45714 (.I(W4632), .ZN(W27852));
  INVX1 G45715 (.I(W4735), .ZN(O2629));
  INVX1 G45716 (.I(W6879), .ZN(O2630));
  INVX1 G45717 (.I(W21246), .ZN(W22934));
  INVX1 G45718 (.I(W20961), .ZN(W22895));
  INVX1 G45719 (.I(W14055), .ZN(W22899));
  INVX1 G45720 (.I(I618), .ZN(W27842));
  INVX1 G45721 (.I(W20161), .ZN(W27841));
  INVX1 G45722 (.I(W17267), .ZN(O4246));
  INVX1 G45723 (.I(W11084), .ZN(W27837));
  INVX1 G45724 (.I(W12374), .ZN(O2633));
  INVX1 G45725 (.I(W18186), .ZN(W27834));
  INVX1 G45726 (.I(W2511), .ZN(W27833));
  INVX1 G45727 (.I(W5342), .ZN(W22979));
  INVX1 G45728 (.I(W157), .ZN(W22963));
  INVX1 G45729 (.I(W9878), .ZN(W22966));
  INVX1 G45730 (.I(I1180), .ZN(O4224));
  INVX1 G45731 (.I(W11505), .ZN(W22967));
  INVX1 G45732 (.I(W7519), .ZN(W22968));
  INVX1 G45733 (.I(W24677), .ZN(W27763));
  INVX1 G45734 (.I(W6736), .ZN(W22973));
  INVX1 G45735 (.I(W20368), .ZN(W22974));
  INVX1 G45736 (.I(W10457), .ZN(W22976));
  INVX1 G45737 (.I(W14582), .ZN(W22962));
  INVX1 G45738 (.I(W1314), .ZN(O2650));
  INVX1 G45739 (.I(W20216), .ZN(W22984));
  INVX1 G45740 (.I(W10017), .ZN(W22988));
  INVX1 G45741 (.I(W14074), .ZN(W22989));
  INVX1 G45742 (.I(I825), .ZN(W22990));
  INVX1 G45743 (.I(W16544), .ZN(O2652));
  INVX1 G45744 (.I(W12356), .ZN(W22992));
  INVX1 G45745 (.I(W7772), .ZN(O2653));
  INVX1 G45746 (.I(W17960), .ZN(W22994));
  INVX1 G45747 (.I(W14961), .ZN(W22955));
  INVX1 G45748 (.I(W3096), .ZN(O2642));
  INVX1 G45749 (.I(W12180), .ZN(W27797));
  INVX1 G45750 (.I(W18933), .ZN(W27796));
  INVX1 G45751 (.I(W11221), .ZN(W27793));
  INVX1 G45752 (.I(W22872), .ZN(W22948));
  INVX1 G45753 (.I(W15091), .ZN(W22949));
  INVX1 G45754 (.I(W18274), .ZN(O4232));
  INVX1 G45755 (.I(W18686), .ZN(W22953));
  INVX1 G45756 (.I(W4693), .ZN(W27785));
  INVX1 G45757 (.I(W3293), .ZN(O2625));
  INVX1 G45758 (.I(W13044), .ZN(O2644));
  INVX1 G45759 (.I(W21572), .ZN(O4229));
  INVX1 G45760 (.I(W2347), .ZN(W27778));
  INVX1 G45761 (.I(W3526), .ZN(O4227));
  INVX1 G45762 (.I(W20403), .ZN(W22959));
  INVX1 G45763 (.I(W20672), .ZN(W22960));
  INVX1 G45764 (.I(W6267), .ZN(W22961));
  INVX1 G45765 (.I(W807), .ZN(W27773));
  INVX1 G45766 (.I(W6947), .ZN(W27772));
  INVX1 G45767 (.I(W6768), .ZN(O4282));
  INVX1 G45768 (.I(W20204), .ZN(W22798));
  INVX1 G45769 (.I(W13927), .ZN(W22799));
  INVX1 G45770 (.I(W5781), .ZN(O4288));
  INVX1 G45771 (.I(W11349), .ZN(W22800));
  INVX1 G45772 (.I(W19946), .ZN(W22810));
  INVX1 G45773 (.I(W20389), .ZN(W22812));
  INVX1 G45774 (.I(W20641), .ZN(W27931));
  INVX1 G45775 (.I(W12357), .ZN(W27930));
  INVX1 G45776 (.I(W7566), .ZN(W22813));
  INVX1 G45777 (.I(W9004), .ZN(W22795));
  INVX1 G45778 (.I(I1518), .ZN(W22816));
  INVX1 G45779 (.I(W11233), .ZN(W22819));
  INVX1 G45780 (.I(I1569), .ZN(W22821));
  INVX1 G45781 (.I(W16477), .ZN(W22823));
  INVX1 G45782 (.I(W13524), .ZN(O4278));
  INVX1 G45783 (.I(W16360), .ZN(W27916));
  INVX1 G45784 (.I(W18680), .ZN(W27914));
  INVX1 G45785 (.I(W5236), .ZN(W22829));
  INVX1 G45786 (.I(W13663), .ZN(O4275));
  INVX1 G45787 (.I(W1675), .ZN(O2613));
  INVX1 G45788 (.I(W27134), .ZN(O4299));
  INVX1 G45789 (.I(W1914), .ZN(W22772));
  INVX1 G45790 (.I(W3900), .ZN(W27969));
  INVX1 G45791 (.I(W7825), .ZN(O2610));
  INVX1 G45792 (.I(W6039), .ZN(O2611));
  INVX1 G45793 (.I(W13249), .ZN(O2612));
  INVX1 G45794 (.I(W19845), .ZN(W27964));
  INVX1 G45795 (.I(W3341), .ZN(W27963));
  INVX1 G45796 (.I(W8706), .ZN(W22779));
  INVX1 G45797 (.I(I344), .ZN(W22830));
  INVX1 G45798 (.I(W1565), .ZN(W22788));
  INVX1 G45799 (.I(W22454), .ZN(W22789));
  INVX1 G45800 (.I(W19529), .ZN(W22790));
  INVX1 G45801 (.I(W18275), .ZN(O2616));
  INVX1 G45802 (.I(W3605), .ZN(W27952));
  INVX1 G45803 (.I(W10145), .ZN(O4291));
  INVX1 G45804 (.I(W17711), .ZN(W27948));
  INVX1 G45805 (.I(W1833), .ZN(W27946));
  INVX1 G45806 (.I(W27810), .ZN(W27945));
  INVX1 G45807 (.I(W9545), .ZN(W27875));
  INVX1 G45808 (.I(W13705), .ZN(W27884));
  INVX1 G45809 (.I(W22587), .ZN(W22852));
  INVX1 G45810 (.I(W19496), .ZN(W27882));
  INVX1 G45811 (.I(W5264), .ZN(O4266));
  INVX1 G45812 (.I(W1369), .ZN(W22854));
  INVX1 G45813 (.I(W15601), .ZN(W27879));
  INVX1 G45814 (.I(W9495), .ZN(W27878));
  INVX1 G45815 (.I(W17953), .ZN(O4265));
  INVX1 G45816 (.I(I240), .ZN(W22855));
  INVX1 G45817 (.I(W12682), .ZN(W22851));
  INVX1 G45818 (.I(W11487), .ZN(O4263));
  INVX1 G45819 (.I(W14959), .ZN(W22860));
  INVX1 G45820 (.I(W3274), .ZN(W27870));
  INVX1 G45821 (.I(W15564), .ZN(W22866));
  INVX1 G45822 (.I(W13444), .ZN(W22868));
  INVX1 G45823 (.I(W3758), .ZN(W27865));
  INVX1 G45824 (.I(W1096), .ZN(O4259));
  INVX1 G45825 (.I(W957), .ZN(W22873));
  INVX1 G45826 (.I(W911), .ZN(O2624));
  INVX1 G45827 (.I(W18340), .ZN(W22839));
  INVX1 G45828 (.I(W18225), .ZN(W27910));
  INVX1 G45829 (.I(W4408), .ZN(O4274));
  INVX1 G45830 (.I(W15463), .ZN(W27907));
  INVX1 G45831 (.I(W19749), .ZN(W22835));
  INVX1 G45832 (.I(W7475), .ZN(W22836));
  INVX1 G45833 (.I(W11597), .ZN(O4271));
  INVX1 G45834 (.I(W23344), .ZN(W27901));
  INVX1 G45835 (.I(W4832), .ZN(O4270));
  INVX1 G45836 (.I(W12531), .ZN(O4269));
  INVX1 G45837 (.I(W6328), .ZN(W17911));
  INVX1 G45838 (.I(W20870), .ZN(W27896));
  INVX1 G45839 (.I(W5914), .ZN(W22843));
  INVX1 G45840 (.I(I1801), .ZN(O2620));
  INVX1 G45841 (.I(W11368), .ZN(W22845));
  INVX1 G45842 (.I(W4769), .ZN(W22848));
  INVX1 G45843 (.I(W5644), .ZN(W22849));
  INVX1 G45844 (.I(W24826), .ZN(O4267));
  INVX1 G45845 (.I(W21063), .ZN(W27887));
  INVX1 G45846 (.I(W15481), .ZN(W27886));
  INVX1 G45847 (.I(W27228), .ZN(W38143));
  INVX1 G45848 (.I(W7459), .ZN(W12677));
  INVX1 G45849 (.I(W12119), .ZN(W12679));
  INVX1 G45850 (.I(I347), .ZN(W38151));
  INVX1 G45851 (.I(W18680), .ZN(O9405));
  INVX1 G45852 (.I(W31592), .ZN(O9404));
  INVX1 G45853 (.I(W25507), .ZN(W38148));
  INVX1 G45854 (.I(W17558), .ZN(O9403));
  INVX1 G45855 (.I(W5575), .ZN(W12680));
  INVX1 G45856 (.I(W33696), .ZN(O9401));
  INVX1 G45857 (.I(W1407), .ZN(O9400));
  INVX1 G45858 (.I(W13619), .ZN(O9408));
  INVX1 G45859 (.I(W8469), .ZN(O634));
  INVX1 G45860 (.I(W8136), .ZN(O9398));
  INVX1 G45861 (.I(W36814), .ZN(O9397));
  INVX1 G45862 (.I(W25243), .ZN(W38137));
  INVX1 G45863 (.I(W26742), .ZN(W38136));
  INVX1 G45864 (.I(W4040), .ZN(O9396));
  INVX1 G45865 (.I(W14541), .ZN(W38133));
  INVX1 G45866 (.I(W1123), .ZN(O9395));
  INVX1 G45867 (.I(W16428), .ZN(W38130));
  INVX1 G45868 (.I(W9322), .ZN(W12663));
  INVX1 G45869 (.I(W1663), .ZN(W12643));
  INVX1 G45870 (.I(I156), .ZN(W38183));
  INVX1 G45871 (.I(W5437), .ZN(W12648));
  INVX1 G45872 (.I(W27353), .ZN(W38179));
  INVX1 G45873 (.I(W5293), .ZN(O9421));
  INVX1 G45874 (.I(W10930), .ZN(W12654));
  INVX1 G45875 (.I(W515), .ZN(W38174));
  INVX1 G45876 (.I(W10521), .ZN(W12660));
  INVX1 G45877 (.I(W18359), .ZN(O9417));
  INVX1 G45878 (.I(W20074), .ZN(O9394));
  INVX1 G45879 (.I(W11472), .ZN(W12665));
  INVX1 G45880 (.I(I386), .ZN(O9415));
  INVX1 G45881 (.I(W12054), .ZN(W12669));
  INVX1 G45882 (.I(W22053), .ZN(W38162));
  INVX1 G45883 (.I(W2164), .ZN(O9411));
  INVX1 G45884 (.I(W8026), .ZN(O631));
  INVX1 G45885 (.I(W36467), .ZN(O9409));
  INVX1 G45886 (.I(W7827), .ZN(O632));
  INVX1 G45887 (.I(W38151), .ZN(W38156));
  INVX1 G45888 (.I(I1149), .ZN(W12743));
  INVX1 G45889 (.I(W442), .ZN(W12730));
  INVX1 G45890 (.I(W10842), .ZN(O9367));
  INVX1 G45891 (.I(I687), .ZN(W38092));
  INVX1 G45892 (.I(W30722), .ZN(W38090));
  INVX1 G45893 (.I(W3433), .ZN(W12732));
  INVX1 G45894 (.I(I1865), .ZN(W12735));
  INVX1 G45895 (.I(W14822), .ZN(W38085));
  INVX1 G45896 (.I(W1433), .ZN(W12736));
  INVX1 G45897 (.I(W7618), .ZN(W12742));
  INVX1 G45898 (.I(W2982), .ZN(W12729));
  INVX1 G45899 (.I(W6779), .ZN(W12744));
  INVX1 G45900 (.I(W5684), .ZN(W12750));
  INVX1 G45901 (.I(W14655), .ZN(O9359));
  INVX1 G45902 (.I(W7641), .ZN(W12752));
  INVX1 G45903 (.I(W4333), .ZN(W12753));
  INVX1 G45904 (.I(W13168), .ZN(O9356));
  INVX1 G45905 (.I(W4305), .ZN(W12755));
  INVX1 G45906 (.I(W29883), .ZN(O9355));
  INVX1 G45907 (.I(W10107), .ZN(O9353));
  INVX1 G45908 (.I(W8757), .ZN(W12702));
  INVX1 G45909 (.I(W10024), .ZN(W12688));
  INVX1 G45910 (.I(W12628), .ZN(W12690));
  INVX1 G45911 (.I(W16361), .ZN(W38124));
  INVX1 G45912 (.I(W37952), .ZN(O9386));
  INVX1 G45913 (.I(W9873), .ZN(W12698));
  INVX1 G45914 (.I(W13556), .ZN(O9384));
  INVX1 G45915 (.I(W26156), .ZN(W38116));
  INVX1 G45916 (.I(W18055), .ZN(W38115));
  INVX1 G45917 (.I(W3344), .ZN(W12700));
  INVX1 G45918 (.I(W9874), .ZN(W12642));
  INVX1 G45919 (.I(W13723), .ZN(W38111));
  INVX1 G45920 (.I(W633), .ZN(W12709));
  INVX1 G45921 (.I(W27226), .ZN(W38108));
  INVX1 G45922 (.I(W11166), .ZN(W12713));
  INVX1 G45923 (.I(W4560), .ZN(O638));
  INVX1 G45924 (.I(W5095), .ZN(W12720));
  INVX1 G45925 (.I(W10929), .ZN(O639));
  INVX1 G45926 (.I(W1965), .ZN(O640));
  INVX1 G45927 (.I(I1472), .ZN(O641));
  INVX1 G45928 (.I(W10054), .ZN(O613));
  INVX1 G45929 (.I(W9109), .ZN(O9481));
  INVX1 G45930 (.I(W23255), .ZN(O9480));
  INVX1 G45931 (.I(W10277), .ZN(W12544));
  INVX1 G45932 (.I(W6692), .ZN(O609));
  INVX1 G45933 (.I(W1740), .ZN(W38281));
  INVX1 G45934 (.I(I1006), .ZN(W12548));
  INVX1 G45935 (.I(W1645), .ZN(O9476));
  INVX1 G45936 (.I(W34999), .ZN(O9473));
  INVX1 G45937 (.I(W4485), .ZN(W12562));
  INVX1 G45938 (.I(W10146), .ZN(W12563));
  INVX1 G45939 (.I(W11208), .ZN(W38287));
  INVX1 G45940 (.I(W14757), .ZN(O9468));
  INVX1 G45941 (.I(W6058), .ZN(O615));
  INVX1 G45942 (.I(I140), .ZN(W12570));
  INVX1 G45943 (.I(W8802), .ZN(W38259));
  INVX1 G45944 (.I(W1192), .ZN(W12571));
  INVX1 G45945 (.I(W10868), .ZN(O9465));
  INVX1 G45946 (.I(W26363), .ZN(W38256));
  INVX1 G45947 (.I(W741), .ZN(W12572));
  INVX1 G45948 (.I(W8325), .ZN(W12573));
  INVX1 G45949 (.I(W7224), .ZN(O9489));
  INVX1 G45950 (.I(W7924), .ZN(O9498));
  INVX1 G45951 (.I(W8339), .ZN(W12521));
  INVX1 G45952 (.I(W31121), .ZN(W38311));
  INVX1 G45953 (.I(W8018), .ZN(W12524));
  INVX1 G45954 (.I(W34765), .ZN(O9495));
  INVX1 G45955 (.I(W15454), .ZN(O9494));
  INVX1 G45956 (.I(W8112), .ZN(W12527));
  INVX1 G45957 (.I(W13716), .ZN(O9493));
  INVX1 G45958 (.I(W19016), .ZN(O9490));
  INVX1 G45959 (.I(W3460), .ZN(O617));
  INVX1 G45960 (.I(W4932), .ZN(W12534));
  INVX1 G45961 (.I(I1462), .ZN(W12537));
  INVX1 G45962 (.I(W27025), .ZN(O9487));
  INVX1 G45963 (.I(W7072), .ZN(W38294));
  INVX1 G45964 (.I(W15325), .ZN(O9486));
  INVX1 G45965 (.I(W3648), .ZN(W12539));
  INVX1 G45966 (.I(W4285), .ZN(W12540));
  INVX1 G45967 (.I(W9237), .ZN(O9482));
  INVX1 G45968 (.I(W601), .ZN(W12542));
  INVX1 G45969 (.I(W9719), .ZN(W12633));
  INVX1 G45970 (.I(W7420), .ZN(W12620));
  INVX1 G45971 (.I(I1617), .ZN(W12622));
  INVX1 G45972 (.I(I683), .ZN(W12623));
  INVX1 G45973 (.I(W21598), .ZN(O9435));
  INVX1 G45974 (.I(W22784), .ZN(W38207));
  INVX1 G45975 (.I(W21211), .ZN(W38206));
  INVX1 G45976 (.I(W3887), .ZN(W12625));
  INVX1 G45977 (.I(W21550), .ZN(W38203));
  INVX1 G45978 (.I(W12445), .ZN(W12630));
  INVX1 G45979 (.I(W578), .ZN(O623));
  INVX1 G45980 (.I(W12530), .ZN(W12634));
  INVX1 G45981 (.I(W11151), .ZN(W12636));
  INVX1 G45982 (.I(W4148), .ZN(W12637));
  INVX1 G45983 (.I(W24415), .ZN(W38195));
  INVX1 G45984 (.I(I1289), .ZN(O627));
  INVX1 G45985 (.I(W10626), .ZN(O9426));
  INVX1 G45986 (.I(W29057), .ZN(W38191));
  INVX1 G45987 (.I(I1340), .ZN(W12641));
  INVX1 G45988 (.I(W28315), .ZN(O9424));
  INVX1 G45989 (.I(W294), .ZN(W12592));
  INVX1 G45990 (.I(W31824), .ZN(O9461));
  INVX1 G45991 (.I(W17308), .ZN(O9459));
  INVX1 G45992 (.I(W9578), .ZN(W12581));
  INVX1 G45993 (.I(W24200), .ZN(O9456));
  INVX1 G45994 (.I(W9701), .ZN(O9455));
  INVX1 G45995 (.I(W10879), .ZN(W12583));
  INVX1 G45996 (.I(W1109), .ZN(O619));
  INVX1 G45997 (.I(W38074), .ZN(W38236));
  INVX1 G45998 (.I(W32318), .ZN(O9451));
  INVX1 G45999 (.I(W2802), .ZN(W12758));
  INVX1 G46000 (.I(W518), .ZN(W12593));
  INVX1 G46001 (.I(W9842), .ZN(O9448));
  INVX1 G46002 (.I(W2087), .ZN(W12602));
  INVX1 G46003 (.I(W665), .ZN(W12607));
  INVX1 G46004 (.I(W9315), .ZN(O9442));
  INVX1 G46005 (.I(W6392), .ZN(W12608));
  INVX1 G46006 (.I(W11025), .ZN(W12613));
  INVX1 G46007 (.I(W32093), .ZN(W38215));
  INVX1 G46008 (.I(W11922), .ZN(W12617));
  INVX1 G46009 (.I(I39), .ZN(W12932));
  INVX1 G46010 (.I(W6596), .ZN(W12913));
  INVX1 G46011 (.I(W3110), .ZN(W12914));
  INVX1 G46012 (.I(W3352), .ZN(W12915));
  INVX1 G46013 (.I(W5784), .ZN(W12921));
  INVX1 G46014 (.I(W20330), .ZN(O9264));
  INVX1 G46015 (.I(W6102), .ZN(W37898));
  INVX1 G46016 (.I(W547), .ZN(W12927));
  INVX1 G46017 (.I(W7862), .ZN(W12928));
  INVX1 G46018 (.I(W7180), .ZN(O9260));
  INVX1 G46019 (.I(W25653), .ZN(O9259));
  INVX1 G46020 (.I(W12274), .ZN(O9270));
  INVX1 G46021 (.I(W16762), .ZN(W37890));
  INVX1 G46022 (.I(W12735), .ZN(W12935));
  INVX1 G46023 (.I(W28299), .ZN(W37888));
  INVX1 G46024 (.I(I45), .ZN(O9257));
  INVX1 G46025 (.I(W6599), .ZN(O668));
  INVX1 G46026 (.I(W27455), .ZN(W37883));
  INVX1 G46027 (.I(W2460), .ZN(W12939));
  INVX1 G46028 (.I(I1259), .ZN(W12940));
  INVX1 G46029 (.I(W6703), .ZN(O670));
  INVX1 G46030 (.I(W22428), .ZN(O9279));
  INVX1 G46031 (.I(W7129), .ZN(W12897));
  INVX1 G46032 (.I(W3740), .ZN(O663));
  INVX1 G46033 (.I(W37888), .ZN(O9283));
  INVX1 G46034 (.I(W32408), .ZN(W37930));
  INVX1 G46035 (.I(W864), .ZN(W12900));
  INVX1 G46036 (.I(W13222), .ZN(W37928));
  INVX1 G46037 (.I(W17020), .ZN(O9282));
  INVX1 G46038 (.I(W15019), .ZN(W37925));
  INVX1 G46039 (.I(I1738), .ZN(O9281));
  INVX1 G46040 (.I(W11802), .ZN(W12945));
  INVX1 G46041 (.I(W937), .ZN(W12905));
  INVX1 G46042 (.I(W6004), .ZN(W37919));
  INVX1 G46043 (.I(W6959), .ZN(W12906));
  INVX1 G46044 (.I(W2153), .ZN(W12907));
  INVX1 G46045 (.I(W1874), .ZN(W12908));
  INVX1 G46046 (.I(W21666), .ZN(O9275));
  INVX1 G46047 (.I(W13410), .ZN(O9273));
  INVX1 G46048 (.I(W9385), .ZN(O9272));
  INVX1 G46049 (.I(W21779), .ZN(W37910));
  INVX1 G46050 (.I(W6572), .ZN(W12995));
  INVX1 G46051 (.I(W3898), .ZN(W12983));
  INVX1 G46052 (.I(W992), .ZN(W37850));
  INVX1 G46053 (.I(W7286), .ZN(W12984));
  INVX1 G46054 (.I(W6491), .ZN(O9231));
  INVX1 G46055 (.I(W17951), .ZN(O9230));
  INVX1 G46056 (.I(W34745), .ZN(O9229));
  INVX1 G46057 (.I(W9580), .ZN(O675));
  INVX1 G46058 (.I(W8343), .ZN(O676));
  INVX1 G46059 (.I(W9607), .ZN(W12992));
  INVX1 G46060 (.I(W32230), .ZN(O9235));
  INVX1 G46061 (.I(W3380), .ZN(W12999));
  INVX1 G46062 (.I(W33126), .ZN(O9221));
  INVX1 G46063 (.I(W3663), .ZN(W13003));
  INVX1 G46064 (.I(W1136), .ZN(O678));
  INVX1 G46065 (.I(W9748), .ZN(W13005));
  INVX1 G46066 (.I(W37527), .ZN(O9216));
  INVX1 G46067 (.I(W7690), .ZN(O9215));
  INVX1 G46068 (.I(W7116), .ZN(O679));
  INVX1 G46069 (.I(W8027), .ZN(W13012));
  INVX1 G46070 (.I(W32043), .ZN(O9241));
  INVX1 G46071 (.I(W30773), .ZN(W37877));
  INVX1 G46072 (.I(W17295), .ZN(O9248));
  INVX1 G46073 (.I(W3381), .ZN(W12949));
  INVX1 G46074 (.I(W2595), .ZN(W37873));
  INVX1 G46075 (.I(W11298), .ZN(W37872));
  INVX1 G46076 (.I(W11634), .ZN(W12964));
  INVX1 G46077 (.I(W27732), .ZN(O9244));
  INVX1 G46078 (.I(W32708), .ZN(O9243));
  INVX1 G46079 (.I(W11310), .ZN(W12966));
  INVX1 G46080 (.I(W29054), .ZN(W37935));
  INVX1 G46081 (.I(W22686), .ZN(W37863));
  INVX1 G46082 (.I(W11331), .ZN(W12969));
  INVX1 G46083 (.I(W3275), .ZN(W37861));
  INVX1 G46084 (.I(W12046), .ZN(W12970));
  INVX1 G46085 (.I(W4973), .ZN(W12973));
  INVX1 G46086 (.I(W12278), .ZN(O9238));
  INVX1 G46087 (.I(W3328), .ZN(W37857));
  INVX1 G46088 (.I(W2203), .ZN(W12976));
  INVX1 G46089 (.I(W17495), .ZN(O9237));
  INVX1 G46090 (.I(W10553), .ZN(W12816));
  INVX1 G46091 (.I(W3625), .ZN(W12798));
  INVX1 G46092 (.I(W4911), .ZN(O651));
  INVX1 G46093 (.I(W3922), .ZN(O653));
  INVX1 G46094 (.I(W6686), .ZN(W12809));
  INVX1 G46095 (.I(W4307), .ZN(O9329));
  INVX1 G46096 (.I(I1054), .ZN(W38018));
  INVX1 G46097 (.I(I1573), .ZN(O9328));
  INVX1 G46098 (.I(W2523), .ZN(W12812));
  INVX1 G46099 (.I(W37993), .ZN(W38014));
  INVX1 G46100 (.I(W12553), .ZN(W12794));
  INVX1 G46101 (.I(W13), .ZN(W38011));
  INVX1 G46102 (.I(W790), .ZN(O656));
  INVX1 G46103 (.I(W11076), .ZN(O9325));
  INVX1 G46104 (.I(W28413), .ZN(O9324));
  INVX1 G46105 (.I(W7076), .ZN(W12822));
  INVX1 G46106 (.I(W10355), .ZN(W12824));
  INVX1 G46107 (.I(W12451), .ZN(W12825));
  INVX1 G46108 (.I(W7289), .ZN(O9319));
  INVX1 G46109 (.I(W9231), .ZN(O9318));
  INVX1 G46110 (.I(W29663), .ZN(O9343));
  INVX1 G46111 (.I(W13700), .ZN(W38060));
  INVX1 G46112 (.I(W18309), .ZN(O9350));
  INVX1 G46113 (.I(I1678), .ZN(O9349));
  INVX1 G46114 (.I(W12613), .ZN(W12764));
  INVX1 G46115 (.I(W9645), .ZN(W12768));
  INVX1 G46116 (.I(W5597), .ZN(W12773));
  INVX1 G46117 (.I(W6205), .ZN(W12775));
  INVX1 G46118 (.I(W1436), .ZN(W12778));
  INVX1 G46119 (.I(W11727), .ZN(W12780));
  INVX1 G46120 (.I(W8143), .ZN(W37998));
  INVX1 G46121 (.I(W847), .ZN(W12783));
  INVX1 G46122 (.I(W9885), .ZN(O9342));
  INVX1 G46123 (.I(W10960), .ZN(O649));
  INVX1 G46124 (.I(W6172), .ZN(O9339));
  INVX1 G46125 (.I(W32692), .ZN(W38036));
  INVX1 G46126 (.I(W14), .ZN(W12788));
  INVX1 G46127 (.I(W15396), .ZN(W38031));
  INVX1 G46128 (.I(W5528), .ZN(W12792));
  INVX1 G46129 (.I(W353), .ZN(W38029));
  INVX1 G46130 (.I(W6378), .ZN(W12881));
  INVX1 G46131 (.I(W12738), .ZN(W12864));
  INVX1 G46132 (.I(W27740), .ZN(O9300));
  INVX1 G46133 (.I(W6037), .ZN(W12868));
  INVX1 G46134 (.I(I956), .ZN(W12871));
  INVX1 G46135 (.I(W22586), .ZN(W37960));
  INVX1 G46136 (.I(W9369), .ZN(W12874));
  INVX1 G46137 (.I(W5059), .ZN(O9295));
  INVX1 G46138 (.I(W23264), .ZN(W37954));
  INVX1 G46139 (.I(W11947), .ZN(W12880));
  INVX1 G46140 (.I(W12593), .ZN(W12857));
  INVX1 G46141 (.I(W24244), .ZN(W37950));
  INVX1 G46142 (.I(W10052), .ZN(O9291));
  INVX1 G46143 (.I(W4834), .ZN(W12885));
  INVX1 G46144 (.I(W26904), .ZN(W37945));
  INVX1 G46145 (.I(W7537), .ZN(W12886));
  INVX1 G46146 (.I(W3413), .ZN(W12889));
  INVX1 G46147 (.I(W585), .ZN(O9287));
  INVX1 G46148 (.I(W5618), .ZN(O662));
  INVX1 G46149 (.I(W21367), .ZN(O9286));
  INVX1 G46150 (.I(W14632), .ZN(O9307));
  INVX1 G46151 (.I(W19893), .ZN(W37993));
  INVX1 G46152 (.I(W11027), .ZN(O658));
  INVX1 G46153 (.I(W36205), .ZN(W37991));
  INVX1 G46154 (.I(W15150), .ZN(O9312));
  INVX1 G46155 (.I(W8061), .ZN(W12837));
  INVX1 G46156 (.I(W10154), .ZN(W12839));
  INVX1 G46157 (.I(W4757), .ZN(W12842));
  INVX1 G46158 (.I(W895), .ZN(W12843));
  INVX1 G46159 (.I(W10662), .ZN(O9308));
  INVX1 G46160 (.I(W28882), .ZN(W38315));
  INVX1 G46161 (.I(W25624), .ZN(W37982));
  INVX1 G46162 (.I(W7274), .ZN(O660));
  INVX1 G46163 (.I(W7143), .ZN(W37979));
  INVX1 G46164 (.I(W4755), .ZN(W12850));
  INVX1 G46165 (.I(W1436), .ZN(W37976));
  INVX1 G46166 (.I(I466), .ZN(W12852));
  INVX1 G46167 (.I(W5494), .ZN(W12853));
  INVX1 G46168 (.I(W16089), .ZN(O9302));
  INVX1 G46169 (.I(W24300), .ZN(W37971));
  INVX1 G46170 (.I(W4527), .ZN(O9685));
  INVX1 G46171 (.I(I5), .ZN(W38632));
  INVX1 G46172 (.I(W9352), .ZN(W12229));
  INVX1 G46173 (.I(W14655), .ZN(W38629));
  INVX1 G46174 (.I(W8607), .ZN(W12233));
  INVX1 G46175 (.I(W21032), .ZN(O9690));
  INVX1 G46176 (.I(W15823), .ZN(O9689));
  INVX1 G46177 (.I(I1663), .ZN(W12236));
  INVX1 G46178 (.I(I1703), .ZN(O582));
  INVX1 G46179 (.I(W4932), .ZN(W12241));
  INVX1 G46180 (.I(W38585), .ZN(O9686));
  INVX1 G46181 (.I(W12010), .ZN(W12228));
  INVX1 G46182 (.I(W12850), .ZN(O9684));
  INVX1 G46183 (.I(W15357), .ZN(O9683));
  INVX1 G46184 (.I(W10920), .ZN(O9681));
  INVX1 G46185 (.I(W7847), .ZN(W12245));
  INVX1 G46186 (.I(W25898), .ZN(O9679));
  INVX1 G46187 (.I(W4390), .ZN(W12249));
  INVX1 G46188 (.I(I140), .ZN(O9677));
  INVX1 G46189 (.I(W1563), .ZN(O584));
  INVX1 G46190 (.I(W13421), .ZN(W38605));
  INVX1 G46191 (.I(W33811), .ZN(O9706));
  INVX1 G46192 (.I(W29714), .ZN(O9714));
  INVX1 G46193 (.I(W3465), .ZN(W12205));
  INVX1 G46194 (.I(W32304), .ZN(O9712));
  INVX1 G46195 (.I(W18751), .ZN(O9711));
  INVX1 G46196 (.I(W13693), .ZN(O9710));
  INVX1 G46197 (.I(W25519), .ZN(O9709));
  INVX1 G46198 (.I(I822), .ZN(W38656));
  INVX1 G46199 (.I(W3926), .ZN(W12206));
  INVX1 G46200 (.I(W27014), .ZN(O9707));
  INVX1 G46201 (.I(W7873), .ZN(W12251));
  INVX1 G46202 (.I(W10953), .ZN(W12207));
  INVX1 G46203 (.I(W22785), .ZN(W38646));
  INVX1 G46204 (.I(W7175), .ZN(O9700));
  INVX1 G46205 (.I(W32887), .ZN(O9699));
  INVX1 G46206 (.I(W19488), .ZN(O9698));
  INVX1 G46207 (.I(W8001), .ZN(W12223));
  INVX1 G46208 (.I(I216), .ZN(O9696));
  INVX1 G46209 (.I(W6263), .ZN(W38638));
  INVX1 G46210 (.I(W20562), .ZN(W38637));
  INVX1 G46211 (.I(I1586), .ZN(W12305));
  INVX1 G46212 (.I(W7411), .ZN(W12290));
  INVX1 G46213 (.I(W22215), .ZN(W38562));
  INVX1 G46214 (.I(W4854), .ZN(W12297));
  INVX1 G46215 (.I(W17889), .ZN(O9651));
  INVX1 G46216 (.I(W17746), .ZN(W38557));
  INVX1 G46217 (.I(W37715), .ZN(W38555));
  INVX1 G46218 (.I(W10197), .ZN(W12302));
  INVX1 G46219 (.I(W10390), .ZN(O9648));
  INVX1 G46220 (.I(W10815), .ZN(W12303));
  INVX1 G46221 (.I(W754), .ZN(O9657));
  INVX1 G46222 (.I(I1540), .ZN(W12306));
  INVX1 G46223 (.I(W10298), .ZN(W12307));
  INVX1 G46224 (.I(W35591), .ZN(O9644));
  INVX1 G46225 (.I(W20540), .ZN(O9643));
  INVX1 G46226 (.I(W27753), .ZN(O9642));
  INVX1 G46227 (.I(W10661), .ZN(W38542));
  INVX1 G46228 (.I(W20856), .ZN(O9639));
  INVX1 G46229 (.I(W4811), .ZN(W12313));
  INVX1 G46230 (.I(W19122), .ZN(W38539));
  INVX1 G46231 (.I(W34264), .ZN(O9666));
  INVX1 G46232 (.I(W4694), .ZN(W12256));
  INVX1 G46233 (.I(W10225), .ZN(W12257));
  INVX1 G46234 (.I(W1160), .ZN(O585));
  INVX1 G46235 (.I(W2888), .ZN(W12268));
  INVX1 G46236 (.I(W37455), .ZN(W38592));
  INVX1 G46237 (.I(W5811), .ZN(W12269));
  INVX1 G46238 (.I(W9225), .ZN(W12271));
  INVX1 G46239 (.I(W37175), .ZN(W38587));
  INVX1 G46240 (.I(W15515), .ZN(O9667));
  INVX1 G46241 (.I(W6443), .ZN(W12203));
  INVX1 G46242 (.I(W16694), .ZN(O9665));
  INVX1 G46243 (.I(W28671), .ZN(W38582));
  INVX1 G46244 (.I(W6709), .ZN(W38581));
  INVX1 G46245 (.I(W7773), .ZN(O9664));
  INVX1 G46246 (.I(W23964), .ZN(W38576));
  INVX1 G46247 (.I(W33307), .ZN(O9662));
  INVX1 G46248 (.I(W32288), .ZN(W38572));
  INVX1 G46249 (.I(W7246), .ZN(W12283));
  INVX1 G46250 (.I(W2207), .ZN(O9658));
  INVX1 G46251 (.I(W8763), .ZN(W12106));
  INVX1 G46252 (.I(W11411), .ZN(W38756));
  INVX1 G46253 (.I(W9880), .ZN(W12094));
  INVX1 G46254 (.I(W3375), .ZN(W12095));
  INVX1 G46255 (.I(W2825), .ZN(O9767));
  INVX1 G46256 (.I(W12057), .ZN(W12098));
  INVX1 G46257 (.I(W19871), .ZN(W38750));
  INVX1 G46258 (.I(W2770), .ZN(W12099));
  INVX1 G46259 (.I(W8787), .ZN(O566));
  INVX1 G46260 (.I(W8783), .ZN(W38746));
  INVX1 G46261 (.I(W6701), .ZN(O9769));
  INVX1 G46262 (.I(W4697), .ZN(O9761));
  INVX1 G46263 (.I(W7125), .ZN(W12111));
  INVX1 G46264 (.I(W1362), .ZN(W12112));
  INVX1 G46265 (.I(W34205), .ZN(O9759));
  INVX1 G46266 (.I(W7079), .ZN(O9758));
  INVX1 G46267 (.I(W6113), .ZN(W12119));
  INVX1 G46268 (.I(W729), .ZN(W12121));
  INVX1 G46269 (.I(W8592), .ZN(O570));
  INVX1 G46270 (.I(W33423), .ZN(W38728));
  INVX1 G46271 (.I(W7107), .ZN(W12076));
  INVX1 G46272 (.I(W12148), .ZN(O9784));
  INVX1 G46273 (.I(W8021), .ZN(W12070));
  INVX1 G46274 (.I(W2666), .ZN(W38781));
  INVX1 G46275 (.I(W12175), .ZN(O9783));
  INVX1 G46276 (.I(W17574), .ZN(O9780));
  INVX1 G46277 (.I(W1775), .ZN(W12074));
  INVX1 G46278 (.I(W6594), .ZN(W12075));
  INVX1 G46279 (.I(I600), .ZN(W38774));
  INVX1 G46280 (.I(W8926), .ZN(O9778));
  INVX1 G46281 (.I(W5900), .ZN(W12129));
  INVX1 G46282 (.I(W622), .ZN(O9777));
  INVX1 G46283 (.I(W8765), .ZN(W12085));
  INVX1 G46284 (.I(I1848), .ZN(W12086));
  INVX1 G46285 (.I(W7043), .ZN(W12087));
  INVX1 G46286 (.I(W34878), .ZN(O9774));
  INVX1 G46287 (.I(W2822), .ZN(W12089));
  INVX1 G46288 (.I(W18425), .ZN(W38762));
  INVX1 G46289 (.I(W1621), .ZN(W12090));
  INVX1 G46290 (.I(W12508), .ZN(O9771));
  INVX1 G46291 (.I(W2657), .ZN(O575));
  INVX1 G46292 (.I(W8244), .ZN(O9736));
  INVX1 G46293 (.I(W18759), .ZN(W38694));
  INVX1 G46294 (.I(W4926), .ZN(W12170));
  INVX1 G46295 (.I(W5667), .ZN(W12173));
  INVX1 G46296 (.I(W573), .ZN(O9731));
  INVX1 G46297 (.I(W35420), .ZN(W38689));
  INVX1 G46298 (.I(W11111), .ZN(W12175));
  INVX1 G46299 (.I(W769), .ZN(W12180));
  INVX1 G46300 (.I(W2132), .ZN(W12181));
  INVX1 G46301 (.I(W11713), .ZN(W12163));
  INVX1 G46302 (.I(W429), .ZN(W12191));
  INVX1 G46303 (.I(W34775), .ZN(O9721));
  INVX1 G46304 (.I(W3938), .ZN(W12194));
  INVX1 G46305 (.I(W27279), .ZN(W38672));
  INVX1 G46306 (.I(W7990), .ZN(W12195));
  INVX1 G46307 (.I(W11301), .ZN(W12197));
  INVX1 G46308 (.I(W1549), .ZN(O9718));
  INVX1 G46309 (.I(W9055), .ZN(W12199));
  INVX1 G46310 (.I(W5145), .ZN(O577));
  INVX1 G46311 (.I(W1896), .ZN(W12142));
  INVX1 G46312 (.I(W7067), .ZN(W12130));
  INVX1 G46313 (.I(W7832), .ZN(W12131));
  INVX1 G46314 (.I(W7607), .ZN(W12132));
  INVX1 G46315 (.I(W35181), .ZN(O9750));
  INVX1 G46316 (.I(W1456), .ZN(W12133));
  INVX1 G46317 (.I(W12721), .ZN(W38721));
  INVX1 G46318 (.I(W7394), .ZN(W12134));
  INVX1 G46319 (.I(W7481), .ZN(W12135));
  INVX1 G46320 (.I(W7513), .ZN(W12136));
  INVX1 G46321 (.I(W25372), .ZN(O9638));
  INVX1 G46322 (.I(W6228), .ZN(W12149));
  INVX1 G46323 (.I(W8283), .ZN(W12150));
  INVX1 G46324 (.I(W10208), .ZN(W12151));
  INVX1 G46325 (.I(W38495), .ZN(W38711));
  INVX1 G46326 (.I(W1672), .ZN(W12152));
  INVX1 G46327 (.I(W4810), .ZN(W12155));
  INVX1 G46328 (.I(W9027), .ZN(W12156));
  INVX1 G46329 (.I(W31130), .ZN(W38704));
  INVX1 G46330 (.I(W2651), .ZN(W12162));
  INVX1 G46331 (.I(W29584), .ZN(O9545));
  INVX1 G46332 (.I(W32007), .ZN(O9554));
  INVX1 G46333 (.I(I704), .ZN(O9553));
  INVX1 G46334 (.I(W35947), .ZN(W38406));
  INVX1 G46335 (.I(W11206), .ZN(O9552));
  INVX1 G46336 (.I(W3452), .ZN(O9551));
  INVX1 G46337 (.I(W19539), .ZN(W38403));
  INVX1 G46338 (.I(W3656), .ZN(W12439));
  INVX1 G46339 (.I(W24161), .ZN(O9548));
  INVX1 G46340 (.I(W6252), .ZN(W12443));
  INVX1 G46341 (.I(W11148), .ZN(W12444));
  INVX1 G46342 (.I(W1011), .ZN(W12433));
  INVX1 G46343 (.I(W16533), .ZN(O9543));
  INVX1 G46344 (.I(W10105), .ZN(W12449));
  INVX1 G46345 (.I(W33446), .ZN(O9541));
  INVX1 G46346 (.I(W3905), .ZN(W12450));
  INVX1 G46347 (.I(W22657), .ZN(O9539));
  INVX1 G46348 (.I(W30953), .ZN(O9538));
  INVX1 G46349 (.I(W5277), .ZN(O9537));
  INVX1 G46350 (.I(W32957), .ZN(W38386));
  INVX1 G46351 (.I(W34298), .ZN(O9536));
  INVX1 G46352 (.I(W38315), .ZN(O9562));
  INVX1 G46353 (.I(W33572), .ZN(W38436));
  INVX1 G46354 (.I(W16874), .ZN(O9571));
  INVX1 G46355 (.I(W4100), .ZN(W12407));
  INVX1 G46356 (.I(W26342), .ZN(O9569));
  INVX1 G46357 (.I(W9447), .ZN(W12411));
  INVX1 G46358 (.I(W9890), .ZN(W12414));
  INVX1 G46359 (.I(W31312), .ZN(O9565));
  INVX1 G46360 (.I(W1259), .ZN(W12416));
  INVX1 G46361 (.I(W7052), .ZN(W12420));
  INVX1 G46362 (.I(W10212), .ZN(W12453));
  INVX1 G46363 (.I(W1696), .ZN(W12423));
  INVX1 G46364 (.I(W331), .ZN(W38421));
  INVX1 G46365 (.I(W29697), .ZN(O9559));
  INVX1 G46366 (.I(I988), .ZN(W12426));
  INVX1 G46367 (.I(W35222), .ZN(W38417));
  INVX1 G46368 (.I(W1740), .ZN(W38415));
  INVX1 G46369 (.I(W2106), .ZN(W12430));
  INVX1 G46370 (.I(W5729), .ZN(W12432));
  INVX1 G46371 (.I(W23102), .ZN(W38411));
  INVX1 G46372 (.I(W4750), .ZN(W12499));
  INVX1 G46373 (.I(W10770), .ZN(W12483));
  INVX1 G46374 (.I(W26238), .ZN(W38350));
  INVX1 G46375 (.I(W2343), .ZN(W12484));
  INVX1 G46376 (.I(W10372), .ZN(W38348));
  INVX1 G46377 (.I(W5071), .ZN(W12485));
  INVX1 G46378 (.I(W20689), .ZN(W38345));
  INVX1 G46379 (.I(W5761), .ZN(W12491));
  INVX1 G46380 (.I(W36282), .ZN(W38343));
  INVX1 G46381 (.I(W23399), .ZN(O9517));
  INVX1 G46382 (.I(W20857), .ZN(W38354));
  INVX1 G46383 (.I(W2594), .ZN(O9515));
  INVX1 G46384 (.I(W6992), .ZN(W12501));
  INVX1 G46385 (.I(W2507), .ZN(W12507));
  INVX1 G46386 (.I(W13209), .ZN(O9509));
  INVX1 G46387 (.I(W30146), .ZN(O9508));
  INVX1 G46388 (.I(W22569), .ZN(O9507));
  INVX1 G46389 (.I(W13364), .ZN(O9505));
  INVX1 G46390 (.I(W12403), .ZN(W12513));
  INVX1 G46391 (.I(W31179), .ZN(O9500));
  INVX1 G46392 (.I(W18768), .ZN(W38370));
  INVX1 G46393 (.I(W11874), .ZN(W12458));
  INVX1 G46394 (.I(W2592), .ZN(W38378));
  INVX1 G46395 (.I(W7109), .ZN(W12460));
  INVX1 G46396 (.I(I652), .ZN(O9532));
  INVX1 G46397 (.I(I464), .ZN(W12461));
  INVX1 G46398 (.I(W8226), .ZN(O602));
  INVX1 G46399 (.I(W7166), .ZN(W12463));
  INVX1 G46400 (.I(W24862), .ZN(O9530));
  INVX1 G46401 (.I(W35076), .ZN(W38371));
  INVX1 G46402 (.I(W9301), .ZN(O9576));
  INVX1 G46403 (.I(W8210), .ZN(W12466));
  INVX1 G46404 (.I(W4316), .ZN(W12468));
  INVX1 G46405 (.I(W23628), .ZN(O9527));
  INVX1 G46406 (.I(W1886), .ZN(W12471));
  INVX1 G46407 (.I(W28634), .ZN(O9524));
  INVX1 G46408 (.I(W36023), .ZN(W38362));
  INVX1 G46409 (.I(W5146), .ZN(W12474));
  INVX1 G46410 (.I(W1149), .ZN(O9523));
  INVX1 G46411 (.I(I1305), .ZN(W12479));
  INVX1 G46412 (.I(W17788), .ZN(O9613));
  INVX1 G46413 (.I(W5677), .ZN(W12347));
  INVX1 G46414 (.I(W13361), .ZN(O9619));
  INVX1 G46415 (.I(W7423), .ZN(W12351));
  INVX1 G46416 (.I(I676), .ZN(O9617));
  INVX1 G46417 (.I(W9015), .ZN(W38505));
  INVX1 G46418 (.I(W7946), .ZN(W12353));
  INVX1 G46419 (.I(W37020), .ZN(O9616));
  INVX1 G46420 (.I(W23890), .ZN(W38502));
  INVX1 G46421 (.I(W33227), .ZN(O9614));
  INVX1 G46422 (.I(W23843), .ZN(W38512));
  INVX1 G46423 (.I(W4260), .ZN(O9612));
  INVX1 G46424 (.I(W36452), .ZN(O9611));
  INVX1 G46425 (.I(W6461), .ZN(W12357));
  INVX1 G46426 (.I(W17419), .ZN(W38495));
  INVX1 G46427 (.I(W22072), .ZN(O9609));
  INVX1 G46428 (.I(W4159), .ZN(W12358));
  INVX1 G46429 (.I(W36926), .ZN(O9608));
  INVX1 G46430 (.I(I116), .ZN(W12359));
  INVX1 G46431 (.I(W9388), .ZN(W38490));
  INVX1 G46432 (.I(W535), .ZN(W12326));
  INVX1 G46433 (.I(W8407), .ZN(W12315));
  INVX1 G46434 (.I(W10228), .ZN(W12316));
  INVX1 G46435 (.I(W4779), .ZN(W38535));
  INVX1 G46436 (.I(W35382), .ZN(O9635));
  INVX1 G46437 (.I(W11759), .ZN(W12320));
  INVX1 G46438 (.I(I128), .ZN(W12322));
  INVX1 G46439 (.I(W2892), .ZN(W38529));
  INVX1 G46440 (.I(W8755), .ZN(W12323));
  INVX1 G46441 (.I(W5418), .ZN(W12324));
  INVX1 G46442 (.I(W2689), .ZN(O9607));
  INVX1 G46443 (.I(W3085), .ZN(W12327));
  INVX1 G46444 (.I(W3733), .ZN(W12330));
  INVX1 G46445 (.I(W13851), .ZN(O9628));
  INVX1 G46446 (.I(W922), .ZN(W12331));
  INVX1 G46447 (.I(W769), .ZN(O9626));
  INVX1 G46448 (.I(W32011), .ZN(O9624));
  INVX1 G46449 (.I(W5615), .ZN(O9623));
  INVX1 G46450 (.I(W22427), .ZN(O9622));
  INVX1 G46451 (.I(W5761), .ZN(W12342));
  INVX1 G46452 (.I(W14603), .ZN(O9585));
  INVX1 G46453 (.I(W7375), .ZN(W12379));
  INVX1 G46454 (.I(W5199), .ZN(W12381));
  INVX1 G46455 (.I(W32306), .ZN(O9592));
  INVX1 G46456 (.I(W7944), .ZN(O9591));
  INVX1 G46457 (.I(W5874), .ZN(O9590));
  INVX1 G46458 (.I(W20838), .ZN(O9588));
  INVX1 G46459 (.I(W2528), .ZN(O597));
  INVX1 G46460 (.I(W6998), .ZN(W12385));
  INVX1 G46461 (.I(W1713), .ZN(W12386));
  INVX1 G46462 (.I(W6118), .ZN(W38466));
  INVX1 G46463 (.I(W19443), .ZN(O9582));
  INVX1 G46464 (.I(W11687), .ZN(W12392));
  INVX1 G46465 (.I(W27803), .ZN(O9581));
  INVX1 G46466 (.I(W11217), .ZN(W12393));
  INVX1 G46467 (.I(W2261), .ZN(W12395));
  INVX1 G46468 (.I(W7173), .ZN(O9579));
  INVX1 G46469 (.I(W7082), .ZN(W12397));
  INVX1 G46470 (.I(W35984), .ZN(W38442));
  INVX1 G46471 (.I(W24500), .ZN(O9577));
  INVX1 G46472 (.I(W4329), .ZN(W12368));
  INVX1 G46473 (.I(W19865), .ZN(W38488));
  INVX1 G46474 (.I(W15207), .ZN(W38487));
  INVX1 G46475 (.I(I163), .ZN(O9605));
  INVX1 G46476 (.I(W9397), .ZN(W12361));
  INVX1 G46477 (.I(W5340), .ZN(W12362));
  INVX1 G46478 (.I(W13837), .ZN(W38482));
  INVX1 G46479 (.I(I831), .ZN(O9602));
  INVX1 G46480 (.I(W5959), .ZN(W12363));
  INVX1 G46481 (.I(W258), .ZN(W12365));
  INVX1 G46482 (.I(W4411), .ZN(W13013));
  INVX1 G46483 (.I(W33750), .ZN(O9599));
  INVX1 G46484 (.I(W3970), .ZN(W38475));
  INVX1 G46485 (.I(W8379), .ZN(W12369));
  INVX1 G46486 (.I(W33173), .ZN(O9598));
  INVX1 G46487 (.I(W9607), .ZN(W12374));
  INVX1 G46488 (.I(W9698), .ZN(W12377));
  INVX1 G46489 (.I(W2279), .ZN(W38469));
  INVX1 G46490 (.I(W17992), .ZN(W38468));
  INVX1 G46491 (.I(W1145), .ZN(O9595));
  INVX1 G46492 (.I(W12469), .ZN(W13686));
  INVX1 G46493 (.I(W2949), .ZN(W13675));
  INVX1 G46494 (.I(W10416), .ZN(O8812));
  INVX1 G46495 (.I(W34786), .ZN(W37156));
  INVX1 G46496 (.I(W21024), .ZN(O8811));
  INVX1 G46497 (.I(I940), .ZN(W13677));
  INVX1 G46498 (.I(W10899), .ZN(W13679));
  INVX1 G46499 (.I(W22615), .ZN(O8807));
  INVX1 G46500 (.I(W9126), .ZN(W13680));
  INVX1 G46501 (.I(I1764), .ZN(O775));
  INVX1 G46502 (.I(W26579), .ZN(O8806));
  INVX1 G46503 (.I(W20912), .ZN(O8814));
  INVX1 G46504 (.I(W3970), .ZN(W13688));
  INVX1 G46505 (.I(W12517), .ZN(W13696));
  INVX1 G46506 (.I(W9799), .ZN(W13697));
  INVX1 G46507 (.I(W166), .ZN(W37136));
  INVX1 G46508 (.I(W9868), .ZN(W13700));
  INVX1 G46509 (.I(W11819), .ZN(W13701));
  INVX1 G46510 (.I(W33916), .ZN(O8799));
  INVX1 G46511 (.I(W11154), .ZN(O778));
  INVX1 G46512 (.I(W13287), .ZN(W37128));
  INVX1 G46513 (.I(W471), .ZN(O771));
  INVX1 G46514 (.I(W1724), .ZN(W13641));
  INVX1 G46515 (.I(I240), .ZN(W13642));
  INVX1 G46516 (.I(W25418), .ZN(W37188));
  INVX1 G46517 (.I(W18512), .ZN(W37187));
  INVX1 G46518 (.I(W16019), .ZN(O8830));
  INVX1 G46519 (.I(W9116), .ZN(W13651));
  INVX1 G46520 (.I(W6325), .ZN(W13654));
  INVX1 G46521 (.I(W29988), .ZN(O8827));
  INVX1 G46522 (.I(W12826), .ZN(W13657));
  INVX1 G46523 (.I(W35666), .ZN(O8796));
  INVX1 G46524 (.I(W13635), .ZN(W13660));
  INVX1 G46525 (.I(W30888), .ZN(O8822));
  INVX1 G46526 (.I(W19025), .ZN(O8821));
  INVX1 G46527 (.I(W27102), .ZN(W37170));
  INVX1 G46528 (.I(W18162), .ZN(O8818));
  INVX1 G46529 (.I(W19107), .ZN(O8816));
  INVX1 G46530 (.I(W10004), .ZN(W13666));
  INVX1 G46531 (.I(W7278), .ZN(W13673));
  INVX1 G46532 (.I(W26878), .ZN(W37161));
  INVX1 G46533 (.I(W32119), .ZN(O8771));
  INVX1 G46534 (.I(W4918), .ZN(W13734));
  INVX1 G46535 (.I(W8573), .ZN(W13738));
  INVX1 G46536 (.I(W7916), .ZN(O8778));
  INVX1 G46537 (.I(W15528), .ZN(W37096));
  INVX1 G46538 (.I(I1428), .ZN(O8777));
  INVX1 G46539 (.I(W14553), .ZN(O8776));
  INVX1 G46540 (.I(W31572), .ZN(W37090));
  INVX1 G46541 (.I(W35539), .ZN(O8773));
  INVX1 G46542 (.I(W4702), .ZN(W13744));
  INVX1 G46543 (.I(W3393), .ZN(O8781));
  INVX1 G46544 (.I(W7502), .ZN(W13745));
  INVX1 G46545 (.I(W264), .ZN(W13748));
  INVX1 G46546 (.I(W4216), .ZN(W13749));
  INVX1 G46547 (.I(W5072), .ZN(W13752));
  INVX1 G46548 (.I(W4399), .ZN(W37081));
  INVX1 G46549 (.I(W32598), .ZN(W37080));
  INVX1 G46550 (.I(W6764), .ZN(O8765));
  INVX1 G46551 (.I(W540), .ZN(W13754));
  INVX1 G46552 (.I(W145), .ZN(W13755));
  INVX1 G46553 (.I(W7239), .ZN(O8786));
  INVX1 G46554 (.I(W11083), .ZN(W13709));
  INVX1 G46555 (.I(I1708), .ZN(W13710));
  INVX1 G46556 (.I(W9733), .ZN(W13716));
  INVX1 G46557 (.I(W11342), .ZN(O8792));
  INVX1 G46558 (.I(W3395), .ZN(W13719));
  INVX1 G46559 (.I(W6389), .ZN(W13720));
  INVX1 G46560 (.I(W13616), .ZN(W13721));
  INVX1 G46561 (.I(W2475), .ZN(W13724));
  INVX1 G46562 (.I(W9787), .ZN(O8787));
  INVX1 G46563 (.I(W4238), .ZN(W13640));
  INVX1 G46564 (.I(W5644), .ZN(W13728));
  INVX1 G46565 (.I(W35522), .ZN(W37110));
  INVX1 G46566 (.I(W20280), .ZN(W37109));
  INVX1 G46567 (.I(W22813), .ZN(O8785));
  INVX1 G46568 (.I(I938), .ZN(W37107));
  INVX1 G46569 (.I(W10946), .ZN(W13729));
  INVX1 G46570 (.I(W11358), .ZN(O8784));
  INVX1 G46571 (.I(W23359), .ZN(O8783));
  INVX1 G46572 (.I(W12829), .ZN(O779));
  INVX1 G46573 (.I(W18486), .ZN(O8877));
  INVX1 G46574 (.I(W5550), .ZN(W13542));
  INVX1 G46575 (.I(W7803), .ZN(O8889));
  INVX1 G46576 (.I(W15315), .ZN(O8888));
  INVX1 G46577 (.I(W1717), .ZN(W37281));
  INVX1 G46578 (.I(W10995), .ZN(W13548));
  INVX1 G46579 (.I(W6549), .ZN(O756));
  INVX1 G46580 (.I(W21209), .ZN(O8884));
  INVX1 G46581 (.I(W22032), .ZN(O8883));
  INVX1 G46582 (.I(W5106), .ZN(O8880));
  INVX1 G46583 (.I(W5297), .ZN(O8890));
  INVX1 G46584 (.I(W5736), .ZN(W13566));
  INVX1 G46585 (.I(W26665), .ZN(W37267));
  INVX1 G46586 (.I(W6632), .ZN(O8875));
  INVX1 G46587 (.I(W5013), .ZN(W13574));
  INVX1 G46588 (.I(W2296), .ZN(W37262));
  INVX1 G46589 (.I(I638), .ZN(W13576));
  INVX1 G46590 (.I(W10657), .ZN(O760));
  INVX1 G46591 (.I(W3783), .ZN(W13578));
  INVX1 G46592 (.I(W11478), .ZN(W13580));
  INVX1 G46593 (.I(W4358), .ZN(W13530));
  INVX1 G46594 (.I(W33716), .ZN(O8911));
  INVX1 G46595 (.I(W8009), .ZN(O8909));
  INVX1 G46596 (.I(W11242), .ZN(W13518));
  INVX1 G46597 (.I(W3711), .ZN(W13521));
  INVX1 G46598 (.I(W10349), .ZN(W37312));
  INVX1 G46599 (.I(W7912), .ZN(O752));
  INVX1 G46600 (.I(W1616), .ZN(W13523));
  INVX1 G46601 (.I(W12520), .ZN(W13526));
  INVX1 G46602 (.I(W6012), .ZN(W13528));
  INVX1 G46603 (.I(W3376), .ZN(O761));
  INVX1 G46604 (.I(W18856), .ZN(O8901));
  INVX1 G46605 (.I(I1391), .ZN(O8899));
  INVX1 G46606 (.I(W34936), .ZN(O8897));
  INVX1 G46607 (.I(W33516), .ZN(O8896));
  INVX1 G46608 (.I(I920), .ZN(W13535));
  INVX1 G46609 (.I(W7712), .ZN(W13536));
  INVX1 G46610 (.I(W12446), .ZN(W13539));
  INVX1 G46611 (.I(I1180), .ZN(O8894));
  INVX1 G46612 (.I(W34761), .ZN(O8892));
  INVX1 G46613 (.I(W22136), .ZN(O8842));
  INVX1 G46614 (.I(W4855), .ZN(W37219));
  INVX1 G46615 (.I(W6992), .ZN(W37217));
  INVX1 G46616 (.I(W1322), .ZN(W13619));
  INVX1 G46617 (.I(I1799), .ZN(W13623));
  INVX1 G46618 (.I(W5310), .ZN(W37212));
  INVX1 G46619 (.I(W15011), .ZN(O8845));
  INVX1 G46620 (.I(W8356), .ZN(W37210));
  INVX1 G46621 (.I(I537), .ZN(W13630));
  INVX1 G46622 (.I(I638), .ZN(W13631));
  INVX1 G46623 (.I(W13050), .ZN(W13617));
  INVX1 G46624 (.I(W4875), .ZN(O8841));
  INVX1 G46625 (.I(W32583), .ZN(O8839));
  INVX1 G46626 (.I(W29769), .ZN(O8838));
  INVX1 G46627 (.I(I32), .ZN(W13633));
  INVX1 G46628 (.I(W5140), .ZN(W37199));
  INVX1 G46629 (.I(W9551), .ZN(O767));
  INVX1 G46630 (.I(W29751), .ZN(W37196));
  INVX1 G46631 (.I(W1320), .ZN(W13637));
  INVX1 G46632 (.I(W12450), .ZN(O8835));
  INVX1 G46633 (.I(W19050), .ZN(O8858));
  INVX1 G46634 (.I(W10821), .ZN(W37251));
  INVX1 G46635 (.I(W4655), .ZN(W13587));
  INVX1 G46636 (.I(W33839), .ZN(W37248));
  INVX1 G46637 (.I(I1406), .ZN(W13589));
  INVX1 G46638 (.I(W7862), .ZN(O762));
  INVX1 G46639 (.I(W7779), .ZN(W13594));
  INVX1 G46640 (.I(W7070), .ZN(O8867));
  INVX1 G46641 (.I(W3436), .ZN(O8863));
  INVX1 G46642 (.I(W5909), .ZN(W13599));
  INVX1 G46643 (.I(W22911), .ZN(W37076));
  INVX1 G46644 (.I(I1267), .ZN(W13604));
  INVX1 G46645 (.I(W2019), .ZN(W13606));
  INVX1 G46646 (.I(W12732), .ZN(W13610));
  INVX1 G46647 (.I(W5627), .ZN(O8855));
  INVX1 G46648 (.I(I1336), .ZN(O8854));
  INVX1 G46649 (.I(W30810), .ZN(O8853));
  INVX1 G46650 (.I(W31034), .ZN(O8852));
  INVX1 G46651 (.I(W18202), .ZN(W37226));
  INVX1 G46652 (.I(W13588), .ZN(W37222));
  INVX1 G46653 (.I(W36355), .ZN(O8681));
  INVX1 G46654 (.I(W728), .ZN(W36941));
  INVX1 G46655 (.I(I401), .ZN(W13881));
  INVX1 G46656 (.I(W12254), .ZN(W13883));
  INVX1 G46657 (.I(W6021), .ZN(W13887));
  INVX1 G46658 (.I(W23852), .ZN(O8685));
  INVX1 G46659 (.I(W6994), .ZN(O8684));
  INVX1 G46660 (.I(W12882), .ZN(W13888));
  INVX1 G46661 (.I(W11828), .ZN(W13890));
  INVX1 G46662 (.I(W4460), .ZN(W13892));
  INVX1 G46663 (.I(W22449), .ZN(W36929));
  INVX1 G46664 (.I(W14750), .ZN(O8690));
  INVX1 G46665 (.I(W33653), .ZN(O8680));
  INVX1 G46666 (.I(W1731), .ZN(W13897));
  INVX1 G46667 (.I(W23669), .ZN(O8679));
  INVX1 G46668 (.I(W17641), .ZN(O8678));
  INVX1 G46669 (.I(W830), .ZN(O8677));
  INVX1 G46670 (.I(W12042), .ZN(O800));
  INVX1 G46671 (.I(W26308), .ZN(W36921));
  INVX1 G46672 (.I(W1147), .ZN(O801));
  INVX1 G46673 (.I(W21789), .ZN(O8674));
  INVX1 G46674 (.I(W31091), .ZN(W36952));
  INVX1 G46675 (.I(W5252), .ZN(W36965));
  INVX1 G46676 (.I(W21218), .ZN(O8703));
  INVX1 G46677 (.I(W10974), .ZN(W13871));
  INVX1 G46678 (.I(W30733), .ZN(W36962));
  INVX1 G46679 (.I(W25311), .ZN(O8701));
  INVX1 G46680 (.I(W25268), .ZN(O8700));
  INVX1 G46681 (.I(W22822), .ZN(W36956));
  INVX1 G46682 (.I(W2875), .ZN(W13876));
  INVX1 G46683 (.I(W8171), .ZN(W36953));
  INVX1 G46684 (.I(W20878), .ZN(O8673));
  INVX1 G46685 (.I(W29286), .ZN(O8696));
  INVX1 G46686 (.I(W27594), .ZN(W36950));
  INVX1 G46687 (.I(W1389), .ZN(O8695));
  INVX1 G46688 (.I(W27357), .ZN(O8694));
  INVX1 G46689 (.I(W21064), .ZN(O8693));
  INVX1 G46690 (.I(W9337), .ZN(W13878));
  INVX1 G46691 (.I(W8857), .ZN(W36945));
  INVX1 G46692 (.I(W12223), .ZN(W36944));
  INVX1 G46693 (.I(W33411), .ZN(O8691));
  INVX1 G46694 (.I(W2942), .ZN(W13944));
  INVX1 G46695 (.I(W19917), .ZN(O8654));
  INVX1 G46696 (.I(W8508), .ZN(O8652));
  INVX1 G46697 (.I(W8138), .ZN(W13930));
  INVX1 G46698 (.I(W6631), .ZN(O8651));
  INVX1 G46699 (.I(W1197), .ZN(O806));
  INVX1 G46700 (.I(W1837), .ZN(W13939));
  INVX1 G46701 (.I(W1723), .ZN(O8648));
  INVX1 G46702 (.I(W21793), .ZN(W36878));
  INVX1 G46703 (.I(W19362), .ZN(W36877));
  INVX1 G46704 (.I(W11019), .ZN(W13927));
  INVX1 G46705 (.I(W16696), .ZN(W36873));
  INVX1 G46706 (.I(W36789), .ZN(W36870));
  INVX1 G46707 (.I(W26585), .ZN(W36869));
  INVX1 G46708 (.I(W593), .ZN(W13948));
  INVX1 G46709 (.I(W15625), .ZN(W36867));
  INVX1 G46710 (.I(W36806), .ZN(O8642));
  INVX1 G46711 (.I(W1053), .ZN(O8641));
  INVX1 G46712 (.I(W1304), .ZN(W13949));
  INVX1 G46713 (.I(W12547), .ZN(W36861));
  INVX1 G46714 (.I(W5244), .ZN(O8666));
  INVX1 G46715 (.I(W6654), .ZN(W13905));
  INVX1 G46716 (.I(W13657), .ZN(W13907));
  INVX1 G46717 (.I(W24334), .ZN(W36914));
  INVX1 G46718 (.I(W7329), .ZN(O802));
  INVX1 G46719 (.I(W10590), .ZN(O803));
  INVX1 G46720 (.I(W32659), .ZN(W36910));
  INVX1 G46721 (.I(W650), .ZN(W13911));
  INVX1 G46722 (.I(W166), .ZN(O804));
  INVX1 G46723 (.I(W9515), .ZN(W13913));
  INVX1 G46724 (.I(W9769), .ZN(W13869));
  INVX1 G46725 (.I(W3328), .ZN(W13914));
  INVX1 G46726 (.I(W28839), .ZN(O8664));
  INVX1 G46727 (.I(W14147), .ZN(W36903));
  INVX1 G46728 (.I(W23674), .ZN(O8663));
  INVX1 G46729 (.I(W33803), .ZN(O8662));
  INVX1 G46730 (.I(W11897), .ZN(W36900));
  INVX1 G46731 (.I(W12928), .ZN(W13916));
  INVX1 G46732 (.I(I1807), .ZN(O805));
  INVX1 G46733 (.I(W29012), .ZN(O8656));
  INVX1 G46734 (.I(W6453), .ZN(W13797));
  INVX1 G46735 (.I(W30350), .ZN(O8745));
  INVX1 G46736 (.I(W19165), .ZN(O8744));
  INVX1 G46737 (.I(W206), .ZN(W13781));
  INVX1 G46738 (.I(W5387), .ZN(W13783));
  INVX1 G46739 (.I(W6520), .ZN(W13785));
  INVX1 G46740 (.I(W337), .ZN(W13788));
  INVX1 G46741 (.I(W1324), .ZN(W13790));
  INVX1 G46742 (.I(W3167), .ZN(O786));
  INVX1 G46743 (.I(I1969), .ZN(O8739));
  INVX1 G46744 (.I(W3566), .ZN(W13780));
  INVX1 G46745 (.I(W3300), .ZN(W37036));
  INVX1 G46746 (.I(W10620), .ZN(W13798));
  INVX1 G46747 (.I(I1310), .ZN(O8738));
  INVX1 G46748 (.I(W32186), .ZN(O8737));
  INVX1 G46749 (.I(W541), .ZN(W13802));
  INVX1 G46750 (.I(W9661), .ZN(W13804));
  INVX1 G46751 (.I(W9670), .ZN(O8734));
  INVX1 G46752 (.I(W21930), .ZN(W37029));
  INVX1 G46753 (.I(W8844), .ZN(W37028));
  INVX1 G46754 (.I(W27692), .ZN(O8756));
  INVX1 G46755 (.I(W34400), .ZN(O8762));
  INVX1 G46756 (.I(W18545), .ZN(O8761));
  INVX1 G46757 (.I(W1372), .ZN(W13760));
  INVX1 G46758 (.I(W17423), .ZN(W37070));
  INVX1 G46759 (.I(W14805), .ZN(O8760));
  INVX1 G46760 (.I(W4535), .ZN(W13763));
  INVX1 G46761 (.I(W1329), .ZN(W13764));
  INVX1 G46762 (.I(W2169), .ZN(W13765));
  INVX1 G46763 (.I(W13482), .ZN(W13766));
  INVX1 G46764 (.I(W19350), .ZN(W37027));
  INVX1 G46765 (.I(W7677), .ZN(W37063));
  INVX1 G46766 (.I(W7956), .ZN(O8755));
  INVX1 G46767 (.I(W23627), .ZN(O8754));
  INVX1 G46768 (.I(W4086), .ZN(W13768));
  INVX1 G46769 (.I(W12897), .ZN(W13773));
  INVX1 G46770 (.I(W17536), .ZN(W37055));
  INVX1 G46771 (.I(W10232), .ZN(W13775));
  INVX1 G46772 (.I(W193), .ZN(O8749));
  INVX1 G46773 (.I(W33920), .ZN(O8748));
  INVX1 G46774 (.I(W11515), .ZN(O8716));
  INVX1 G46775 (.I(W35482), .ZN(W36999));
  INVX1 G46776 (.I(W32491), .ZN(O8724));
  INVX1 G46777 (.I(W12945), .ZN(W13837));
  INVX1 G46778 (.I(W25480), .ZN(W36996));
  INVX1 G46779 (.I(W10866), .ZN(W13839));
  INVX1 G46780 (.I(W23680), .ZN(O8721));
  INVX1 G46781 (.I(W12251), .ZN(W13841));
  INVX1 G46782 (.I(I1373), .ZN(O789));
  INVX1 G46783 (.I(W7220), .ZN(O790));
  INVX1 G46784 (.I(W230), .ZN(W13836));
  INVX1 G46785 (.I(W2098), .ZN(W36983));
  INVX1 G46786 (.I(W31439), .ZN(W36982));
  INVX1 G46787 (.I(W11521), .ZN(W13852));
  INVX1 G46788 (.I(W22161), .ZN(O8712));
  INVX1 G46789 (.I(W22099), .ZN(W36978));
  INVX1 G46790 (.I(W8752), .ZN(W13854));
  INVX1 G46791 (.I(W11968), .ZN(W36975));
  INVX1 G46792 (.I(W1600), .ZN(W13858));
  INVX1 G46793 (.I(W12890), .ZN(O794));
  INVX1 G46794 (.I(W20447), .ZN(W37015));
  INVX1 G46795 (.I(W1470), .ZN(O8733));
  INVX1 G46796 (.I(W141), .ZN(W13805));
  INVX1 G46797 (.I(W5218), .ZN(W13807));
  INVX1 G46798 (.I(W2811), .ZN(W13808));
  INVX1 G46799 (.I(W7669), .ZN(W13809));
  INVX1 G46800 (.I(W5243), .ZN(W37021));
  INVX1 G46801 (.I(W12081), .ZN(W37020));
  INVX1 G46802 (.I(W1048), .ZN(W13810));
  INVX1 G46803 (.I(W13337), .ZN(W13815));
  INVX1 G46804 (.I(W17113), .ZN(O8912));
  INVX1 G46805 (.I(W13625), .ZN(O8730));
  INVX1 G46806 (.I(W7907), .ZN(W13817));
  INVX1 G46807 (.I(W12916), .ZN(W37012));
  INVX1 G46808 (.I(W8372), .ZN(W37011));
  INVX1 G46809 (.I(W7130), .ZN(W13822));
  INVX1 G46810 (.I(W2045), .ZN(W13825));
  INVX1 G46811 (.I(W32763), .ZN(W37005));
  INVX1 G46812 (.I(W1361), .ZN(W13833));
  INVX1 G46813 (.I(I1606), .ZN(W13834));
  INVX1 G46814 (.I(W23312), .ZN(O9102));
  INVX1 G46815 (.I(W18767), .ZN(O9114));
  INVX1 G46816 (.I(W7435), .ZN(W13162));
  INVX1 G46817 (.I(W23834), .ZN(O9112));
  INVX1 G46818 (.I(W6920), .ZN(W13163));
  INVX1 G46819 (.I(W39), .ZN(O9110));
  INVX1 G46820 (.I(W10154), .ZN(W13164));
  INVX1 G46821 (.I(W1659), .ZN(O704));
  INVX1 G46822 (.I(W33147), .ZN(O9107));
  INVX1 G46823 (.I(W9838), .ZN(W13169));
  INVX1 G46824 (.I(W282), .ZN(W13172));
  INVX1 G46825 (.I(W26239), .ZN(O9116));
  INVX1 G46826 (.I(W25239), .ZN(W37653));
  INVX1 G46827 (.I(W3905), .ZN(W13175));
  INVX1 G46828 (.I(W5672), .ZN(O706));
  INVX1 G46829 (.I(W36892), .ZN(W37648));
  INVX1 G46830 (.I(W17226), .ZN(W37645));
  INVX1 G46831 (.I(W9384), .ZN(O707));
  INVX1 G46832 (.I(I1361), .ZN(W37643));
  INVX1 G46833 (.I(W9342), .ZN(W13183));
  INVX1 G46834 (.I(W30622), .ZN(O9096));
  INVX1 G46835 (.I(W31288), .ZN(O9125));
  INVX1 G46836 (.I(W11618), .ZN(O701));
  INVX1 G46837 (.I(W1513), .ZN(O9133));
  INVX1 G46838 (.I(W679), .ZN(W13139));
  INVX1 G46839 (.I(W9272), .ZN(W13140));
  INVX1 G46840 (.I(W26025), .ZN(O9131));
  INVX1 G46841 (.I(W9164), .ZN(W13142));
  INVX1 G46842 (.I(W20466), .ZN(O9129));
  INVX1 G46843 (.I(W4998), .ZN(W13145));
  INVX1 G46844 (.I(W5505), .ZN(O702));
  INVX1 G46845 (.I(I1430), .ZN(W13186));
  INVX1 G46846 (.I(W12481), .ZN(W13151));
  INVX1 G46847 (.I(W9070), .ZN(W13153));
  INVX1 G46848 (.I(W33584), .ZN(O9123));
  INVX1 G46849 (.I(W24009), .ZN(O9122));
  INVX1 G46850 (.I(W8211), .ZN(W13158));
  INVX1 G46851 (.I(W7643), .ZN(O9120));
  INVX1 G46852 (.I(I415), .ZN(W13159));
  INVX1 G46853 (.I(W4888), .ZN(W13160));
  INVX1 G46854 (.I(W9404), .ZN(O9117));
  INVX1 G46855 (.I(W12830), .ZN(W13254));
  INVX1 G46856 (.I(W27303), .ZN(W37601));
  INVX1 G46857 (.I(W10748), .ZN(W13231));
  INVX1 G46858 (.I(W22848), .ZN(W37599));
  INVX1 G46859 (.I(I197), .ZN(O715));
  INVX1 G46860 (.I(W4897), .ZN(W13239));
  INVX1 G46861 (.I(I1853), .ZN(W13247));
  INVX1 G46862 (.I(W5306), .ZN(W37590));
  INVX1 G46863 (.I(W3779), .ZN(O718));
  INVX1 G46864 (.I(W11258), .ZN(W13253));
  INVX1 G46865 (.I(W34622), .ZN(W37603));
  INVX1 G46866 (.I(W16914), .ZN(W37583));
  INVX1 G46867 (.I(W30864), .ZN(W37582));
  INVX1 G46868 (.I(W16974), .ZN(O9063));
  INVX1 G46869 (.I(W2641), .ZN(W37577));
  INVX1 G46870 (.I(W22223), .ZN(O9060));
  INVX1 G46871 (.I(W28627), .ZN(W37575));
  INVX1 G46872 (.I(W14286), .ZN(W37570));
  INVX1 G46873 (.I(W6428), .ZN(W13271));
  INVX1 G46874 (.I(W31205), .ZN(O9056));
  INVX1 G46875 (.I(I764), .ZN(W13212));
  INVX1 G46876 (.I(W14298), .ZN(W37638));
  INVX1 G46877 (.I(W17730), .ZN(W37637));
  INVX1 G46878 (.I(W12747), .ZN(W13191));
  INVX1 G46879 (.I(W24959), .ZN(O9093));
  INVX1 G46880 (.I(W11182), .ZN(O709));
  INVX1 G46881 (.I(W14554), .ZN(O9087));
  INVX1 G46882 (.I(W3307), .ZN(O710));
  INVX1 G46883 (.I(W4988), .ZN(O711));
  INVX1 G46884 (.I(W4651), .ZN(W37620));
  INVX1 G46885 (.I(W25165), .ZN(O9135));
  INVX1 G46886 (.I(W11342), .ZN(W13214));
  INVX1 G46887 (.I(W5486), .ZN(W13218));
  INVX1 G46888 (.I(W34679), .ZN(O9078));
  INVX1 G46889 (.I(W2798), .ZN(W13221));
  INVX1 G46890 (.I(W20223), .ZN(W37609));
  INVX1 G46891 (.I(W8967), .ZN(W13226));
  INVX1 G46892 (.I(W32599), .ZN(W37607));
  INVX1 G46893 (.I(W22730), .ZN(O9075));
  INVX1 G46894 (.I(W36576), .ZN(O9074));
  INVX1 G46895 (.I(I639), .ZN(O690));
  INVX1 G46896 (.I(W31576), .ZN(W37783));
  INVX1 G46897 (.I(W32132), .ZN(O9184));
  INVX1 G46898 (.I(W16501), .ZN(W37781));
  INVX1 G46899 (.I(W2877), .ZN(W13060));
  INVX1 G46900 (.I(I1504), .ZN(W13063));
  INVX1 G46901 (.I(W427), .ZN(W13066));
  INVX1 G46902 (.I(W10684), .ZN(O9179));
  INVX1 G46903 (.I(W5294), .ZN(W13073));
  INVX1 G46904 (.I(W31367), .ZN(O9176));
  INVX1 G46905 (.I(W6063), .ZN(W13056));
  INVX1 G46906 (.I(W901), .ZN(O9175));
  INVX1 G46907 (.I(W25179), .ZN(O9174));
  INVX1 G46908 (.I(W33045), .ZN(W37763));
  INVX1 G46909 (.I(W26582), .ZN(W37761));
  INVX1 G46910 (.I(W32862), .ZN(O9172));
  INVX1 G46911 (.I(W31937), .ZN(O9171));
  INVX1 G46912 (.I(W6187), .ZN(W37758));
  INVX1 G46913 (.I(W4912), .ZN(W13078));
  INVX1 G46914 (.I(W12839), .ZN(W37755));
  INVX1 G46915 (.I(W29141), .ZN(W37812));
  INVX1 G46916 (.I(W2922), .ZN(W13016));
  INVX1 G46917 (.I(W7031), .ZN(W13018));
  INVX1 G46918 (.I(W3247), .ZN(W13020));
  INVX1 G46919 (.I(W13101), .ZN(O9210));
  INVX1 G46920 (.I(W28708), .ZN(O9209));
  INVX1 G46921 (.I(W10478), .ZN(O9208));
  INVX1 G46922 (.I(W29445), .ZN(W37815));
  INVX1 G46923 (.I(W24090), .ZN(O9206));
  INVX1 G46924 (.I(W4340), .ZN(O9205));
  INVX1 G46925 (.I(W37278), .ZN(O9167));
  INVX1 G46926 (.I(W29680), .ZN(O9204));
  INVX1 G46927 (.I(W5321), .ZN(W13023));
  INVX1 G46928 (.I(W22328), .ZN(O9201));
  INVX1 G46929 (.I(W8167), .ZN(W13034));
  INVX1 G46930 (.I(W9238), .ZN(W13036));
  INVX1 G46931 (.I(W1551), .ZN(W13037));
  INVX1 G46932 (.I(W1733), .ZN(W13045));
  INVX1 G46933 (.I(W32640), .ZN(O9191));
  INVX1 G46934 (.I(W8420), .ZN(W13051));
  INVX1 G46935 (.I(W2722), .ZN(W13119));
  INVX1 G46936 (.I(W1428), .ZN(W13113));
  INVX1 G46937 (.I(I1535), .ZN(W37722));
  INVX1 G46938 (.I(W32716), .ZN(W37721));
  INVX1 G46939 (.I(W17942), .ZN(O9146));
  INVX1 G46940 (.I(W36299), .ZN(O9145));
  INVX1 G46941 (.I(I1638), .ZN(W13115));
  INVX1 G46942 (.I(W3647), .ZN(O9144));
  INVX1 G46943 (.I(W8697), .ZN(O9143));
  INVX1 G46944 (.I(W6207), .ZN(O697));
  INVX1 G46945 (.I(W9687), .ZN(O9148));
  INVX1 G46946 (.I(W1924), .ZN(O700));
  INVX1 G46947 (.I(W5077), .ZN(W13121));
  INVX1 G46948 (.I(W629), .ZN(W13122));
  INVX1 G46949 (.I(W30814), .ZN(O9139));
  INVX1 G46950 (.I(W34005), .ZN(O9138));
  INVX1 G46951 (.I(W15341), .ZN(W37704));
  INVX1 G46952 (.I(W12314), .ZN(W13126));
  INVX1 G46953 (.I(W25553), .ZN(W37700));
  INVX1 G46954 (.I(W1014), .ZN(W13130));
  INVX1 G46955 (.I(W2668), .ZN(O9157));
  INVX1 G46956 (.I(W4301), .ZN(W13084));
  INVX1 G46957 (.I(W23196), .ZN(O9165));
  INVX1 G46958 (.I(W7154), .ZN(W13087));
  INVX1 G46959 (.I(W26318), .ZN(O9163));
  INVX1 G46960 (.I(W29439), .ZN(O9162));
  INVX1 G46961 (.I(W8524), .ZN(O9161));
  INVX1 G46962 (.I(W1633), .ZN(W13089));
  INVX1 G46963 (.I(W3609), .ZN(W13093));
  INVX1 G46964 (.I(I877), .ZN(W13094));
  INVX1 G46965 (.I(W4766), .ZN(W13275));
  INVX1 G46966 (.I(W16060), .ZN(W37739));
  INVX1 G46967 (.I(W8528), .ZN(W13097));
  INVX1 G46968 (.I(W37191), .ZN(W37735));
  INVX1 G46969 (.I(W4929), .ZN(W13103));
  INVX1 G46970 (.I(W5764), .ZN(O695));
  INVX1 G46971 (.I(W1999), .ZN(W13106));
  INVX1 G46972 (.I(W10597), .ZN(W13109));
  INVX1 G46973 (.I(W8930), .ZN(W13110));
  INVX1 G46974 (.I(W12743), .ZN(O696));
  INVX1 G46975 (.I(W5098), .ZN(O743));
  INVX1 G46976 (.I(W20066), .ZN(W37411));
  INVX1 G46977 (.I(W3409), .ZN(O8966));
  INVX1 G46978 (.I(W8116), .ZN(W37409));
  INVX1 G46979 (.I(W9826), .ZN(W37408));
  INVX1 G46980 (.I(W24908), .ZN(O8964));
  INVX1 G46981 (.I(W19855), .ZN(W37403));
  INVX1 G46982 (.I(W4892), .ZN(W13441));
  INVX1 G46983 (.I(I737), .ZN(O8959));
  INVX1 G46984 (.I(W17259), .ZN(W37395));
  INVX1 G46985 (.I(W23412), .ZN(W37393));
  INVX1 G46986 (.I(I90), .ZN(W13431));
  INVX1 G46987 (.I(I1259), .ZN(W13454));
  INVX1 G46988 (.I(W6632), .ZN(W13455));
  INVX1 G46989 (.I(W34035), .ZN(O8954));
  INVX1 G46990 (.I(W11937), .ZN(W13458));
  INVX1 G46991 (.I(W7041), .ZN(W13460));
  INVX1 G46992 (.I(I1347), .ZN(O745));
  INVX1 G46993 (.I(W33959), .ZN(W37380));
  INVX1 G46994 (.I(W2950), .ZN(O8949));
  INVX1 G46995 (.I(W1070), .ZN(W13464));
  INVX1 G46996 (.I(W2362), .ZN(O8978));
  INVX1 G46997 (.I(W5197), .ZN(W13395));
  INVX1 G46998 (.I(W7703), .ZN(W13399));
  INVX1 G46999 (.I(W12528), .ZN(O738));
  INVX1 G47000 (.I(W5940), .ZN(W13403));
  INVX1 G47001 (.I(W14007), .ZN(W37439));
  INVX1 G47002 (.I(W6635), .ZN(O8981));
  INVX1 G47003 (.I(I1011), .ZN(W13405));
  INVX1 G47004 (.I(W29865), .ZN(O8979));
  INVX1 G47005 (.I(I1472), .ZN(W37434));
  INVX1 G47006 (.I(W17181), .ZN(W37376));
  INVX1 G47007 (.I(W9942), .ZN(W37431));
  INVX1 G47008 (.I(W23191), .ZN(W37430));
  INVX1 G47009 (.I(W4899), .ZN(W13421));
  INVX1 G47010 (.I(W5588), .ZN(W13422));
  INVX1 G47011 (.I(W34650), .ZN(W37421));
  INVX1 G47012 (.I(W7298), .ZN(W13428));
  INVX1 G47013 (.I(W34730), .ZN(O8969));
  INVX1 G47014 (.I(W36084), .ZN(O8968));
  INVX1 G47015 (.I(W17427), .ZN(W37413));
  INVX1 G47016 (.I(W66), .ZN(W37333));
  INVX1 G47017 (.I(W5270), .ZN(W13492));
  INVX1 G47018 (.I(W14189), .ZN(O8925));
  INVX1 G47019 (.I(W8144), .ZN(W13497));
  INVX1 G47020 (.I(W15014), .ZN(O8924));
  INVX1 G47021 (.I(I406), .ZN(W13498));
  INVX1 G47022 (.I(W2529), .ZN(O749));
  INVX1 G47023 (.I(W6969), .ZN(O8921));
  INVX1 G47024 (.I(W5738), .ZN(O750));
  INVX1 G47025 (.I(W9321), .ZN(W13503));
  INVX1 G47026 (.I(W1772), .ZN(O8928));
  INVX1 G47027 (.I(W7018), .ZN(W37332));
  INVX1 G47028 (.I(I290), .ZN(W37331));
  INVX1 G47029 (.I(W14878), .ZN(W37330));
  INVX1 G47030 (.I(I342), .ZN(W37329));
  INVX1 G47031 (.I(W37109), .ZN(O8918));
  INVX1 G47032 (.I(W26175), .ZN(O8915));
  INVX1 G47033 (.I(W12756), .ZN(W13506));
  INVX1 G47034 (.I(W6148), .ZN(W13509));
  INVX1 G47035 (.I(W3361), .ZN(W13513));
  INVX1 G47036 (.I(W15358), .ZN(W37359));
  INVX1 G47037 (.I(W8650), .ZN(W13466));
  INVX1 G47038 (.I(W35312), .ZN(W37374));
  INVX1 G47039 (.I(W392), .ZN(O746));
  INVX1 G47040 (.I(W12658), .ZN(W13471));
  INVX1 G47041 (.I(W3078), .ZN(W13477));
  INVX1 G47042 (.I(W34861), .ZN(O8940));
  INVX1 G47043 (.I(W11710), .ZN(W13479));
  INVX1 G47044 (.I(W17304), .ZN(O8939));
  INVX1 G47045 (.I(W17985), .ZN(O8938));
  INVX1 G47046 (.I(W24437), .ZN(W37447));
  INVX1 G47047 (.I(I1030), .ZN(O8937));
  INVX1 G47048 (.I(W13791), .ZN(O8936));
  INVX1 G47049 (.I(W9558), .ZN(O748));
  INVX1 G47050 (.I(W32654), .ZN(W37355));
  INVX1 G47051 (.I(I1696), .ZN(W13482));
  INVX1 G47052 (.I(W11722), .ZN(W13483));
  INVX1 G47053 (.I(W12368), .ZN(W13485));
  INVX1 G47054 (.I(W12481), .ZN(W37350));
  INVX1 G47055 (.I(W9135), .ZN(O8930));
  INVX1 G47056 (.I(W5364), .ZN(W37519));
  INVX1 G47057 (.I(W27390), .ZN(W37533));
  INVX1 G47058 (.I(W9766), .ZN(W13313));
  INVX1 G47059 (.I(W19073), .ZN(O9033));
  INVX1 G47060 (.I(W11120), .ZN(W13317));
  INVX1 G47061 (.I(W32575), .ZN(O9030));
  INVX1 G47062 (.I(W8461), .ZN(W13324));
  INVX1 G47063 (.I(W6775), .ZN(W37522));
  INVX1 G47064 (.I(W1452), .ZN(O9027));
  INVX1 G47065 (.I(W8367), .ZN(O9026));
  INVX1 G47066 (.I(W16932), .ZN(O9037));
  INVX1 G47067 (.I(I103), .ZN(O728));
  INVX1 G47068 (.I(W19999), .ZN(W37516));
  INVX1 G47069 (.I(W3991), .ZN(W13328));
  INVX1 G47070 (.I(W23041), .ZN(O9024));
  INVX1 G47071 (.I(W3655), .ZN(O731));
  INVX1 G47072 (.I(W6626), .ZN(W13337));
  INVX1 G47073 (.I(W22724), .ZN(W37507));
  INVX1 G47074 (.I(W6985), .ZN(W13338));
  INVX1 G47075 (.I(W30630), .ZN(O9020));
  INVX1 G47076 (.I(W12352), .ZN(O9044));
  INVX1 G47077 (.I(W8202), .ZN(W13276));
  INVX1 G47078 (.I(W25247), .ZN(O9054));
  INVX1 G47079 (.I(W16743), .ZN(O9053));
  INVX1 G47080 (.I(W3362), .ZN(W13279));
  INVX1 G47081 (.I(W6280), .ZN(W13284));
  INVX1 G47082 (.I(W1523), .ZN(W13295));
  INVX1 G47083 (.I(W2907), .ZN(W13296));
  INVX1 G47084 (.I(W7251), .ZN(W13297));
  INVX1 G47085 (.I(W9108), .ZN(O9045));
  INVX1 G47086 (.I(W23032), .ZN(W37504));
  INVX1 G47087 (.I(W6997), .ZN(O9043));
  INVX1 G47088 (.I(W10564), .ZN(W13298));
  INVX1 G47089 (.I(W35658), .ZN(W37546));
  INVX1 G47090 (.I(W1518), .ZN(W13301));
  INVX1 G47091 (.I(I622), .ZN(W13302));
  INVX1 G47092 (.I(I917), .ZN(W13309));
  INVX1 G47093 (.I(W33213), .ZN(O9040));
  INVX1 G47094 (.I(W14793), .ZN(W37538));
  INVX1 G47095 (.I(W13574), .ZN(O9039));
  INVX1 G47096 (.I(W1006), .ZN(W13382));
  INVX1 G47097 (.I(W1661), .ZN(W37476));
  INVX1 G47098 (.I(W20294), .ZN(W37475));
  INVX1 G47099 (.I(I861), .ZN(W13362));
  INVX1 G47100 (.I(W3034), .ZN(W13367));
  INVX1 G47101 (.I(W1738), .ZN(W13371));
  INVX1 G47102 (.I(W20574), .ZN(O8995));
  INVX1 G47103 (.I(W4666), .ZN(W13375));
  INVX1 G47104 (.I(W6342), .ZN(W13379));
  INVX1 G47105 (.I(W35925), .ZN(O8994));
  INVX1 G47106 (.I(W30718), .ZN(O9003));
  INVX1 G47107 (.I(W2332), .ZN(W37460));
  INVX1 G47108 (.I(W5755), .ZN(W13383));
  INVX1 G47109 (.I(W28211), .ZN(O8991));
  INVX1 G47110 (.I(W4039), .ZN(W13384));
  INVX1 G47111 (.I(W3806), .ZN(W13387));
  INVX1 G47112 (.I(I1343), .ZN(W13390));
  INVX1 G47113 (.I(W15547), .ZN(O8989));
  INVX1 G47114 (.I(W17804), .ZN(O8988));
  INVX1 G47115 (.I(W2260), .ZN(W13392));
  INVX1 G47116 (.I(W6459), .ZN(O9010));
  INVX1 G47117 (.I(W3970), .ZN(W13339));
  INVX1 G47118 (.I(W9897), .ZN(W13340));
  INVX1 G47119 (.I(W10910), .ZN(W37500));
  INVX1 G47120 (.I(W997), .ZN(W13345));
  INVX1 G47121 (.I(W4384), .ZN(W13346));
  INVX1 G47122 (.I(W21443), .ZN(O9014));
  INVX1 G47123 (.I(W25579), .ZN(O9012));
  INVX1 G47124 (.I(W31536), .ZN(W37493));
  INVX1 G47125 (.I(W3327), .ZN(W13349));
  INVX1 G47126 (.I(W27331), .ZN(O9785));
  INVX1 G47127 (.I(I990), .ZN(W13350));
  INVX1 G47128 (.I(W8898), .ZN(W37489));
  INVX1 G47129 (.I(W1397), .ZN(W37488));
  INVX1 G47130 (.I(W11731), .ZN(W37487));
  INVX1 G47131 (.I(W321), .ZN(O733));
  INVX1 G47132 (.I(W26783), .ZN(O9007));
  INVX1 G47133 (.I(W11259), .ZN(O734));
  INVX1 G47134 (.I(W11038), .ZN(W13355));
  INVX1 G47135 (.I(W293), .ZN(O9004));
  INVX1 G47136 (.I(W4091), .ZN(W10829));
  INVX1 G47137 (.I(W6328), .ZN(W10821));
  INVX1 G47138 (.I(I887), .ZN(W10823));
  INVX1 G47139 (.I(W3770), .ZN(W10825));
  INVX1 G47140 (.I(W1844), .ZN(W10826));
  INVX1 G47141 (.I(W1315), .ZN(W10827));
  INVX1 G47142 (.I(W10321), .ZN(O10632));
  INVX1 G47143 (.I(W973), .ZN(W10828));
  INVX1 G47144 (.I(W16127), .ZN(O10630));
  INVX1 G47145 (.I(W3091), .ZN(O10629));
  INVX1 G47146 (.I(W5388), .ZN(O10628));
  INVX1 G47147 (.I(W30305), .ZN(O10634));
  INVX1 G47148 (.I(W3784), .ZN(W10830));
  INVX1 G47149 (.I(W7052), .ZN(O10626));
  INVX1 G47150 (.I(W2151), .ZN(O10625));
  INVX1 G47151 (.I(W10465), .ZN(W10837));
  INVX1 G47152 (.I(W264), .ZN(O440));
  INVX1 G47153 (.I(W18927), .ZN(W40031));
  INVX1 G47154 (.I(I1407), .ZN(W10844));
  INVX1 G47155 (.I(W835), .ZN(W10845));
  INVX1 G47156 (.I(W8027), .ZN(W10846));
  INVX1 G47157 (.I(W20843), .ZN(O10644));
  INVX1 G47158 (.I(W5693), .ZN(W40082));
  INVX1 G47159 (.I(W4965), .ZN(W10789));
  INVX1 G47160 (.I(W1986), .ZN(W10793));
  INVX1 G47161 (.I(W6019), .ZN(W10798));
  INVX1 G47162 (.I(W4749), .ZN(W10799));
  INVX1 G47163 (.I(W4948), .ZN(W10800));
  INVX1 G47164 (.I(W4313), .ZN(W40068));
  INVX1 G47165 (.I(I1665), .ZN(W40065));
  INVX1 G47166 (.I(W10493), .ZN(W10805));
  INVX1 G47167 (.I(W34692), .ZN(W40024));
  INVX1 G47168 (.I(W19274), .ZN(O10642));
  INVX1 G47169 (.I(I1844), .ZN(W10807));
  INVX1 G47170 (.I(W4448), .ZN(O438));
  INVX1 G47171 (.I(I748), .ZN(W10809));
  INVX1 G47172 (.I(I1030), .ZN(W10810));
  INVX1 G47173 (.I(W2557), .ZN(W10812));
  INVX1 G47174 (.I(W8637), .ZN(W10813));
  INVX1 G47175 (.I(W28616), .ZN(W40054));
  INVX1 G47176 (.I(I1134), .ZN(W10815));
  INVX1 G47177 (.I(W14628), .ZN(O10585));
  INVX1 G47178 (.I(W765), .ZN(W10874));
  INVX1 G47179 (.I(W5912), .ZN(W10881));
  INVX1 G47180 (.I(I1463), .ZN(W39987));
  INVX1 G47181 (.I(W3212), .ZN(O447));
  INVX1 G47182 (.I(I188), .ZN(W10883));
  INVX1 G47183 (.I(W17431), .ZN(O10590));
  INVX1 G47184 (.I(W17375), .ZN(W39983));
  INVX1 G47185 (.I(W24447), .ZN(O10588));
  INVX1 G47186 (.I(W5103), .ZN(W10888));
  INVX1 G47187 (.I(W6099), .ZN(O10596));
  INVX1 G47188 (.I(W4238), .ZN(O450));
  INVX1 G47189 (.I(W1614), .ZN(W10891));
  INVX1 G47190 (.I(W1733), .ZN(W10893));
  INVX1 G47191 (.I(W646), .ZN(O10581));
  INVX1 G47192 (.I(W2949), .ZN(O451));
  INVX1 G47193 (.I(W24767), .ZN(O10580));
  INVX1 G47194 (.I(W37475), .ZN(O10577));
  INVX1 G47195 (.I(I1391), .ZN(O10574));
  INVX1 G47196 (.I(I163), .ZN(W10912));
  INVX1 G47197 (.I(W3700), .ZN(O10608));
  INVX1 G47198 (.I(W21319), .ZN(W40023));
  INVX1 G47199 (.I(I718), .ZN(W10848));
  INVX1 G47200 (.I(W11329), .ZN(O10617));
  INVX1 G47201 (.I(W11), .ZN(O10616));
  INVX1 G47202 (.I(W2691), .ZN(O10615));
  INVX1 G47203 (.I(W9154), .ZN(W10852));
  INVX1 G47204 (.I(W4724), .ZN(W10854));
  INVX1 G47205 (.I(W6656), .ZN(W10855));
  INVX1 G47206 (.I(W9711), .ZN(O443));
  INVX1 G47207 (.I(W28433), .ZN(O10654));
  INVX1 G47208 (.I(W9745), .ZN(W10858));
  INVX1 G47209 (.I(W3591), .ZN(W10860));
  INVX1 G47210 (.I(W23031), .ZN(O10605));
  INVX1 G47211 (.I(W34302), .ZN(O10603));
  INVX1 G47212 (.I(W22156), .ZN(W40001));
  INVX1 G47213 (.I(W10864), .ZN(W10866));
  INVX1 G47214 (.I(W461), .ZN(W10867));
  INVX1 G47215 (.I(W2519), .ZN(W10869));
  INVX1 G47216 (.I(W1026), .ZN(O444));
  INVX1 G47217 (.I(W37003), .ZN(O10717));
  INVX1 G47218 (.I(W18745), .ZN(O10724));
  INVX1 G47219 (.I(W5362), .ZN(W40178));
  INVX1 G47220 (.I(W13369), .ZN(W40176));
  INVX1 G47221 (.I(W13220), .ZN(W40175));
  INVX1 G47222 (.I(W3290), .ZN(W10693));
  INVX1 G47223 (.I(W9370), .ZN(W10698));
  INVX1 G47224 (.I(W35132), .ZN(O10720));
  INVX1 G47225 (.I(W22006), .ZN(W40169));
  INVX1 G47226 (.I(W31644), .ZN(O10719));
  INVX1 G47227 (.I(W3382), .ZN(O10718));
  INVX1 G47228 (.I(W29220), .ZN(O10725));
  INVX1 G47229 (.I(W5121), .ZN(O425));
  INVX1 G47230 (.I(W22471), .ZN(O10715));
  INVX1 G47231 (.I(W3054), .ZN(W10703));
  INVX1 G47232 (.I(W28541), .ZN(O10713));
  INVX1 G47233 (.I(W9293), .ZN(O10712));
  INVX1 G47234 (.I(W6559), .ZN(W10706));
  INVX1 G47235 (.I(W9831), .ZN(W10712));
  INVX1 G47236 (.I(W6529), .ZN(W10714));
  INVX1 G47237 (.I(W7485), .ZN(W10715));
  INVX1 G47238 (.I(W38714), .ZN(W40202));
  INVX1 G47239 (.I(W8677), .ZN(O10750));
  INVX1 G47240 (.I(W4439), .ZN(O10748));
  INVX1 G47241 (.I(W4262), .ZN(W10655));
  INVX1 G47242 (.I(W3076), .ZN(O417));
  INVX1 G47243 (.I(W29639), .ZN(O10746));
  INVX1 G47244 (.I(W3190), .ZN(W10662));
  INVX1 G47245 (.I(W26929), .ZN(O10742));
  INVX1 G47246 (.I(W30654), .ZN(O10740));
  INVX1 G47247 (.I(W7561), .ZN(W10669));
  INVX1 G47248 (.I(W14945), .ZN(W40147));
  INVX1 G47249 (.I(I463), .ZN(W10671));
  INVX1 G47250 (.I(W13954), .ZN(O10736));
  INVX1 G47251 (.I(I1858), .ZN(O420));
  INVX1 G47252 (.I(W9678), .ZN(W10677));
  INVX1 G47253 (.I(I511), .ZN(O421));
  INVX1 G47254 (.I(W21319), .ZN(O10727));
  INVX1 G47255 (.I(W30973), .ZN(W40185));
  INVX1 G47256 (.I(W3690), .ZN(W40184));
  INVX1 G47257 (.I(W37856), .ZN(O10726));
  INVX1 G47258 (.I(W1192), .ZN(W10766));
  INVX1 G47259 (.I(W2054), .ZN(O10681));
  INVX1 G47260 (.I(W10451), .ZN(W10750));
  INVX1 G47261 (.I(W10917), .ZN(W40114));
  INVX1 G47262 (.I(W4625), .ZN(O10677));
  INVX1 G47263 (.I(W31998), .ZN(W40111));
  INVX1 G47264 (.I(W26609), .ZN(O10676));
  INVX1 G47265 (.I(W33890), .ZN(O10675));
  INVX1 G47266 (.I(W3050), .ZN(W10756));
  INVX1 G47267 (.I(W4498), .ZN(O10669));
  INVX1 G47268 (.I(W19826), .ZN(O10684));
  INVX1 G47269 (.I(W28260), .ZN(O10668));
  INVX1 G47270 (.I(I866), .ZN(W10770));
  INVX1 G47271 (.I(W35139), .ZN(O10665));
  INVX1 G47272 (.I(W21417), .ZN(O10664));
  INVX1 G47273 (.I(W4086), .ZN(W10774));
  INVX1 G47274 (.I(W9294), .ZN(W10775));
  INVX1 G47275 (.I(I615), .ZN(W10776));
  INVX1 G47276 (.I(W23804), .ZN(W40086));
  INVX1 G47277 (.I(W5079), .ZN(W10780));
  INVX1 G47278 (.I(W9400), .ZN(W10732));
  INVX1 G47279 (.I(W28076), .ZN(O10703));
  INVX1 G47280 (.I(W35862), .ZN(O10702));
  INVX1 G47281 (.I(I745), .ZN(W10727));
  INVX1 G47282 (.I(I505), .ZN(W10728));
  INVX1 G47283 (.I(W35962), .ZN(O10700));
  INVX1 G47284 (.I(W1181), .ZN(O10698));
  INVX1 G47285 (.I(I135), .ZN(O427));
  INVX1 G47286 (.I(W9837), .ZN(W40137));
  INVX1 G47287 (.I(W38980), .ZN(O10696));
  INVX1 G47288 (.I(W2737), .ZN(W39955));
  INVX1 G47289 (.I(W7153), .ZN(W10734));
  INVX1 G47290 (.I(W24069), .ZN(O10694));
  INVX1 G47291 (.I(W562), .ZN(W10737));
  INVX1 G47292 (.I(W5223), .ZN(W10741));
  INVX1 G47293 (.I(W37440), .ZN(O10691));
  INVX1 G47294 (.I(W30275), .ZN(W40128));
  INVX1 G47295 (.I(W18802), .ZN(O10690));
  INVX1 G47296 (.I(W36877), .ZN(O10689));
  INVX1 G47297 (.I(W4533), .ZN(O10687));
  INVX1 G47298 (.I(W1203), .ZN(W11071));
  INVX1 G47299 (.I(W394), .ZN(W39810));
  INVX1 G47300 (.I(I752), .ZN(O475));
  INVX1 G47301 (.I(W8705), .ZN(O476));
  INVX1 G47302 (.I(W2407), .ZN(W11060));
  INVX1 G47303 (.I(W38669), .ZN(O10460));
  INVX1 G47304 (.I(I1892), .ZN(O10458));
  INVX1 G47305 (.I(W9039), .ZN(W11065));
  INVX1 G47306 (.I(W6839), .ZN(W11066));
  INVX1 G47307 (.I(W16988), .ZN(W39799));
  INVX1 G47308 (.I(I192), .ZN(W11067));
  INVX1 G47309 (.I(W9544), .ZN(O10465));
  INVX1 G47310 (.I(W24435), .ZN(O10454));
  INVX1 G47311 (.I(W34583), .ZN(O10453));
  INVX1 G47312 (.I(W8257), .ZN(W11075));
  INVX1 G47313 (.I(I1339), .ZN(W11078));
  INVX1 G47314 (.I(W10173), .ZN(O477));
  INVX1 G47315 (.I(W492), .ZN(W11084));
  INVX1 G47316 (.I(W1880), .ZN(W39788));
  INVX1 G47317 (.I(W5214), .ZN(O10448));
  INVX1 G47318 (.I(W32364), .ZN(W39786));
  INVX1 G47319 (.I(W6750), .ZN(W11030));
  INVX1 G47320 (.I(W7932), .ZN(W11016));
  INVX1 G47321 (.I(W8425), .ZN(W11020));
  INVX1 G47322 (.I(W14791), .ZN(O10488));
  INVX1 G47323 (.I(I1726), .ZN(O10487));
  INVX1 G47324 (.I(W4899), .ZN(O468));
  INVX1 G47325 (.I(W8494), .ZN(W11025));
  INVX1 G47326 (.I(W12169), .ZN(O10482));
  INVX1 G47327 (.I(W3081), .ZN(W39831));
  INVX1 G47328 (.I(I647), .ZN(W11027));
  INVX1 G47329 (.I(W887), .ZN(O480));
  INVX1 G47330 (.I(W7141), .ZN(O471));
  INVX1 G47331 (.I(W910), .ZN(W11037));
  INVX1 G47332 (.I(W9883), .ZN(O473));
  INVX1 G47333 (.I(W9247), .ZN(W39819));
  INVX1 G47334 (.I(W21731), .ZN(O10470));
  INVX1 G47335 (.I(I987), .ZN(W11042));
  INVX1 G47336 (.I(W6812), .ZN(W11046));
  INVX1 G47337 (.I(W2499), .ZN(W11047));
  INVX1 G47338 (.I(W9612), .ZN(W11049));
  INVX1 G47339 (.I(W32440), .ZN(O10423));
  INVX1 G47340 (.I(W29265), .ZN(O10430));
  INVX1 G47341 (.I(W5734), .ZN(W11117));
  INVX1 G47342 (.I(W10651), .ZN(O10428));
  INVX1 G47343 (.I(W11679), .ZN(W39752));
  INVX1 G47344 (.I(W32071), .ZN(O10427));
  INVX1 G47345 (.I(W14220), .ZN(O10426));
  INVX1 G47346 (.I(W32913), .ZN(O10425));
  INVX1 G47347 (.I(W21263), .ZN(W39748));
  INVX1 G47348 (.I(W1157), .ZN(W11120));
  INVX1 G47349 (.I(W3417), .ZN(W11116));
  INVX1 G47350 (.I(W34946), .ZN(W39745));
  INVX1 G47351 (.I(W9939), .ZN(W11121));
  INVX1 G47352 (.I(W4358), .ZN(W11122));
  INVX1 G47353 (.I(W7883), .ZN(W11124));
  INVX1 G47354 (.I(W6162), .ZN(O483));
  INVX1 G47355 (.I(W5160), .ZN(W11126));
  INVX1 G47356 (.I(W6875), .ZN(W11127));
  INVX1 G47357 (.I(W12161), .ZN(O10416));
  INVX1 G47358 (.I(W16937), .ZN(O10415));
  INVX1 G47359 (.I(I1026), .ZN(W11110));
  INVX1 G47360 (.I(I1575), .ZN(O10444));
  INVX1 G47361 (.I(W1279), .ZN(W11092));
  INVX1 G47362 (.I(W9519), .ZN(W11093));
  INVX1 G47363 (.I(W6636), .ZN(W11094));
  INVX1 G47364 (.I(W1820), .ZN(W11095));
  INVX1 G47365 (.I(W3071), .ZN(W11098));
  INVX1 G47366 (.I(W3268), .ZN(W11104));
  INVX1 G47367 (.I(W7530), .ZN(W11107));
  INVX1 G47368 (.I(W2593), .ZN(W11108));
  INVX1 G47369 (.I(W34540), .ZN(O10493));
  INVX1 G47370 (.I(W18596), .ZN(W39767));
  INVX1 G47371 (.I(W38455), .ZN(W39766));
  INVX1 G47372 (.I(W21833), .ZN(W39765));
  INVX1 G47373 (.I(W6409), .ZN(W11113));
  INVX1 G47374 (.I(W31721), .ZN(O10435));
  INVX1 G47375 (.I(W7770), .ZN(W11115));
  INVX1 G47376 (.I(W2534), .ZN(O10433));
  INVX1 G47377 (.I(W5488), .ZN(O10432));
  INVX1 G47378 (.I(W18309), .ZN(W39757));
  INVX1 G47379 (.I(W21964), .ZN(O10545));
  INVX1 G47380 (.I(W24179), .ZN(O10556));
  INVX1 G47381 (.I(W38744), .ZN(O10555));
  INVX1 G47382 (.I(W31482), .ZN(O10554));
  INVX1 G47383 (.I(W24941), .ZN(O10551));
  INVX1 G47384 (.I(I1960), .ZN(W10936));
  INVX1 G47385 (.I(W17721), .ZN(O10548));
  INVX1 G47386 (.I(W30420), .ZN(W39918));
  INVX1 G47387 (.I(W979), .ZN(W10941));
  INVX1 G47388 (.I(W875), .ZN(W10943));
  INVX1 G47389 (.I(W2432), .ZN(W10927));
  INVX1 G47390 (.I(W38505), .ZN(W39914));
  INVX1 G47391 (.I(W31379), .ZN(O10544));
  INVX1 G47392 (.I(W15856), .ZN(O10543));
  INVX1 G47393 (.I(W35620), .ZN(W39909));
  INVX1 G47394 (.I(W4378), .ZN(W10948));
  INVX1 G47395 (.I(W36680), .ZN(W39906));
  INVX1 G47396 (.I(W7100), .ZN(W10949));
  INVX1 G47397 (.I(I1016), .ZN(W10953));
  INVX1 G47398 (.I(W1380), .ZN(W10954));
  INVX1 G47399 (.I(W3903), .ZN(W10918));
  INVX1 G47400 (.I(W9323), .ZN(W10913));
  INVX1 G47401 (.I(W14879), .ZN(O10570));
  INVX1 G47402 (.I(W4559), .ZN(W10914));
  INVX1 G47403 (.I(W36104), .ZN(O10569));
  INVX1 G47404 (.I(W9922), .ZN(O10568));
  INVX1 G47405 (.I(W1202), .ZN(O453));
  INVX1 G47406 (.I(W12773), .ZN(W39948));
  INVX1 G47407 (.I(W34049), .ZN(O10566));
  INVX1 G47408 (.I(W18148), .ZN(W39946));
  INVX1 G47409 (.I(W8083), .ZN(W10959));
  INVX1 G47410 (.I(W19838), .ZN(W39942));
  INVX1 G47411 (.I(W8337), .ZN(W10921));
  INVX1 G47412 (.I(W25679), .ZN(O10561));
  INVX1 G47413 (.I(W20220), .ZN(O10560));
  INVX1 G47414 (.I(W544), .ZN(W10925));
  INVX1 G47415 (.I(W22509), .ZN(O10559));
  INVX1 G47416 (.I(W23627), .ZN(W39934));
  INVX1 G47417 (.I(W9176), .ZN(W39933));
  INVX1 G47418 (.I(W1532), .ZN(W10926));
  INVX1 G47419 (.I(W2628), .ZN(W11007));
  INVX1 G47420 (.I(W4950), .ZN(W11001));
  INVX1 G47421 (.I(W34040), .ZN(O10510));
  INVX1 G47422 (.I(W3217), .ZN(W11003));
  INVX1 G47423 (.I(W33373), .ZN(O10508));
  INVX1 G47424 (.I(W36870), .ZN(O10507));
  INVX1 G47425 (.I(W2521), .ZN(O10506));
  INVX1 G47426 (.I(W10783), .ZN(O10505));
  INVX1 G47427 (.I(W9069), .ZN(O462));
  INVX1 G47428 (.I(W39314), .ZN(W39858));
  INVX1 G47429 (.I(W5180), .ZN(W11000));
  INVX1 G47430 (.I(W25708), .ZN(O10502));
  INVX1 G47431 (.I(I596), .ZN(O10501));
  INVX1 G47432 (.I(W33141), .ZN(W39854));
  INVX1 G47433 (.I(I1620), .ZN(O10498));
  INVX1 G47434 (.I(W6681), .ZN(O465));
  INVX1 G47435 (.I(W10690), .ZN(W39848));
  INVX1 G47436 (.I(W10141), .ZN(O10496));
  INVX1 G47437 (.I(W38982), .ZN(O10495));
  INVX1 G47438 (.I(W4446), .ZN(W11013));
  INVX1 G47439 (.I(W25138), .ZN(O10523));
  INVX1 G47440 (.I(W23775), .ZN(W39897));
  INVX1 G47441 (.I(W6454), .ZN(W10961));
  INVX1 G47442 (.I(W2518), .ZN(W10969));
  INVX1 G47443 (.I(W5085), .ZN(W10970));
  INVX1 G47444 (.I(W2759), .ZN(O458));
  INVX1 G47445 (.I(W32205), .ZN(W39890));
  INVX1 G47446 (.I(W8559), .ZN(W10974));
  INVX1 G47447 (.I(W10137), .ZN(O10525));
  INVX1 G47448 (.I(W5208), .ZN(W10977));
  INVX1 G47449 (.I(I549), .ZN(W10646));
  INVX1 G47450 (.I(I1482), .ZN(W10980));
  INVX1 G47451 (.I(W9159), .ZN(W10983));
  INVX1 G47452 (.I(W33424), .ZN(W39879));
  INVX1 G47453 (.I(W634), .ZN(W10990));
  INVX1 G47454 (.I(W338), .ZN(O461));
  INVX1 G47455 (.I(W13136), .ZN(O10517));
  INVX1 G47456 (.I(W9800), .ZN(O10516));
  INVX1 G47457 (.I(I1739), .ZN(W10994));
  INVX1 G47458 (.I(W5498), .ZN(W39870));
  INVX1 G47459 (.I(I1697), .ZN(W10351));
  INVX1 G47460 (.I(W14042), .ZN(O10982));
  INVX1 G47461 (.I(W5448), .ZN(W10329));
  INVX1 G47462 (.I(W28018), .ZN(W40552));
  INVX1 G47463 (.I(W13868), .ZN(W40550));
  INVX1 G47464 (.I(W3012), .ZN(O10979));
  INVX1 G47465 (.I(W5320), .ZN(W10341));
  INVX1 G47466 (.I(W7912), .ZN(W10342));
  INVX1 G47467 (.I(W6331), .ZN(W10345));
  INVX1 G47468 (.I(W40519), .ZN(O10973));
  INVX1 G47469 (.I(W3254), .ZN(W10350));
  INVX1 G47470 (.I(W9423), .ZN(W10327));
  INVX1 G47471 (.I(W10331), .ZN(W40538));
  INVX1 G47472 (.I(W34636), .ZN(W40536));
  INVX1 G47473 (.I(W1306), .ZN(W10356));
  INVX1 G47474 (.I(W1805), .ZN(W10363));
  INVX1 G47475 (.I(W7797), .ZN(W40529));
  INVX1 G47476 (.I(W6980), .ZN(O10964));
  INVX1 G47477 (.I(W6900), .ZN(W10371));
  INVX1 G47478 (.I(W26270), .ZN(W40524));
  INVX1 G47479 (.I(I169), .ZN(W10376));
  INVX1 G47480 (.I(W20970), .ZN(W40566));
  INVX1 G47481 (.I(W9731), .ZN(W10306));
  INVX1 G47482 (.I(W7152), .ZN(W10307));
  INVX1 G47483 (.I(I1698), .ZN(O381));
  INVX1 G47484 (.I(W3443), .ZN(W10310));
  INVX1 G47485 (.I(I370), .ZN(W10311));
  INVX1 G47486 (.I(W25314), .ZN(W40570));
  INVX1 G47487 (.I(W5441), .ZN(O382));
  INVX1 G47488 (.I(W9531), .ZN(W10313));
  INVX1 G47489 (.I(W9183), .ZN(W10314));
  INVX1 G47490 (.I(W35981), .ZN(W40521));
  INVX1 G47491 (.I(W37465), .ZN(O10989));
  INVX1 G47492 (.I(W33775), .ZN(O10988));
  INVX1 G47493 (.I(W6896), .ZN(W10320));
  INVX1 G47494 (.I(W6220), .ZN(W10322));
  INVX1 G47495 (.I(W8045), .ZN(O10985));
  INVX1 G47496 (.I(W16109), .ZN(W40559));
  INVX1 G47497 (.I(W4298), .ZN(W10325));
  INVX1 G47498 (.I(W5450), .ZN(W10326));
  INVX1 G47499 (.I(W28846), .ZN(W40556));
  INVX1 G47500 (.I(W9150), .ZN(W10414));
  INVX1 G47501 (.I(W4463), .ZN(W10398));
  INVX1 G47502 (.I(W29657), .ZN(W40488));
  INVX1 G47503 (.I(W722), .ZN(O10934));
  INVX1 G47504 (.I(W7060), .ZN(W10405));
  INVX1 G47505 (.I(W686), .ZN(W10406));
  INVX1 G47506 (.I(W23725), .ZN(O10931));
  INVX1 G47507 (.I(W3411), .ZN(O388));
  INVX1 G47508 (.I(W8734), .ZN(W10408));
  INVX1 G47509 (.I(W7086), .ZN(W10411));
  INVX1 G47510 (.I(W33157), .ZN(O10936));
  INVX1 G47511 (.I(W15796), .ZN(W40474));
  INVX1 G47512 (.I(W20745), .ZN(O10926));
  INVX1 G47513 (.I(W8157), .ZN(W10418));
  INVX1 G47514 (.I(W8474), .ZN(W10420));
  INVX1 G47515 (.I(I1347), .ZN(W10421));
  INVX1 G47516 (.I(W8448), .ZN(W10425));
  INVX1 G47517 (.I(W30603), .ZN(W40466));
  INVX1 G47518 (.I(W18960), .ZN(O10920));
  INVX1 G47519 (.I(W6893), .ZN(W10426));
  INVX1 G47520 (.I(W36328), .ZN(O10946));
  INVX1 G47521 (.I(W29087), .ZN(O10956));
  INVX1 G47522 (.I(W153), .ZN(O385));
  INVX1 G47523 (.I(W37977), .ZN(W40510));
  INVX1 G47524 (.I(W8183), .ZN(O386));
  INVX1 G47525 (.I(W12628), .ZN(O10951));
  INVX1 G47526 (.I(W10585), .ZN(O10950));
  INVX1 G47527 (.I(W3935), .ZN(O387));
  INVX1 G47528 (.I(W13956), .ZN(O10947));
  INVX1 G47529 (.I(W35972), .ZN(W40502));
  INVX1 G47530 (.I(W9069), .ZN(W10303));
  INVX1 G47531 (.I(W10331), .ZN(W10391));
  INVX1 G47532 (.I(W8570), .ZN(W10392));
  INVX1 G47533 (.I(I1011), .ZN(W10393));
  INVX1 G47534 (.I(W5610), .ZN(O10943));
  INVX1 G47535 (.I(I1811), .ZN(O10942));
  INVX1 G47536 (.I(W372), .ZN(W10394));
  INVX1 G47537 (.I(W1817), .ZN(W10395));
  INVX1 G47538 (.I(I1356), .ZN(W10397));
  INVX1 G47539 (.I(W10949), .ZN(O10937));
  INVX1 G47540 (.I(W10183), .ZN(W10228));
  INVX1 G47541 (.I(W2559), .ZN(O11060));
  INVX1 G47542 (.I(W11600), .ZN(O11059));
  INVX1 G47543 (.I(W30471), .ZN(O11058));
  INVX1 G47544 (.I(W34048), .ZN(O11057));
  INVX1 G47545 (.I(W2777), .ZN(O372));
  INVX1 G47546 (.I(I464), .ZN(W10218));
  INVX1 G47547 (.I(W8994), .ZN(W10219));
  INVX1 G47548 (.I(W2222), .ZN(W10220));
  INVX1 G47549 (.I(W4604), .ZN(W10227));
  INVX1 G47550 (.I(W3265), .ZN(O371));
  INVX1 G47551 (.I(W16834), .ZN(W40649));
  INVX1 G47552 (.I(W10019), .ZN(W10229));
  INVX1 G47553 (.I(W31789), .ZN(W40647));
  INVX1 G47554 (.I(W34331), .ZN(O11049));
  INVX1 G47555 (.I(W8434), .ZN(W10231));
  INVX1 G47556 (.I(I1682), .ZN(W40643));
  INVX1 G47557 (.I(W23590), .ZN(O11047));
  INVX1 G47558 (.I(W3581), .ZN(W10233));
  INVX1 G47559 (.I(W3288), .ZN(W10234));
  INVX1 G47560 (.I(W1200), .ZN(W10201));
  INVX1 G47561 (.I(W22969), .ZN(O11074));
  INVX1 G47562 (.I(W5372), .ZN(W10188));
  INVX1 G47563 (.I(W489), .ZN(O370));
  INVX1 G47564 (.I(W37025), .ZN(O11073));
  INVX1 G47565 (.I(W9409), .ZN(W10193));
  INVX1 G47566 (.I(I1002), .ZN(W10195));
  INVX1 G47567 (.I(W1026), .ZN(W10196));
  INVX1 G47568 (.I(W7911), .ZN(W10198));
  INVX1 G47569 (.I(W19810), .ZN(W40679));
  INVX1 G47570 (.I(W3257), .ZN(W10236));
  INVX1 G47571 (.I(W30297), .ZN(W40674));
  INVX1 G47572 (.I(I1870), .ZN(W10205));
  INVX1 G47573 (.I(W2717), .ZN(W10206));
  INVX1 G47574 (.I(W28298), .ZN(W40670));
  INVX1 G47575 (.I(W3558), .ZN(O11066));
  INVX1 G47576 (.I(W2306), .ZN(W10210));
  INVX1 G47577 (.I(W37658), .ZN(O11064));
  INVX1 G47578 (.I(W7589), .ZN(O11063));
  INVX1 G47579 (.I(W22263), .ZN(W40664));
  INVX1 G47580 (.I(W39831), .ZN(O11007));
  INVX1 G47581 (.I(W1908), .ZN(O375));
  INVX1 G47582 (.I(W28090), .ZN(O11019));
  INVX1 G47583 (.I(W212), .ZN(O11018));
  INVX1 G47584 (.I(W8979), .ZN(W10278));
  INVX1 G47585 (.I(W29721), .ZN(O11015));
  INVX1 G47586 (.I(W32382), .ZN(O11014));
  INVX1 G47587 (.I(W7361), .ZN(W10280));
  INVX1 G47588 (.I(W27421), .ZN(W40594));
  INVX1 G47589 (.I(W3858), .ZN(W10289));
  INVX1 G47590 (.I(W10218), .ZN(W10273));
  INVX1 G47591 (.I(W4058), .ZN(W10291));
  INVX1 G47592 (.I(W7324), .ZN(W10296));
  INVX1 G47593 (.I(W8037), .ZN(O11003));
  INVX1 G47594 (.I(W10454), .ZN(O11002));
  INVX1 G47595 (.I(W7367), .ZN(W10297));
  INVX1 G47596 (.I(W6495), .ZN(W10300));
  INVX1 G47597 (.I(W26776), .ZN(O10999));
  INVX1 G47598 (.I(W11766), .ZN(O10997));
  INVX1 G47599 (.I(W9287), .ZN(W10302));
  INVX1 G47600 (.I(W6485), .ZN(W10255));
  INVX1 G47601 (.I(W9462), .ZN(O11044));
  INVX1 G47602 (.I(W4215), .ZN(W10238));
  INVX1 G47603 (.I(W33419), .ZN(O11042));
  INVX1 G47604 (.I(W9544), .ZN(W10239));
  INVX1 G47605 (.I(W8745), .ZN(W10240));
  INVX1 G47606 (.I(W6053), .ZN(W10248));
  INVX1 G47607 (.I(W10709), .ZN(W40626));
  INVX1 G47608 (.I(W19512), .ZN(W40625));
  INVX1 G47609 (.I(W21561), .ZN(O11032));
  INVX1 G47610 (.I(W3843), .ZN(W10427));
  INVX1 G47611 (.I(I1502), .ZN(W10261));
  INVX1 G47612 (.I(W6615), .ZN(O11028));
  INVX1 G47613 (.I(I1814), .ZN(W10262));
  INVX1 G47614 (.I(W7293), .ZN(W10264));
  INVX1 G47615 (.I(W27501), .ZN(O11026));
  INVX1 G47616 (.I(W1580), .ZN(W10267));
  INVX1 G47617 (.I(W2714), .ZN(W10268));
  INVX1 G47618 (.I(W1858), .ZN(O374));
  INVX1 G47619 (.I(I1053), .ZN(O11022));
  INVX1 G47620 (.I(I494), .ZN(W10572));
  INVX1 G47621 (.I(W830), .ZN(W10566));
  INVX1 G47622 (.I(W16628), .ZN(W40311));
  INVX1 G47623 (.I(W13199), .ZN(W40310));
  INVX1 G47624 (.I(W261), .ZN(O10807));
  INVX1 G47625 (.I(W8276), .ZN(W10568));
  INVX1 G47626 (.I(W39848), .ZN(W40307));
  INVX1 G47627 (.I(W9327), .ZN(O10806));
  INVX1 G47628 (.I(W2716), .ZN(W40305));
  INVX1 G47629 (.I(W439), .ZN(W10569));
  INVX1 G47630 (.I(W28803), .ZN(O10805));
  INVX1 G47631 (.I(W30100), .ZN(W40314));
  INVX1 G47632 (.I(W14308), .ZN(O10803));
  INVX1 G47633 (.I(W31409), .ZN(W40299));
  INVX1 G47634 (.I(W36859), .ZN(O10802));
  INVX1 G47635 (.I(W4655), .ZN(W10575));
  INVX1 G47636 (.I(W20426), .ZN(O10800));
  INVX1 G47637 (.I(W23679), .ZN(O10799));
  INVX1 G47638 (.I(W3070), .ZN(O408));
  INVX1 G47639 (.I(W7418), .ZN(W10579));
  INVX1 G47640 (.I(W3904), .ZN(W10581));
  INVX1 G47641 (.I(W182), .ZN(O10817));
  INVX1 G47642 (.I(W6559), .ZN(W10532));
  INVX1 G47643 (.I(W4418), .ZN(W10534));
  INVX1 G47644 (.I(W23395), .ZN(W40340));
  INVX1 G47645 (.I(W9514), .ZN(W10539));
  INVX1 G47646 (.I(W5025), .ZN(W10541));
  INVX1 G47647 (.I(W6155), .ZN(W10542));
  INVX1 G47648 (.I(W7733), .ZN(W10546));
  INVX1 G47649 (.I(W6918), .ZN(O10819));
  INVX1 G47650 (.I(W10483), .ZN(W40333));
  INVX1 G47651 (.I(W5973), .ZN(O10796));
  INVX1 G47652 (.I(W10201), .ZN(W10548));
  INVX1 G47653 (.I(W19450), .ZN(O10815));
  INVX1 G47654 (.I(W39146), .ZN(O10813));
  INVX1 G47655 (.I(W8818), .ZN(W10557));
  INVX1 G47656 (.I(W34471), .ZN(W40320));
  INVX1 G47657 (.I(W2539), .ZN(W10558));
  INVX1 G47658 (.I(I1000), .ZN(W10559));
  INVX1 G47659 (.I(W14664), .ZN(O10810));
  INVX1 G47660 (.I(W6988), .ZN(O405));
  INVX1 G47661 (.I(W6404), .ZN(O10763));
  INVX1 G47662 (.I(W104), .ZN(W10622));
  INVX1 G47663 (.I(W5217), .ZN(O10771));
  INVX1 G47664 (.I(I530), .ZN(O412));
  INVX1 G47665 (.I(W8372), .ZN(O10767));
  INVX1 G47666 (.I(W28896), .ZN(W40243));
  INVX1 G47667 (.I(W39137), .ZN(W40241));
  INVX1 G47668 (.I(W37937), .ZN(W40240));
  INVX1 G47669 (.I(W8001), .ZN(W10635));
  INVX1 G47670 (.I(W15398), .ZN(O10764));
  INVX1 G47671 (.I(W22977), .ZN(O10773));
  INVX1 G47672 (.I(W3084), .ZN(W10637));
  INVX1 G47673 (.I(W2749), .ZN(O414));
  INVX1 G47674 (.I(W6867), .ZN(W10640));
  INVX1 G47675 (.I(W38646), .ZN(O10759));
  INVX1 G47676 (.I(W13493), .ZN(O10758));
  INVX1 G47677 (.I(W14745), .ZN(O10757));
  INVX1 G47678 (.I(W8157), .ZN(O10756));
  INVX1 G47679 (.I(W38822), .ZN(W40226));
  INVX1 G47680 (.I(W3655), .ZN(W10645));
  INVX1 G47681 (.I(W2457), .ZN(W10595));
  INVX1 G47682 (.I(I1500), .ZN(W10582));
  INVX1 G47683 (.I(W5118), .ZN(W40286));
  INVX1 G47684 (.I(W8173), .ZN(W40284));
  INVX1 G47685 (.I(W24997), .ZN(O10793));
  INVX1 G47686 (.I(W1953), .ZN(W10587));
  INVX1 G47687 (.I(W7311), .ZN(W10589));
  INVX1 G47688 (.I(W34053), .ZN(O10788));
  INVX1 G47689 (.I(W3462), .ZN(W10594));
  INVX1 G47690 (.I(W32794), .ZN(O10786));
  INVX1 G47691 (.I(W9612), .ZN(W10530));
  INVX1 G47692 (.I(W9776), .ZN(W40271));
  INVX1 G47693 (.I(W8864), .ZN(W10597));
  INVX1 G47694 (.I(W32448), .ZN(W40267));
  INVX1 G47695 (.I(I455), .ZN(W10604));
  INVX1 G47696 (.I(W28092), .ZN(W40262));
  INVX1 G47697 (.I(W28498), .ZN(W40260));
  INVX1 G47698 (.I(W5130), .ZN(W10607));
  INVX1 G47699 (.I(I732), .ZN(O409));
  INVX1 G47700 (.I(W11145), .ZN(O10774));
  INVX1 G47701 (.I(W6202), .ZN(W10463));
  INVX1 G47702 (.I(W5154), .ZN(O10898));
  INVX1 G47703 (.I(W6555), .ZN(O391));
  INVX1 G47704 (.I(W31080), .ZN(O10895));
  INVX1 G47705 (.I(W7228), .ZN(W10448));
  INVX1 G47706 (.I(W36270), .ZN(W40431));
  INVX1 G47707 (.I(W8362), .ZN(W10455));
  INVX1 G47708 (.I(W11273), .ZN(O10890));
  INVX1 G47709 (.I(W869), .ZN(O393));
  INVX1 G47710 (.I(W16324), .ZN(O10886));
  INVX1 G47711 (.I(W5651), .ZN(O10899));
  INVX1 G47712 (.I(W20570), .ZN(W40423));
  INVX1 G47713 (.I(W8502), .ZN(W10464));
  INVX1 G47714 (.I(W35242), .ZN(O10883));
  INVX1 G47715 (.I(W10328), .ZN(O395));
  INVX1 G47716 (.I(W36737), .ZN(O10881));
  INVX1 G47717 (.I(W3912), .ZN(W10471));
  INVX1 G47718 (.I(W6270), .ZN(W10472));
  INVX1 G47719 (.I(W9924), .ZN(W10473));
  INVX1 G47720 (.I(W25795), .ZN(O10877));
  INVX1 G47721 (.I(W8813), .ZN(O10909));
  INVX1 G47722 (.I(W2007), .ZN(W10428));
  INVX1 G47723 (.I(W3952), .ZN(W10430));
  INVX1 G47724 (.I(W20268), .ZN(O10916));
  INVX1 G47725 (.I(W3421), .ZN(W10431));
  INVX1 G47726 (.I(W276), .ZN(O389));
  INVX1 G47727 (.I(W16104), .ZN(O10913));
  INVX1 G47728 (.I(W18748), .ZN(O10912));
  INVX1 G47729 (.I(W34372), .ZN(O10911));
  INVX1 G47730 (.I(W15442), .ZN(O10910));
  INVX1 G47731 (.I(W10138), .ZN(O397));
  INVX1 G47732 (.I(W7166), .ZN(W10433));
  INVX1 G47733 (.I(W13890), .ZN(W40450));
  INVX1 G47734 (.I(W28275), .ZN(O10906));
  INVX1 G47735 (.I(W7144), .ZN(W10436));
  INVX1 G47736 (.I(W7952), .ZN(W10438));
  INVX1 G47737 (.I(W22512), .ZN(O10903));
  INVX1 G47738 (.I(W7293), .ZN(W10439));
  INVX1 G47739 (.I(W2248), .ZN(O10900));
  INVX1 G47740 (.I(I1357), .ZN(W40440));
  INVX1 G47741 (.I(W885), .ZN(W10521));
  INVX1 G47742 (.I(W31204), .ZN(W40374));
  INVX1 G47743 (.I(W20503), .ZN(O10846));
  INVX1 G47744 (.I(W6196), .ZN(O402));
  INVX1 G47745 (.I(W32897), .ZN(O10844));
  INVX1 G47746 (.I(W7699), .ZN(O10843));
  INVX1 G47747 (.I(W9522), .ZN(W10517));
  INVX1 G47748 (.I(W1875), .ZN(W40364));
  INVX1 G47749 (.I(I1866), .ZN(W10518));
  INVX1 G47750 (.I(W5402), .ZN(W10519));
  INVX1 G47751 (.I(I1092), .ZN(W10510));
  INVX1 G47752 (.I(I1686), .ZN(W10522));
  INVX1 G47753 (.I(I1566), .ZN(W10523));
  INVX1 G47754 (.I(I1044), .ZN(W10527));
  INVX1 G47755 (.I(W9815), .ZN(W10528));
  INVX1 G47756 (.I(W39637), .ZN(W40354));
  INVX1 G47757 (.I(W14492), .ZN(O10830));
  INVX1 G47758 (.I(W30267), .ZN(O10829));
  INVX1 G47759 (.I(W39790), .ZN(O10828));
  INVX1 G47760 (.I(W15339), .ZN(W40349));
  INVX1 G47761 (.I(W6324), .ZN(W10493));
  INVX1 G47762 (.I(W6253), .ZN(O10870));
  INVX1 G47763 (.I(W4080), .ZN(W40404));
  INVX1 G47764 (.I(W28692), .ZN(O10869));
  INVX1 G47765 (.I(W1788), .ZN(W10484));
  INVX1 G47766 (.I(W33311), .ZN(O10867));
  INVX1 G47767 (.I(W13893), .ZN(O10866));
  INVX1 G47768 (.I(W6604), .ZN(O10863));
  INVX1 G47769 (.I(I619), .ZN(W10492));
  INVX1 G47770 (.I(W678), .ZN(W40392));
  INVX1 G47771 (.I(W32183), .ZN(O10414));
  INVX1 G47772 (.I(W37126), .ZN(O10859));
  INVX1 G47773 (.I(W9442), .ZN(W10495));
  INVX1 G47774 (.I(W24454), .ZN(O10857));
  INVX1 G47775 (.I(W4893), .ZN(O10856));
  INVX1 G47776 (.I(W4679), .ZN(W10496));
  INVX1 G47777 (.I(W19612), .ZN(O10854));
  INVX1 G47778 (.I(W5550), .ZN(O10853));
  INVX1 G47779 (.I(W9051), .ZN(W10501));
  INVX1 G47780 (.I(W2436), .ZN(W10509));
  INVX1 G47781 (.I(W8769), .ZN(W11750));
  INVX1 G47782 (.I(W8714), .ZN(W11737));
  INVX1 G47783 (.I(W18178), .ZN(O9985));
  INVX1 G47784 (.I(W16162), .ZN(O9984));
  INVX1 G47785 (.I(W8289), .ZN(W11739));
  INVX1 G47786 (.I(W10940), .ZN(W11740));
  INVX1 G47787 (.I(W10016), .ZN(O9980));
  INVX1 G47788 (.I(W2592), .ZN(O9979));
  INVX1 G47789 (.I(W3649), .ZN(W11746));
  INVX1 G47790 (.I(W5061), .ZN(W11748));
  INVX1 G47791 (.I(W18685), .ZN(O9975));
  INVX1 G47792 (.I(W29372), .ZN(O9987));
  INVX1 G47793 (.I(W2049), .ZN(W11755));
  INVX1 G47794 (.I(W9621), .ZN(W11756));
  INVX1 G47795 (.I(W31896), .ZN(O9971));
  INVX1 G47796 (.I(W28779), .ZN(O9970));
  INVX1 G47797 (.I(W9272), .ZN(W11760));
  INVX1 G47798 (.I(W4699), .ZN(W39094));
  INVX1 G47799 (.I(W739), .ZN(W39092));
  INVX1 G47800 (.I(W3823), .ZN(W11762));
  INVX1 G47801 (.I(W6340), .ZN(W11763));
  INVX1 G47802 (.I(W7451), .ZN(W11718));
  INVX1 G47803 (.I(W23754), .ZN(O10011));
  INVX1 G47804 (.I(W10834), .ZN(W11703));
  INVX1 G47805 (.I(W6818), .ZN(W11708));
  INVX1 G47806 (.I(W6037), .ZN(O10006));
  INVX1 G47807 (.I(W20094), .ZN(W39144));
  INVX1 G47808 (.I(W3547), .ZN(O10003));
  INVX1 G47809 (.I(W3677), .ZN(W11715));
  INVX1 G47810 (.I(W6422), .ZN(W11717));
  INVX1 G47811 (.I(W9499), .ZN(O10000));
  INVX1 G47812 (.I(W11680), .ZN(W11765));
  INVX1 G47813 (.I(I1636), .ZN(W11721));
  INVX1 G47814 (.I(W10782), .ZN(W11723));
  INVX1 G47815 (.I(I1348), .ZN(W11725));
  INVX1 G47816 (.I(W10250), .ZN(W11726));
  INVX1 G47817 (.I(W22214), .ZN(O9994));
  INVX1 G47818 (.I(W3709), .ZN(W11727));
  INVX1 G47819 (.I(W6587), .ZN(W11731));
  INVX1 G47820 (.I(W10041), .ZN(O534));
  INVX1 G47821 (.I(W11614), .ZN(W11735));
  INVX1 G47822 (.I(W2868), .ZN(W11841));
  INVX1 G47823 (.I(W7138), .ZN(W11811));
  INVX1 G47824 (.I(W3048), .ZN(W39049));
  INVX1 G47825 (.I(W9002), .ZN(W11821));
  INVX1 G47826 (.I(I439), .ZN(W11824));
  INVX1 G47827 (.I(I79), .ZN(O9934));
  INVX1 G47828 (.I(W26814), .ZN(W39040));
  INVX1 G47829 (.I(W10874), .ZN(O541));
  INVX1 G47830 (.I(W20080), .ZN(W39038));
  INVX1 G47831 (.I(W7989), .ZN(W11834));
  INVX1 G47832 (.I(W36037), .ZN(W39052));
  INVX1 G47833 (.I(W11768), .ZN(O9930));
  INVX1 G47834 (.I(W5533), .ZN(W11843));
  INVX1 G47835 (.I(I1614), .ZN(O9929));
  INVX1 G47836 (.I(W14609), .ZN(W39028));
  INVX1 G47837 (.I(W11331), .ZN(W11845));
  INVX1 G47838 (.I(W32315), .ZN(W39023));
  INVX1 G47839 (.I(W78), .ZN(W11852));
  INVX1 G47840 (.I(W24221), .ZN(O9926));
  INVX1 G47841 (.I(W197), .ZN(W11853));
  INVX1 G47842 (.I(I202), .ZN(W11791));
  INVX1 G47843 (.I(W11691), .ZN(O9961));
  INVX1 G47844 (.I(W2583), .ZN(W11774));
  INVX1 G47845 (.I(W25286), .ZN(W39079));
  INVX1 G47846 (.I(W6547), .ZN(W11778));
  INVX1 G47847 (.I(W27404), .ZN(O9957));
  INVX1 G47848 (.I(W553), .ZN(O9956));
  INVX1 G47849 (.I(W9243), .ZN(W11779));
  INVX1 G47850 (.I(W4654), .ZN(W11785));
  INVX1 G47851 (.I(W560), .ZN(W11787));
  INVX1 G47852 (.I(W6973), .ZN(W11702));
  INVX1 G47853 (.I(W10056), .ZN(W11792));
  INVX1 G47854 (.I(W13363), .ZN(O9948));
  INVX1 G47855 (.I(W6895), .ZN(W11793));
  INVX1 G47856 (.I(W2108), .ZN(W39061));
  INVX1 G47857 (.I(W25028), .ZN(O9945));
  INVX1 G47858 (.I(W1707), .ZN(W11802));
  INVX1 G47859 (.I(W37567), .ZN(O9942));
  INVX1 G47860 (.I(W1464), .ZN(W11803));
  INVX1 G47861 (.I(I530), .ZN(W11806));
  INVX1 G47862 (.I(W2973), .ZN(W11614));
  INVX1 G47863 (.I(W10782), .ZN(W11603));
  INVX1 G47864 (.I(W1441), .ZN(O10078));
  INVX1 G47865 (.I(W239), .ZN(W11606));
  INVX1 G47866 (.I(W393), .ZN(O10074));
  INVX1 G47867 (.I(W12562), .ZN(O10073));
  INVX1 G47868 (.I(W34559), .ZN(O10072));
  INVX1 G47869 (.I(W30547), .ZN(O10070));
  INVX1 G47870 (.I(W6500), .ZN(W11612));
  INVX1 G47871 (.I(W1137), .ZN(W11613));
  INVX1 G47872 (.I(W33527), .ZN(W39251));
  INVX1 G47873 (.I(W35236), .ZN(O10068));
  INVX1 G47874 (.I(I1514), .ZN(W39229));
  INVX1 G47875 (.I(W4114), .ZN(O10066));
  INVX1 G47876 (.I(W2559), .ZN(W11617));
  INVX1 G47877 (.I(W3412), .ZN(W11622));
  INVX1 G47878 (.I(W4457), .ZN(O10061));
  INVX1 G47879 (.I(I1159), .ZN(W11625));
  INVX1 G47880 (.I(W1416), .ZN(W11627));
  INVX1 G47881 (.I(W36415), .ZN(O10054));
  INVX1 G47882 (.I(W1742), .ZN(W11588));
  INVX1 G47883 (.I(W9245), .ZN(O10097));
  INVX1 G47884 (.I(W22984), .ZN(W39276));
  INVX1 G47885 (.I(W13036), .ZN(W39275));
  INVX1 G47886 (.I(W3925), .ZN(W11573));
  INVX1 G47887 (.I(W3731), .ZN(W11575));
  INVX1 G47888 (.I(W31331), .ZN(O10091));
  INVX1 G47889 (.I(I1814), .ZN(W11583));
  INVX1 G47890 (.I(W6199), .ZN(W11585));
  INVX1 G47891 (.I(W9336), .ZN(W11587));
  INVX1 G47892 (.I(W32294), .ZN(O10053));
  INVX1 G47893 (.I(W3752), .ZN(W11589));
  INVX1 G47894 (.I(W3412), .ZN(W11591));
  INVX1 G47895 (.I(W6159), .ZN(W11593));
  INVX1 G47896 (.I(W25325), .ZN(W39258));
  INVX1 G47897 (.I(W4536), .ZN(W11595));
  INVX1 G47898 (.I(W2549), .ZN(W11596));
  INVX1 G47899 (.I(W8797), .ZN(O523));
  INVX1 G47900 (.I(W35787), .ZN(O10084));
  INVX1 G47901 (.I(W36650), .ZN(O10083));
  INVX1 G47902 (.I(W5453), .ZN(O10022));
  INVX1 G47903 (.I(W25976), .ZN(O10034));
  INVX1 G47904 (.I(I1336), .ZN(O529));
  INVX1 G47905 (.I(W8665), .ZN(W11671));
  INVX1 G47906 (.I(W876), .ZN(W11676));
  INVX1 G47907 (.I(W5902), .ZN(W11677));
  INVX1 G47908 (.I(W4638), .ZN(O10028));
  INVX1 G47909 (.I(W9215), .ZN(W11679));
  INVX1 G47910 (.I(W1338), .ZN(W11682));
  INVX1 G47911 (.I(W9624), .ZN(W11687));
  INVX1 G47912 (.I(W31888), .ZN(W39183));
  INVX1 G47913 (.I(W36211), .ZN(O10021));
  INVX1 G47914 (.I(W20234), .ZN(O10020));
  INVX1 G47915 (.I(W5277), .ZN(O10018));
  INVX1 G47916 (.I(W3187), .ZN(O10017));
  INVX1 G47917 (.I(W7000), .ZN(W11689));
  INVX1 G47918 (.I(W307), .ZN(W11695));
  INVX1 G47919 (.I(W1742), .ZN(W11698));
  INVX1 G47920 (.I(W6761), .ZN(W11700));
  INVX1 G47921 (.I(W28546), .ZN(O10012));
  INVX1 G47922 (.I(W4370), .ZN(O10044));
  INVX1 G47923 (.I(W20169), .ZN(O10051));
  INVX1 G47924 (.I(W7325), .ZN(W11634));
  INVX1 G47925 (.I(W31057), .ZN(O10050));
  INVX1 G47926 (.I(W2674), .ZN(W39206));
  INVX1 G47927 (.I(W6007), .ZN(W11636));
  INVX1 G47928 (.I(W38), .ZN(W11637));
  INVX1 G47929 (.I(I1700), .ZN(W11643));
  INVX1 G47930 (.I(W27578), .ZN(O10046));
  INVX1 G47931 (.I(W8020), .ZN(W11648));
  INVX1 G47932 (.I(W5102), .ZN(W11855));
  INVX1 G47933 (.I(W2739), .ZN(O10043));
  INVX1 G47934 (.I(W2799), .ZN(W11652));
  INVX1 G47935 (.I(W7619), .ZN(W11657));
  INVX1 G47936 (.I(W572), .ZN(W11658));
  INVX1 G47937 (.I(W2081), .ZN(O10039));
  INVX1 G47938 (.I(W22138), .ZN(O10038));
  INVX1 G47939 (.I(W365), .ZN(O528));
  INVX1 G47940 (.I(W2690), .ZN(W11665));
  INVX1 G47941 (.I(W9395), .ZN(W11668));
  INVX1 G47942 (.I(W11130), .ZN(W12007));
  INVX1 G47943 (.I(I552), .ZN(W11993));
  INVX1 G47944 (.I(W35030), .ZN(W38868));
  INVX1 G47945 (.I(W32562), .ZN(O9837));
  INVX1 G47946 (.I(W11498), .ZN(O9836));
  INVX1 G47947 (.I(W13), .ZN(W12000));
  INVX1 G47948 (.I(W18245), .ZN(W38862));
  INVX1 G47949 (.I(W5808), .ZN(O556));
  INVX1 G47950 (.I(W21455), .ZN(O9832));
  INVX1 G47951 (.I(W4125), .ZN(W12004));
  INVX1 G47952 (.I(W263), .ZN(W12005));
  INVX1 G47953 (.I(I1298), .ZN(W11992));
  INVX1 G47954 (.I(W3317), .ZN(W12008));
  INVX1 G47955 (.I(W15229), .ZN(O9828));
  INVX1 G47956 (.I(W11908), .ZN(W12014));
  INVX1 G47957 (.I(W3591), .ZN(O9826));
  INVX1 G47958 (.I(I1284), .ZN(W12016));
  INVX1 G47959 (.I(W24484), .ZN(O9823));
  INVX1 G47960 (.I(W11278), .ZN(W12021));
  INVX1 G47961 (.I(W17022), .ZN(W38843));
  INVX1 G47962 (.I(W6155), .ZN(O561));
  INVX1 G47963 (.I(I604), .ZN(W11981));
  INVX1 G47964 (.I(W3627), .ZN(W11972));
  INVX1 G47965 (.I(W36798), .ZN(O9851));
  INVX1 G47966 (.I(W15933), .ZN(O9850));
  INVX1 G47967 (.I(W11262), .ZN(W11973));
  INVX1 G47968 (.I(W21594), .ZN(O9849));
  INVX1 G47969 (.I(W7557), .ZN(W11975));
  INVX1 G47970 (.I(W4874), .ZN(W11978));
  INVX1 G47971 (.I(W2729), .ZN(W11979));
  INVX1 G47972 (.I(W1944), .ZN(O9846));
  INVX1 G47973 (.I(W4826), .ZN(W12027));
  INVX1 G47974 (.I(W4927), .ZN(W11982));
  INVX1 G47975 (.I(W1661), .ZN(O555));
  INVX1 G47976 (.I(W3038), .ZN(W38882));
  INVX1 G47977 (.I(W25401), .ZN(O9842));
  INVX1 G47978 (.I(W761), .ZN(W11987));
  INVX1 G47979 (.I(W11467), .ZN(W11989));
  INVX1 G47980 (.I(W8853), .ZN(W11990));
  INVX1 G47981 (.I(W4927), .ZN(O9840));
  INVX1 G47982 (.I(W10208), .ZN(W38873));
  INVX1 G47983 (.I(W5129), .ZN(O9793));
  INVX1 G47984 (.I(W8250), .ZN(W12046));
  INVX1 G47985 (.I(W33172), .ZN(W38806));
  INVX1 G47986 (.I(W8801), .ZN(W12049));
  INVX1 G47987 (.I(W9028), .ZN(O564));
  INVX1 G47988 (.I(W25933), .ZN(O9797));
  INVX1 G47989 (.I(W1872), .ZN(W12052));
  INVX1 G47990 (.I(W8768), .ZN(W12054));
  INVX1 G47991 (.I(W6152), .ZN(O9794));
  INVX1 G47992 (.I(W25073), .ZN(W38798));
  INVX1 G47993 (.I(W27628), .ZN(O9800));
  INVX1 G47994 (.I(W11867), .ZN(W38796));
  INVX1 G47995 (.I(W9453), .ZN(W12055));
  INVX1 G47996 (.I(W9256), .ZN(W12056));
  INVX1 G47997 (.I(W10925), .ZN(W12061));
  INVX1 G47998 (.I(W4806), .ZN(W12063));
  INVX1 G47999 (.I(W22622), .ZN(W38789));
  INVX1 G48000 (.I(W6643), .ZN(W12064));
  INVX1 G48001 (.I(W18544), .ZN(O9786));
  INVX1 G48002 (.I(W11827), .ZN(W12068));
  INVX1 G48003 (.I(I647), .ZN(W12034));
  INVX1 G48004 (.I(W7542), .ZN(O562));
  INVX1 G48005 (.I(W36405), .ZN(O9815));
  INVX1 G48006 (.I(W16330), .ZN(O9814));
  INVX1 G48007 (.I(W33876), .ZN(W38831));
  INVX1 G48008 (.I(W5350), .ZN(O9813));
  INVX1 G48009 (.I(W35475), .ZN(O9812));
  INVX1 G48010 (.I(W11381), .ZN(W12033));
  INVX1 G48011 (.I(W37421), .ZN(O9810));
  INVX1 G48012 (.I(W31447), .ZN(W38825));
  INVX1 G48013 (.I(W766), .ZN(W11971));
  INVX1 G48014 (.I(W4110), .ZN(W12035));
  INVX1 G48015 (.I(W34624), .ZN(W38822));
  INVX1 G48016 (.I(W32733), .ZN(O9807));
  INVX1 G48017 (.I(W178), .ZN(W12039));
  INVX1 G48018 (.I(W23892), .ZN(O9806));
  INVX1 G48019 (.I(W910), .ZN(O563));
  INVX1 G48020 (.I(W10550), .ZN(W38814));
  INVX1 G48021 (.I(W14654), .ZN(O9804));
  INVX1 G48022 (.I(W21730), .ZN(O9802));
  INVX1 G48023 (.I(W9345), .ZN(W11910));
  INVX1 G48024 (.I(W10386), .ZN(W11897));
  INVX1 G48025 (.I(W31221), .ZN(W38986));
  INVX1 G48026 (.I(W18075), .ZN(O9905));
  INVX1 G48027 (.I(W6984), .ZN(O9904));
  INVX1 G48028 (.I(I1307), .ZN(W11900));
  INVX1 G48029 (.I(W16729), .ZN(O9903));
  INVX1 G48030 (.I(I1780), .ZN(W11903));
  INVX1 G48031 (.I(W1667), .ZN(O547));
  INVX1 G48032 (.I(W33016), .ZN(W38973));
  INVX1 G48033 (.I(W10986), .ZN(W11893));
  INVX1 G48034 (.I(W23717), .ZN(W38970));
  INVX1 G48035 (.I(W6825), .ZN(O9894));
  INVX1 G48036 (.I(W26776), .ZN(O9892));
  INVX1 G48037 (.I(W23944), .ZN(O9891));
  INVX1 G48038 (.I(W27224), .ZN(W38963));
  INVX1 G48039 (.I(W10782), .ZN(W11917));
  INVX1 G48040 (.I(W33031), .ZN(O9890));
  INVX1 G48041 (.I(W19300), .ZN(W38959));
  INVX1 G48042 (.I(W34641), .ZN(W38958));
  INVX1 G48043 (.I(W4311), .ZN(W11872));
  INVX1 G48044 (.I(I450), .ZN(W11856));
  INVX1 G48045 (.I(W11222), .ZN(W11858));
  INVX1 G48046 (.I(W21160), .ZN(O9921));
  INVX1 G48047 (.I(W3031), .ZN(W11860));
  INVX1 G48048 (.I(W25685), .ZN(W39010));
  INVX1 G48049 (.I(W29099), .ZN(O9919));
  INVX1 G48050 (.I(I819), .ZN(W11866));
  INVX1 G48051 (.I(I1618), .ZN(W11869));
  INVX1 G48052 (.I(W21687), .ZN(O9915));
  INVX1 G48053 (.I(W10746), .ZN(W38957));
  INVX1 G48054 (.I(W623), .ZN(W11875));
  INVX1 G48055 (.I(W6153), .ZN(W11877));
  INVX1 G48056 (.I(W135), .ZN(W11881));
  INVX1 G48057 (.I(W3374), .ZN(O9911));
  INVX1 G48058 (.I(W19468), .ZN(W38996));
  INVX1 G48059 (.I(W7815), .ZN(O545));
  INVX1 G48060 (.I(W27218), .ZN(W38993));
  INVX1 G48061 (.I(W8970), .ZN(W11890));
  INVX1 G48062 (.I(W15118), .ZN(O9909));
  INVX1 G48063 (.I(W2595), .ZN(W11955));
  INVX1 G48064 (.I(W32595), .ZN(O9867));
  INVX1 G48065 (.I(W3801), .ZN(W38926));
  INVX1 G48066 (.I(W9214), .ZN(W11946));
  INVX1 G48067 (.I(W13033), .ZN(W38922));
  INVX1 G48068 (.I(W3932), .ZN(W11948));
  INVX1 G48069 (.I(W33826), .ZN(W38920));
  INVX1 G48070 (.I(W20313), .ZN(O9863));
  INVX1 G48071 (.I(W21811), .ZN(O9862));
  INVX1 G48072 (.I(W2421), .ZN(W38913));
  INVX1 G48073 (.I(W8406), .ZN(O9869));
  INVX1 G48074 (.I(W13842), .ZN(O9860));
  INVX1 G48075 (.I(W3057), .ZN(W11959));
  INVX1 G48076 (.I(W5189), .ZN(W11960));
  INVX1 G48077 (.I(W8489), .ZN(W11962));
  INVX1 G48078 (.I(W8646), .ZN(W11963));
  INVX1 G48079 (.I(W35685), .ZN(O9856));
  INVX1 G48080 (.I(W4285), .ZN(O553));
  INVX1 G48081 (.I(I1014), .ZN(W11967));
  INVX1 G48082 (.I(W10002), .ZN(W11968));
  INVX1 G48083 (.I(W36252), .ZN(O9880));
  INVX1 G48084 (.I(W34114), .ZN(O9889));
  INVX1 G48085 (.I(W7066), .ZN(W11925));
  INVX1 G48086 (.I(W10735), .ZN(W11926));
  INVX1 G48087 (.I(W1422), .ZN(W11928));
  INVX1 G48088 (.I(W1165), .ZN(W11929));
  INVX1 G48089 (.I(W20020), .ZN(O9885));
  INVX1 G48090 (.I(W20961), .ZN(O9883));
  INVX1 G48091 (.I(W17626), .ZN(O9882));
  INVX1 G48092 (.I(W33121), .ZN(W38944));
  INVX1 G48093 (.I(W2413), .ZN(O10098));
  INVX1 G48094 (.I(W2728), .ZN(O9879));
  INVX1 G48095 (.I(W28002), .ZN(O9878));
  INVX1 G48096 (.I(W8054), .ZN(W11934));
  INVX1 G48097 (.I(W26781), .ZN(O9877));
  INVX1 G48098 (.I(W38260), .ZN(O9875));
  INVX1 G48099 (.I(W6438), .ZN(O9874));
  INVX1 G48100 (.I(W2641), .ZN(W11938));
  INVX1 G48101 (.I(W1404), .ZN(W11940));
  INVX1 G48102 (.I(W2727), .ZN(W38932));
  INVX1 G48103 (.I(W10268), .ZN(W11288));
  INVX1 G48104 (.I(W8101), .ZN(W11262));
  INVX1 G48105 (.I(W2761), .ZN(W11264));
  INVX1 G48106 (.I(W7908), .ZN(W11268));
  INVX1 G48107 (.I(I622), .ZN(W11271));
  INVX1 G48108 (.I(W8142), .ZN(W11273));
  INVX1 G48109 (.I(W25957), .ZN(O10320));
  INVX1 G48110 (.I(W10204), .ZN(O10319));
  INVX1 G48111 (.I(W10640), .ZN(W11279));
  INVX1 G48112 (.I(W8009), .ZN(O10314));
  INVX1 G48113 (.I(W5552), .ZN(W11283));
  INVX1 G48114 (.I(W7659), .ZN(W11261));
  INVX1 G48115 (.I(W10739), .ZN(W11289));
  INVX1 G48116 (.I(I366), .ZN(W11290));
  INVX1 G48117 (.I(I6), .ZN(W11291));
  INVX1 G48118 (.I(W30032), .ZN(O10308));
  INVX1 G48119 (.I(W33325), .ZN(W39581));
  INVX1 G48120 (.I(W2695), .ZN(O10306));
  INVX1 G48121 (.I(W34968), .ZN(O10305));
  INVX1 G48122 (.I(I1401), .ZN(O10304));
  INVX1 G48123 (.I(W7906), .ZN(O10303));
  INVX1 G48124 (.I(W1190), .ZN(W11248));
  INVX1 G48125 (.I(W33679), .ZN(O10348));
  INVX1 G48126 (.I(W32764), .ZN(O10346));
  INVX1 G48127 (.I(W22439), .ZN(O10345));
  INVX1 G48128 (.I(W50), .ZN(W11238));
  INVX1 G48129 (.I(W4981), .ZN(W39629));
  INVX1 G48130 (.I(W2185), .ZN(W11239));
  INVX1 G48131 (.I(W331), .ZN(W11240));
  INVX1 G48132 (.I(W824), .ZN(W11242));
  INVX1 G48133 (.I(W13816), .ZN(O10337));
  INVX1 G48134 (.I(W4376), .ZN(W11294));
  INVX1 G48135 (.I(W34579), .ZN(W39619));
  INVX1 G48136 (.I(W3350), .ZN(W11249));
  INVX1 G48137 (.I(W8613), .ZN(W11250));
  INVX1 G48138 (.I(W22785), .ZN(W39616));
  INVX1 G48139 (.I(W36435), .ZN(O10334));
  INVX1 G48140 (.I(W2708), .ZN(W11254));
  INVX1 G48141 (.I(I20), .ZN(O494));
  INVX1 G48142 (.I(W9181), .ZN(O495));
  INVX1 G48143 (.I(W2070), .ZN(W11260));
  INVX1 G48144 (.I(W4557), .ZN(W11335));
  INVX1 G48145 (.I(W6366), .ZN(W11320));
  INVX1 G48146 (.I(I1100), .ZN(W11321));
  INVX1 G48147 (.I(W20916), .ZN(W39545));
  INVX1 G48148 (.I(W10546), .ZN(O10283));
  INVX1 G48149 (.I(W11313), .ZN(W11323));
  INVX1 G48150 (.I(W27481), .ZN(O10279));
  INVX1 G48151 (.I(W8163), .ZN(W39536));
  INVX1 G48152 (.I(W3960), .ZN(W11332));
  INVX1 G48153 (.I(W177), .ZN(O10275));
  INVX1 G48154 (.I(W10444), .ZN(O10286));
  INVX1 G48155 (.I(W1282), .ZN(O10271));
  INVX1 G48156 (.I(W6431), .ZN(W11338));
  INVX1 G48157 (.I(W6849), .ZN(W11339));
  INVX1 G48158 (.I(W32776), .ZN(W39525));
  INVX1 G48159 (.I(W36645), .ZN(O10269));
  INVX1 G48160 (.I(W17606), .ZN(O10268));
  INVX1 G48161 (.I(W27546), .ZN(O10266));
  INVX1 G48162 (.I(W9303), .ZN(W11343));
  INVX1 G48163 (.I(I1337), .ZN(O10264));
  INVX1 G48164 (.I(W8771), .ZN(O499));
  INVX1 G48165 (.I(I1440), .ZN(W11295));
  INVX1 G48166 (.I(W10154), .ZN(W11296));
  INVX1 G48167 (.I(W32138), .ZN(O10300));
  INVX1 G48168 (.I(W8205), .ZN(W11300));
  INVX1 G48169 (.I(W9320), .ZN(O10298));
  INVX1 G48170 (.I(W4794), .ZN(W11301));
  INVX1 G48171 (.I(W4902), .ZN(W11302));
  INVX1 G48172 (.I(W7096), .ZN(W11303));
  INVX1 G48173 (.I(W7729), .ZN(W11304));
  INVX1 G48174 (.I(W14737), .ZN(W39635));
  INVX1 G48175 (.I(W3562), .ZN(W11309));
  INVX1 G48176 (.I(W626), .ZN(W11310));
  INVX1 G48177 (.I(W7778), .ZN(W11312));
  INVX1 G48178 (.I(W4752), .ZN(W11314));
  INVX1 G48179 (.I(W9044), .ZN(W11315));
  INVX1 G48180 (.I(W36196), .ZN(O10288));
  INVX1 G48181 (.I(W7682), .ZN(W39552));
  INVX1 G48182 (.I(W10255), .ZN(O10287));
  INVX1 G48183 (.I(W9549), .ZN(W11318));
  INVX1 G48184 (.I(W7643), .ZN(W11173));
  INVX1 G48185 (.I(W6910), .ZN(W11151));
  INVX1 G48186 (.I(W28248), .ZN(W39705));
  INVX1 G48187 (.I(I884), .ZN(W11158));
  INVX1 G48188 (.I(W4487), .ZN(W11159));
  INVX1 G48189 (.I(W2610), .ZN(W11164));
  INVX1 G48190 (.I(W6734), .ZN(W11165));
  INVX1 G48191 (.I(W4072), .ZN(O10388));
  INVX1 G48192 (.I(W2647), .ZN(W11167));
  INVX1 G48193 (.I(W35140), .ZN(W39695));
  INVX1 G48194 (.I(W1108), .ZN(O485));
  INVX1 G48195 (.I(W5802), .ZN(W11176));
  INVX1 G48196 (.I(W7834), .ZN(W11184));
  INVX1 G48197 (.I(W28762), .ZN(O10382));
  INVX1 G48198 (.I(W998), .ZN(W11185));
  INVX1 G48199 (.I(W8384), .ZN(W11187));
  INVX1 G48200 (.I(W9866), .ZN(W11192));
  INVX1 G48201 (.I(W1874), .ZN(W11193));
  INVX1 G48202 (.I(W12266), .ZN(O10378));
  INVX1 G48203 (.I(W10488), .ZN(W11195));
  INVX1 G48204 (.I(I796), .ZN(O10406));
  INVX1 G48205 (.I(W14696), .ZN(W39734));
  INVX1 G48206 (.I(W6238), .ZN(W11135));
  INVX1 G48207 (.I(W31269), .ZN(O10409));
  INVX1 G48208 (.I(W5748), .ZN(W11136));
  INVX1 G48209 (.I(W27393), .ZN(O10408));
  INVX1 G48210 (.I(W37706), .ZN(W39726));
  INVX1 G48211 (.I(W8750), .ZN(W11137));
  INVX1 G48212 (.I(W11313), .ZN(W39724));
  INVX1 G48213 (.I(W32210), .ZN(O10407));
  INVX1 G48214 (.I(W6715), .ZN(W11198));
  INVX1 G48215 (.I(W13966), .ZN(O10405));
  INVX1 G48216 (.I(W17366), .ZN(W39719));
  INVX1 G48217 (.I(W30374), .ZN(O10404));
  INVX1 G48218 (.I(I1389), .ZN(W11140));
  INVX1 G48219 (.I(W12412), .ZN(O10402));
  INVX1 G48220 (.I(W14819), .ZN(O10401));
  INVX1 G48221 (.I(W4714), .ZN(W11145));
  INVX1 G48222 (.I(W9060), .ZN(W11146));
  INVX1 G48223 (.I(W16362), .ZN(O10397));
  INVX1 G48224 (.I(W22107), .ZN(O10355));
  INVX1 G48225 (.I(W2854), .ZN(W11217));
  INVX1 G48226 (.I(W25334), .ZN(W39655));
  INVX1 G48227 (.I(W10727), .ZN(W11218));
  INVX1 G48228 (.I(W26203), .ZN(O10359));
  INVX1 G48229 (.I(W5437), .ZN(W11219));
  INVX1 G48230 (.I(W858), .ZN(O10358));
  INVX1 G48231 (.I(W1443), .ZN(W11224));
  INVX1 G48232 (.I(W28947), .ZN(O10356));
  INVX1 G48233 (.I(W38469), .ZN(W39648));
  INVX1 G48234 (.I(W14590), .ZN(O10362));
  INVX1 G48235 (.I(I62), .ZN(W11225));
  INVX1 G48236 (.I(W4965), .ZN(W11228));
  INVX1 G48237 (.I(I1982), .ZN(O489));
  INVX1 G48238 (.I(W21926), .ZN(O10352));
  INVX1 G48239 (.I(W31318), .ZN(O10351));
  INVX1 G48240 (.I(W6136), .ZN(O10350));
  INVX1 G48241 (.I(W3193), .ZN(W11234));
  INVX1 G48242 (.I(W25613), .ZN(W39637));
  INVX1 G48243 (.I(W7936), .ZN(O490));
  INVX1 G48244 (.I(W7987), .ZN(W11210));
  INVX1 G48245 (.I(W5578), .ZN(O10376));
  INVX1 G48246 (.I(W27826), .ZN(O10374));
  INVX1 G48247 (.I(W3130), .ZN(W11204));
  INVX1 G48248 (.I(W8616), .ZN(W11205));
  INVX1 G48249 (.I(W5683), .ZN(W11206));
  INVX1 G48250 (.I(W3194), .ZN(W11207));
  INVX1 G48251 (.I(I1756), .ZN(W11208));
  INVX1 G48252 (.I(W4150), .ZN(W11209));
  INVX1 G48253 (.I(W17795), .ZN(O10369));
  INVX1 G48254 (.I(W11300), .ZN(W11347));
  INVX1 G48255 (.I(W32854), .ZN(W39666));
  INVX1 G48256 (.I(W22995), .ZN(O10368));
  INVX1 G48257 (.I(W631), .ZN(W11211));
  INVX1 G48258 (.I(W30509), .ZN(O10366));
  INVX1 G48259 (.I(W37553), .ZN(O10365));
  INVX1 G48260 (.I(W10388), .ZN(W11212));
  INVX1 G48261 (.I(W6202), .ZN(W11214));
  INVX1 G48262 (.I(W25355), .ZN(O10364));
  INVX1 G48263 (.I(W8877), .ZN(W11215));
  INVX1 G48264 (.I(W11201), .ZN(W11501));
  INVX1 G48265 (.I(W19333), .ZN(O10159));
  INVX1 G48266 (.I(W27388), .ZN(O10157));
  INVX1 G48267 (.I(W1674), .ZN(O10156));
  INVX1 G48268 (.I(W36484), .ZN(O10155));
  INVX1 G48269 (.I(W8497), .ZN(W11485));
  INVX1 G48270 (.I(W8346), .ZN(W11489));
  INVX1 G48271 (.I(W3550), .ZN(W39359));
  INVX1 G48272 (.I(W6799), .ZN(W11494));
  INVX1 G48273 (.I(W4273), .ZN(W11499));
  INVX1 G48274 (.I(W9318), .ZN(W39353));
  INVX1 G48275 (.I(W4263), .ZN(W11481));
  INVX1 G48276 (.I(W22360), .ZN(O10143));
  INVX1 G48277 (.I(W7904), .ZN(W39349));
  INVX1 G48278 (.I(W9747), .ZN(O10141));
  INVX1 G48279 (.I(W8271), .ZN(W11504));
  INVX1 G48280 (.I(W10997), .ZN(W11506));
  INVX1 G48281 (.I(W1630), .ZN(W11507));
  INVX1 G48282 (.I(W37850), .ZN(O10138));
  INVX1 G48283 (.I(W11292), .ZN(W11509));
  INVX1 G48284 (.I(W553), .ZN(O10137));
  INVX1 G48285 (.I(W6061), .ZN(W11457));
  INVX1 G48286 (.I(W38844), .ZN(O10182));
  INVX1 G48287 (.I(W6555), .ZN(W11452));
  INVX1 G48288 (.I(W10962), .ZN(W39398));
  INVX1 G48289 (.I(W6307), .ZN(W39397));
  INVX1 G48290 (.I(W36718), .ZN(W39396));
  INVX1 G48291 (.I(W4854), .ZN(O10179));
  INVX1 G48292 (.I(W5833), .ZN(W11454));
  INVX1 G48293 (.I(W10836), .ZN(O10178));
  INVX1 G48294 (.I(W8636), .ZN(W11455));
  INVX1 G48295 (.I(W21625), .ZN(O10136));
  INVX1 G48296 (.I(W33704), .ZN(O10174));
  INVX1 G48297 (.I(W35929), .ZN(O10173));
  INVX1 G48298 (.I(W8107), .ZN(O10170));
  INVX1 G48299 (.I(W13417), .ZN(O10169));
  INVX1 G48300 (.I(W23518), .ZN(W39382));
  INVX1 G48301 (.I(W7552), .ZN(W11472));
  INVX1 G48302 (.I(W7833), .ZN(W11473));
  INVX1 G48303 (.I(W26831), .ZN(O10162));
  INVX1 G48304 (.I(W7557), .ZN(W11479));
  INVX1 G48305 (.I(W2909), .ZN(W11547));
  INVX1 G48306 (.I(W30231), .ZN(O10118));
  INVX1 G48307 (.I(I1998), .ZN(W11529));
  INVX1 G48308 (.I(W6484), .ZN(O516));
  INVX1 G48309 (.I(W7100), .ZN(W11537));
  INVX1 G48310 (.I(W7192), .ZN(W11539));
  INVX1 G48311 (.I(W30529), .ZN(O10112));
  INVX1 G48312 (.I(W3543), .ZN(W11540));
  INVX1 G48313 (.I(W38352), .ZN(O10110));
  INVX1 G48314 (.I(W719), .ZN(O10109));
  INVX1 G48315 (.I(W32532), .ZN(W39312));
  INVX1 G48316 (.I(W5273), .ZN(O518));
  INVX1 G48317 (.I(W24248), .ZN(O10105));
  INVX1 G48318 (.I(W7786), .ZN(O10104));
  INVX1 G48319 (.I(W9543), .ZN(W11556));
  INVX1 G48320 (.I(W1630), .ZN(W39285));
  INVX1 G48321 (.I(W3862), .ZN(W11561));
  INVX1 G48322 (.I(W752), .ZN(W11565));
  INVX1 G48323 (.I(W7993), .ZN(W11566));
  INVX1 G48324 (.I(W15291), .ZN(W39280));
  INVX1 G48325 (.I(W9177), .ZN(W11518));
  INVX1 G48326 (.I(W7876), .ZN(W11510));
  INVX1 G48327 (.I(W34453), .ZN(W39336));
  INVX1 G48328 (.I(W32983), .ZN(W39335));
  INVX1 G48329 (.I(W3611), .ZN(O10133));
  INVX1 G48330 (.I(W5425), .ZN(W11512));
  INVX1 G48331 (.I(I340), .ZN(O10131));
  INVX1 G48332 (.I(W22733), .ZN(O10129));
  INVX1 G48333 (.I(I668), .ZN(W11516));
  INVX1 G48334 (.I(W5872), .ZN(O10127));
  INVX1 G48335 (.I(W5481), .ZN(O511));
  INVX1 G48336 (.I(W35986), .ZN(O10125));
  INVX1 G48337 (.I(W1625), .ZN(O10124));
  INVX1 G48338 (.I(W1710), .ZN(O10123));
  INVX1 G48339 (.I(W2764), .ZN(W11523));
  INVX1 G48340 (.I(I1748), .ZN(W11525));
  INVX1 G48341 (.I(W8757), .ZN(O10121));
  INVX1 G48342 (.I(W1334), .ZN(W11526));
  INVX1 G48343 (.I(W797), .ZN(O10119));
  INVX1 G48344 (.I(W889), .ZN(W39315));
  INVX1 G48345 (.I(W1242), .ZN(W11390));
  INVX1 G48346 (.I(W15972), .ZN(O10244));
  INVX1 G48347 (.I(W5334), .ZN(W11371));
  INVX1 G48348 (.I(W9116), .ZN(O10243));
  INVX1 G48349 (.I(W8309), .ZN(W11373));
  INVX1 G48350 (.I(W2597), .ZN(W11374));
  INVX1 G48351 (.I(W4417), .ZN(W11383));
  INVX1 G48352 (.I(W8044), .ZN(O10237));
  INVX1 G48353 (.I(W34367), .ZN(W39476));
  INVX1 G48354 (.I(W524), .ZN(W11389));
  INVX1 G48355 (.I(W3493), .ZN(W11370));
  INVX1 G48356 (.I(I1820), .ZN(W11394));
  INVX1 G48357 (.I(W32254), .ZN(W39469));
  INVX1 G48358 (.I(I1738), .ZN(W11397));
  INVX1 G48359 (.I(W7475), .ZN(W11398));
  INVX1 G48360 (.I(W12459), .ZN(O10227));
  INVX1 G48361 (.I(W5203), .ZN(O10226));
  INVX1 G48362 (.I(W16298), .ZN(O10225));
  INVX1 G48363 (.I(W11809), .ZN(O10224));
  INVX1 G48364 (.I(I1876), .ZN(W39460));
  INVX1 G48365 (.I(W6920), .ZN(W39503));
  INVX1 G48366 (.I(W14611), .ZN(O10261));
  INVX1 G48367 (.I(W3030), .ZN(W11349));
  INVX1 G48368 (.I(W5837), .ZN(O502));
  INVX1 G48369 (.I(W29243), .ZN(W39511));
  INVX1 G48370 (.I(W8060), .ZN(W11353));
  INVX1 G48371 (.I(W788), .ZN(W11358));
  INVX1 G48372 (.I(W3515), .ZN(W39508));
  INVX1 G48373 (.I(W33206), .ZN(O10256));
  INVX1 G48374 (.I(W672), .ZN(W11361));
  INVX1 G48375 (.I(W9406), .ZN(W11399));
  INVX1 G48376 (.I(W25390), .ZN(O10254));
  INVX1 G48377 (.I(W7100), .ZN(W11365));
  INVX1 G48378 (.I(W21756), .ZN(O10252));
  INVX1 G48379 (.I(W12354), .ZN(O10251));
  INVX1 G48380 (.I(I241), .ZN(W11366));
  INVX1 G48381 (.I(W3271), .ZN(O10249));
  INVX1 G48382 (.I(W26083), .ZN(O10247));
  INVX1 G48383 (.I(W9812), .ZN(W11369));
  INVX1 G48384 (.I(W32705), .ZN(O10245));
  INVX1 G48385 (.I(W2387), .ZN(W11437));
  INVX1 G48386 (.I(W508), .ZN(W39427));
  INVX1 G48387 (.I(W31133), .ZN(W39426));
  INVX1 G48388 (.I(W20756), .ZN(O10198));
  INVX1 G48389 (.I(W32408), .ZN(O10197));
  INVX1 G48390 (.I(W21516), .ZN(O10196));
  INVX1 G48391 (.I(W38075), .ZN(W39421));
  INVX1 G48392 (.I(W10848), .ZN(W11432));
  INVX1 G48393 (.I(W5654), .ZN(W11435));
  INVX1 G48394 (.I(W22710), .ZN(W39417));
  INVX1 G48395 (.I(W9603), .ZN(W11428));
  INVX1 G48396 (.I(W1762), .ZN(W11440));
  INVX1 G48397 (.I(W31581), .ZN(O10191));
  INVX1 G48398 (.I(W9329), .ZN(W11441));
  INVX1 G48399 (.I(W15959), .ZN(O10189));
  INVX1 G48400 (.I(W9424), .ZN(W11442));
  INVX1 G48401 (.I(W2552), .ZN(O10187));
  INVX1 G48402 (.I(W10936), .ZN(W11443));
  INVX1 G48403 (.I(W24134), .ZN(O10186));
  INVX1 G48404 (.I(W10991), .ZN(O510));
  INVX1 G48405 (.I(W37519), .ZN(O10213));
  INVX1 G48406 (.I(W225), .ZN(W11400));
  INVX1 G48407 (.I(W6635), .ZN(O505));
  INVX1 G48408 (.I(W959), .ZN(O10221));
  INVX1 G48409 (.I(W3500), .ZN(W11403));
  INVX1 G48410 (.I(W10997), .ZN(O10220));
  INVX1 G48411 (.I(W9121), .ZN(W11404));
  INVX1 G48412 (.I(W8603), .ZN(W11407));
  INVX1 G48413 (.I(W39176), .ZN(O10217));
  INVX1 G48414 (.I(W5723), .ZN(O10216));
  INVX1 G48415 (.I(W31784), .ZN(O8639));
  INVX1 G48416 (.I(W365), .ZN(O507));
  INVX1 G48417 (.I(W32277), .ZN(W39439));
  INVX1 G48418 (.I(W1481), .ZN(W11419));
  INVX1 G48419 (.I(W1441), .ZN(W11420));
  INVX1 G48420 (.I(W29721), .ZN(O10203));
  INVX1 G48421 (.I(I424), .ZN(O10202));
  INVX1 G48422 (.I(W10703), .ZN(W11426));
  INVX1 G48423 (.I(W25779), .ZN(W39431));
  INVX1 G48424 (.I(W12514), .ZN(O10201));
  INVX1 G48425 (.I(W15014), .ZN(O7145));
  INVX1 G48426 (.I(I1695), .ZN(O7155));
  INVX1 G48427 (.I(W7274), .ZN(W16635));
  INVX1 G48428 (.I(W573), .ZN(W16639));
  INVX1 G48429 (.I(W32220), .ZN(W34251));
  INVX1 G48430 (.I(W32015), .ZN(O7152));
  INVX1 G48431 (.I(I1978), .ZN(W16641));
  INVX1 G48432 (.I(W312), .ZN(W16643));
  INVX1 G48433 (.I(W9184), .ZN(W16644));
  INVX1 G48434 (.I(W4005), .ZN(O7147));
  INVX1 G48435 (.I(W22141), .ZN(O7146));
  INVX1 G48436 (.I(W905), .ZN(W16633));
  INVX1 G48437 (.I(W3613), .ZN(O7144));
  INVX1 G48438 (.I(W15925), .ZN(O7143));
  INVX1 G48439 (.I(W15723), .ZN(W16647));
  INVX1 G48440 (.I(W316), .ZN(W16650));
  INVX1 G48441 (.I(W5352), .ZN(O1221));
  INVX1 G48442 (.I(I1782), .ZN(W16653));
  INVX1 G48443 (.I(W25689), .ZN(O7142));
  INVX1 G48444 (.I(W15709), .ZN(O1222));
  INVX1 G48445 (.I(W31014), .ZN(O7140));
  INVX1 G48446 (.I(W29971), .ZN(O7159));
  INVX1 G48447 (.I(W20851), .ZN(O7170));
  INVX1 G48448 (.I(W3877), .ZN(O7169));
  INVX1 G48449 (.I(W9558), .ZN(O7168));
  INVX1 G48450 (.I(W27033), .ZN(O7167));
  INVX1 G48451 (.I(W24854), .ZN(O7166));
  INVX1 G48452 (.I(W8433), .ZN(W16606));
  INVX1 G48453 (.I(W7788), .ZN(O7164));
  INVX1 G48454 (.I(I1993), .ZN(W16612));
  INVX1 G48455 (.I(W10951), .ZN(W16613));
  INVX1 G48456 (.I(W9986), .ZN(W16662));
  INVX1 G48457 (.I(W29389), .ZN(W34269));
  INVX1 G48458 (.I(W6746), .ZN(W16620));
  INVX1 G48459 (.I(W23987), .ZN(W34267));
  INVX1 G48460 (.I(W4861), .ZN(O1216));
  INVX1 G48461 (.I(I680), .ZN(W16626));
  INVX1 G48462 (.I(W28700), .ZN(O7156));
  INVX1 G48463 (.I(W11856), .ZN(W16629));
  INVX1 G48464 (.I(I1639), .ZN(W34259));
  INVX1 G48465 (.I(W6687), .ZN(O1217));
  INVX1 G48466 (.I(W19383), .ZN(W34189));
  INVX1 G48467 (.I(W3320), .ZN(O7121));
  INVX1 G48468 (.I(W17288), .ZN(W34202));
  INVX1 G48469 (.I(W20788), .ZN(O7120));
  INVX1 G48470 (.I(W2728), .ZN(O7119));
  INVX1 G48471 (.I(W14472), .ZN(W16694));
  INVX1 G48472 (.I(W19210), .ZN(W34197));
  INVX1 G48473 (.I(W31492), .ZN(W34196));
  INVX1 G48474 (.I(W16046), .ZN(W16697));
  INVX1 G48475 (.I(W12216), .ZN(O1232));
  INVX1 G48476 (.I(W16556), .ZN(O1230));
  INVX1 G48477 (.I(W8792), .ZN(O7115));
  INVX1 G48478 (.I(W14430), .ZN(W16706));
  INVX1 G48479 (.I(W6435), .ZN(O1233));
  INVX1 G48480 (.I(W17221), .ZN(O7110));
  INVX1 G48481 (.I(W19618), .ZN(W34178));
  INVX1 G48482 (.I(W1243), .ZN(W16717));
  INVX1 G48483 (.I(W13341), .ZN(W16718));
  INVX1 G48484 (.I(W6785), .ZN(O7108));
  INVX1 G48485 (.I(W8999), .ZN(O1237));
  INVX1 G48486 (.I(W13050), .ZN(W16677));
  INVX1 G48487 (.I(W646), .ZN(W16663));
  INVX1 G48488 (.I(W14278), .ZN(W16664));
  INVX1 G48489 (.I(W6345), .ZN(W16667));
  INVX1 G48490 (.I(W1762), .ZN(W34227));
  INVX1 G48491 (.I(W111), .ZN(W16672));
  INVX1 G48492 (.I(W7089), .ZN(O7134));
  INVX1 G48493 (.I(W15180), .ZN(W16673));
  INVX1 G48494 (.I(W15550), .ZN(W16675));
  INVX1 G48495 (.I(W9304), .ZN(W34220));
  INVX1 G48496 (.I(W33936), .ZN(W34286));
  INVX1 G48497 (.I(W4337), .ZN(O7129));
  INVX1 G48498 (.I(W8895), .ZN(W16683));
  INVX1 G48499 (.I(W20908), .ZN(W34213));
  INVX1 G48500 (.I(W12126), .ZN(W16685));
  INVX1 G48501 (.I(W1946), .ZN(W16686));
  INVX1 G48502 (.I(W1340), .ZN(O7125));
  INVX1 G48503 (.I(W31512), .ZN(O7124));
  INVX1 G48504 (.I(W14760), .ZN(O7123));
  INVX1 G48505 (.I(W8356), .ZN(O1228));
  INVX1 G48506 (.I(W13861), .ZN(W16513));
  INVX1 G48507 (.I(W5483), .ZN(W34383));
  INVX1 G48508 (.I(W699), .ZN(O7222));
  INVX1 G48509 (.I(W8625), .ZN(W16501));
  INVX1 G48510 (.I(I1156), .ZN(W34377));
  INVX1 G48511 (.I(I843), .ZN(O1187));
  INVX1 G48512 (.I(W5246), .ZN(W16505));
  INVX1 G48513 (.I(W14922), .ZN(W16506));
  INVX1 G48514 (.I(W11716), .ZN(W34373));
  INVX1 G48515 (.I(W29221), .ZN(W34370));
  INVX1 G48516 (.I(W15245), .ZN(O7216));
  INVX1 G48517 (.I(W31007), .ZN(O7223));
  INVX1 G48518 (.I(W4469), .ZN(W16515));
  INVX1 G48519 (.I(W25648), .ZN(O7214));
  INVX1 G48520 (.I(W3209), .ZN(O1190));
  INVX1 G48521 (.I(W2225), .ZN(W34361));
  INVX1 G48522 (.I(W373), .ZN(W34360));
  INVX1 G48523 (.I(W10696), .ZN(W16522));
  INVX1 G48524 (.I(W6464), .ZN(W16527));
  INVX1 G48525 (.I(W11811), .ZN(W16529));
  INVX1 G48526 (.I(I1634), .ZN(W34353));
  INVX1 G48527 (.I(W9002), .ZN(W16477));
  INVX1 G48528 (.I(W26832), .ZN(O7249));
  INVX1 G48529 (.I(W5677), .ZN(W16447));
  INVX1 G48530 (.I(W13000), .ZN(W34416));
  INVX1 G48531 (.I(W28929), .ZN(O7243));
  INVX1 G48532 (.I(W1868), .ZN(O7242));
  INVX1 G48533 (.I(W16157), .ZN(W16459));
  INVX1 G48534 (.I(W8559), .ZN(O1181));
  INVX1 G48535 (.I(W1476), .ZN(W16467));
  INVX1 G48536 (.I(W2662), .ZN(W16471));
  INVX1 G48537 (.I(W8840), .ZN(O1193));
  INVX1 G48538 (.I(I1454), .ZN(W16478));
  INVX1 G48539 (.I(W15230), .ZN(W16481));
  INVX1 G48540 (.I(W17673), .ZN(O7230));
  INVX1 G48541 (.I(I81), .ZN(O1184));
  INVX1 G48542 (.I(W745), .ZN(W16486));
  INVX1 G48543 (.I(W7890), .ZN(O1185));
  INVX1 G48544 (.I(I315), .ZN(W16492));
  INVX1 G48545 (.I(W7693), .ZN(W16493));
  INVX1 G48546 (.I(W14843), .ZN(O7224));
  INVX1 G48547 (.I(W3597), .ZN(W16591));
  INVX1 G48548 (.I(W4272), .ZN(W16576));
  INVX1 G48549 (.I(W10754), .ZN(O7190));
  INVX1 G48550 (.I(W8568), .ZN(W16577));
  INVX1 G48551 (.I(W15714), .ZN(W16578));
  INVX1 G48552 (.I(W8748), .ZN(O7187));
  INVX1 G48553 (.I(W1968), .ZN(W34310));
  INVX1 G48554 (.I(W7665), .ZN(W16585));
  INVX1 G48555 (.I(W31472), .ZN(W34305));
  INVX1 G48556 (.I(W7941), .ZN(W34304));
  INVX1 G48557 (.I(W6974), .ZN(W16575));
  INVX1 G48558 (.I(W27244), .ZN(O7182));
  INVX1 G48559 (.I(W30121), .ZN(W34298));
  INVX1 G48560 (.I(W28266), .ZN(O7178));
  INVX1 G48561 (.I(W21161), .ZN(O7177));
  INVX1 G48562 (.I(W7714), .ZN(W16598));
  INVX1 G48563 (.I(I378), .ZN(O1212));
  INVX1 G48564 (.I(W7140), .ZN(W16601));
  INVX1 G48565 (.I(W12828), .ZN(W16605));
  INVX1 G48566 (.I(W6576), .ZN(O7171));
  INVX1 G48567 (.I(W6415), .ZN(W16558));
  INVX1 G48568 (.I(W29783), .ZN(O7206));
  INVX1 G48569 (.I(W11398), .ZN(W16538));
  INVX1 G48570 (.I(W6026), .ZN(W16540));
  INVX1 G48571 (.I(W2498), .ZN(O7203));
  INVX1 G48572 (.I(W10213), .ZN(W16546));
  INVX1 G48573 (.I(W15368), .ZN(O1198));
  INVX1 G48574 (.I(W1451), .ZN(O1199));
  INVX1 G48575 (.I(W284), .ZN(W16550));
  INVX1 G48576 (.I(W2364), .ZN(O1201));
  INVX1 G48577 (.I(W10616), .ZN(O1238));
  INVX1 G48578 (.I(W20510), .ZN(W34331));
  INVX1 G48579 (.I(W2265), .ZN(O1204));
  INVX1 G48580 (.I(W6144), .ZN(O1205));
  INVX1 G48581 (.I(W24801), .ZN(O7196));
  INVX1 G48582 (.I(W3503), .ZN(W16566));
  INVX1 G48583 (.I(W12433), .ZN(W34325));
  INVX1 G48584 (.I(W5520), .ZN(W16567));
  INVX1 G48585 (.I(W30310), .ZN(O7194));
  INVX1 G48586 (.I(W12242), .ZN(W16572));
  INVX1 G48587 (.I(W15895), .ZN(W16898));
  INVX1 G48588 (.I(W7052), .ZN(W34018));
  INVX1 G48589 (.I(W467), .ZN(O7015));
  INVX1 G48590 (.I(W123), .ZN(O7014));
  INVX1 G48591 (.I(W4321), .ZN(W16881));
  INVX1 G48592 (.I(W4025), .ZN(W16886));
  INVX1 G48593 (.I(W3987), .ZN(W34012));
  INVX1 G48594 (.I(W6198), .ZN(O7012));
  INVX1 G48595 (.I(W6322), .ZN(W16892));
  INVX1 G48596 (.I(W17698), .ZN(W34005));
  INVX1 G48597 (.I(W24999), .ZN(W34003));
  INVX1 G48598 (.I(W23897), .ZN(O7016));
  INVX1 G48599 (.I(W20646), .ZN(O7005));
  INVX1 G48600 (.I(W16144), .ZN(O1278));
  INVX1 G48601 (.I(W10282), .ZN(W16905));
  INVX1 G48602 (.I(W33755), .ZN(O7002));
  INVX1 G48603 (.I(W9459), .ZN(W16907));
  INVX1 G48604 (.I(I508), .ZN(W16910));
  INVX1 G48605 (.I(W18604), .ZN(W33991));
  INVX1 G48606 (.I(W15037), .ZN(O7000));
  INVX1 G48607 (.I(W28547), .ZN(W33989));
  INVX1 G48608 (.I(W30872), .ZN(O7027));
  INVX1 G48609 (.I(W24413), .ZN(O7037));
  INVX1 G48610 (.I(W13083), .ZN(W16845));
  INVX1 G48611 (.I(W23985), .ZN(W34049));
  INVX1 G48612 (.I(W7875), .ZN(W16852));
  INVX1 G48613 (.I(W26840), .ZN(O7032));
  INVX1 G48614 (.I(W16640), .ZN(O1273));
  INVX1 G48615 (.I(W5558), .ZN(O7029));
  INVX1 G48616 (.I(W8171), .ZN(W16864));
  INVX1 G48617 (.I(W828), .ZN(W16866));
  INVX1 G48618 (.I(W5331), .ZN(W16912));
  INVX1 G48619 (.I(W2037), .ZN(W16869));
  INVX1 G48620 (.I(W12162), .ZN(W16870));
  INVX1 G48621 (.I(W2661), .ZN(W16872));
  INVX1 G48622 (.I(W12194), .ZN(W16873));
  INVX1 G48623 (.I(W31258), .ZN(O7024));
  INVX1 G48624 (.I(W32528), .ZN(O7023));
  INVX1 G48625 (.I(W12986), .ZN(O7021));
  INVX1 G48626 (.I(W29246), .ZN(O7019));
  INVX1 G48627 (.I(W24081), .ZN(O7017));
  INVX1 G48628 (.I(W30939), .ZN(O6968));
  INVX1 G48629 (.I(W13395), .ZN(W16952));
  INVX1 G48630 (.I(W28853), .ZN(O6974));
  INVX1 G48631 (.I(W10393), .ZN(W16954));
  INVX1 G48632 (.I(W23017), .ZN(W33949));
  INVX1 G48633 (.I(W14678), .ZN(W16957));
  INVX1 G48634 (.I(W13477), .ZN(W16959));
  INVX1 G48635 (.I(W5115), .ZN(W16960));
  INVX1 G48636 (.I(W5379), .ZN(W16962));
  INVX1 G48637 (.I(W9312), .ZN(W16964));
  INVX1 G48638 (.I(W9169), .ZN(W16948));
  INVX1 G48639 (.I(W7541), .ZN(O6967));
  INVX1 G48640 (.I(W5650), .ZN(O1289));
  INVX1 G48641 (.I(W16452), .ZN(W33937));
  INVX1 G48642 (.I(W10549), .ZN(W16970));
  INVX1 G48643 (.I(W2950), .ZN(W16974));
  INVX1 G48644 (.I(W15078), .ZN(W33931));
  INVX1 G48645 (.I(W3615), .ZN(W33929));
  INVX1 G48646 (.I(W10346), .ZN(O1292));
  INVX1 G48647 (.I(W26253), .ZN(W33927));
  INVX1 G48648 (.I(W7427), .ZN(W33970));
  INVX1 G48649 (.I(W27431), .ZN(O6999));
  INVX1 G48650 (.I(W2394), .ZN(W16913));
  INVX1 G48651 (.I(W698), .ZN(W16917));
  INVX1 G48652 (.I(W3800), .ZN(W16922));
  INVX1 G48653 (.I(W10205), .ZN(O6992));
  INVX1 G48654 (.I(W9952), .ZN(O6990));
  INVX1 G48655 (.I(W3386), .ZN(O6986));
  INVX1 G48656 (.I(W19610), .ZN(W33972));
  INVX1 G48657 (.I(I1895), .ZN(W33971));
  INVX1 G48658 (.I(W5330), .ZN(W34057));
  INVX1 G48659 (.I(W2234), .ZN(W33968));
  INVX1 G48660 (.I(W654), .ZN(O1286));
  INVX1 G48661 (.I(I906), .ZN(O6984));
  INVX1 G48662 (.I(W7036), .ZN(O6983));
  INVX1 G48663 (.I(W7912), .ZN(O6982));
  INVX1 G48664 (.I(W4930), .ZN(W16939));
  INVX1 G48665 (.I(W15670), .ZN(W16942));
  INVX1 G48666 (.I(W5341), .ZN(W16943));
  INVX1 G48667 (.I(W26439), .ZN(O6979));
  INVX1 G48668 (.I(W7952), .ZN(O7083));
  INVX1 G48669 (.I(W9403), .ZN(W16741));
  INVX1 G48670 (.I(W17377), .ZN(W34145));
  INVX1 G48671 (.I(W15318), .ZN(O1247));
  INVX1 G48672 (.I(W8712), .ZN(W34140));
  INVX1 G48673 (.I(W11993), .ZN(O7086));
  INVX1 G48674 (.I(W25290), .ZN(O7085));
  INVX1 G48675 (.I(W5640), .ZN(O1251));
  INVX1 G48676 (.I(W8195), .ZN(W16753));
  INVX1 G48677 (.I(W4863), .ZN(W34132));
  INVX1 G48678 (.I(W27023), .ZN(O7090));
  INVX1 G48679 (.I(W5740), .ZN(O1253));
  INVX1 G48680 (.I(W6737), .ZN(O1254));
  INVX1 G48681 (.I(W18841), .ZN(O7079));
  INVX1 G48682 (.I(W10822), .ZN(W16771));
  INVX1 G48683 (.I(W23488), .ZN(W34121));
  INVX1 G48684 (.I(W7003), .ZN(W16774));
  INVX1 G48685 (.I(W14374), .ZN(W16777));
  INVX1 G48686 (.I(W6750), .ZN(O1258));
  INVX1 G48687 (.I(W7289), .ZN(W34115));
  INVX1 G48688 (.I(W19136), .ZN(W34158));
  INVX1 G48689 (.I(W10811), .ZN(W16723));
  INVX1 G48690 (.I(W11285), .ZN(W16725));
  INVX1 G48691 (.I(W28996), .ZN(O7103));
  INVX1 G48692 (.I(W7579), .ZN(W16726));
  INVX1 G48693 (.I(W1778), .ZN(W16727));
  INVX1 G48694 (.I(W4117), .ZN(W16731));
  INVX1 G48695 (.I(W2792), .ZN(O7101));
  INVX1 G48696 (.I(W17820), .ZN(O7100));
  INVX1 G48697 (.I(W4528), .ZN(O7097));
  INVX1 G48698 (.I(W8532), .ZN(O1259));
  INVX1 G48699 (.I(W27479), .ZN(W34157));
  INVX1 G48700 (.I(W1841), .ZN(W16736));
  INVX1 G48701 (.I(W8375), .ZN(O7095));
  INVX1 G48702 (.I(W30215), .ZN(W34153));
  INVX1 G48703 (.I(W5753), .ZN(W16738));
  INVX1 G48704 (.I(W16461), .ZN(O7092));
  INVX1 G48705 (.I(W25639), .ZN(W34150));
  INVX1 G48706 (.I(I836), .ZN(W34149));
  INVX1 G48707 (.I(W8648), .ZN(O1245));
  INVX1 G48708 (.I(W2897), .ZN(W16825));
  INVX1 G48709 (.I(W14031), .ZN(W16812));
  INVX1 G48710 (.I(I488), .ZN(W16815));
  INVX1 G48711 (.I(W8987), .ZN(W16817));
  INVX1 G48712 (.I(W15831), .ZN(W16818));
  INVX1 G48713 (.I(I958), .ZN(W34078));
  INVX1 G48714 (.I(W9535), .ZN(O7056));
  INVX1 G48715 (.I(W16509), .ZN(W16820));
  INVX1 G48716 (.I(W20320), .ZN(W34073));
  INVX1 G48717 (.I(W4865), .ZN(W16823));
  INVX1 G48718 (.I(W2959), .ZN(O1268));
  INVX1 G48719 (.I(W18604), .ZN(O7049));
  INVX1 G48720 (.I(W30294), .ZN(O7048));
  INVX1 G48721 (.I(W14817), .ZN(O1270));
  INVX1 G48722 (.I(W1184), .ZN(W16829));
  INVX1 G48723 (.I(W6139), .ZN(O1271));
  INVX1 G48724 (.I(W15747), .ZN(W16834));
  INVX1 G48725 (.I(W24753), .ZN(O7043));
  INVX1 G48726 (.I(W26193), .ZN(W34059));
  INVX1 G48727 (.I(W11771), .ZN(O7041));
  INVX1 G48728 (.I(W8674), .ZN(O1263));
  INVX1 G48729 (.I(W8642), .ZN(O7073));
  INVX1 G48730 (.I(W13164), .ZN(W16781));
  INVX1 G48731 (.I(I52), .ZN(W16785));
  INVX1 G48732 (.I(W11365), .ZN(O1261));
  INVX1 G48733 (.I(W14543), .ZN(O7069));
  INVX1 G48734 (.I(W5686), .ZN(W34105));
  INVX1 G48735 (.I(W27772), .ZN(W34104));
  INVX1 G48736 (.I(W4096), .ZN(W16794));
  INVX1 G48737 (.I(W7310), .ZN(O7066));
  INVX1 G48738 (.I(W5858), .ZN(O7250));
  INVX1 G48739 (.I(W4168), .ZN(W16796));
  INVX1 G48740 (.I(W4139), .ZN(W16798));
  INVX1 G48741 (.I(W2993), .ZN(O1266));
  INVX1 G48742 (.I(W7869), .ZN(W16804));
  INVX1 G48743 (.I(W11254), .ZN(W34093));
  INVX1 G48744 (.I(W17529), .ZN(W34091));
  INVX1 G48745 (.I(W33865), .ZN(W34089));
  INVX1 G48746 (.I(W12673), .ZN(W16808));
  INVX1 G48747 (.I(W14187), .ZN(O7060));
  INVX1 G48748 (.I(W9095), .ZN(W16082));
  INVX1 G48749 (.I(W481), .ZN(W16072));
  INVX1 G48750 (.I(I448), .ZN(O7426));
  INVX1 G48751 (.I(W15182), .ZN(W34747));
  INVX1 G48752 (.I(W20928), .ZN(W34746));
  INVX1 G48753 (.I(W15362), .ZN(W34745));
  INVX1 G48754 (.I(W9494), .ZN(W16074));
  INVX1 G48755 (.I(W12133), .ZN(O7423));
  INVX1 G48756 (.I(W4470), .ZN(W16081));
  INVX1 G48757 (.I(W16442), .ZN(O7421));
  INVX1 G48758 (.I(W23043), .ZN(O7420));
  INVX1 G48759 (.I(W12294), .ZN(W16071));
  INVX1 G48760 (.I(W33817), .ZN(W34736));
  INVX1 G48761 (.I(W14956), .ZN(W16087));
  INVX1 G48762 (.I(W9029), .ZN(W16091));
  INVX1 G48763 (.I(W30496), .ZN(W34730));
  INVX1 G48764 (.I(W9899), .ZN(O1119));
  INVX1 G48765 (.I(W25236), .ZN(W34728));
  INVX1 G48766 (.I(W7905), .ZN(W16093));
  INVX1 G48767 (.I(W9150), .ZN(W34725));
  INVX1 G48768 (.I(W22230), .ZN(O7412));
  INVX1 G48769 (.I(W9743), .ZN(W16062));
  INVX1 G48770 (.I(W3477), .ZN(W34775));
  INVX1 G48771 (.I(W21527), .ZN(O7441));
  INVX1 G48772 (.I(W8865), .ZN(W16047));
  INVX1 G48773 (.I(W3230), .ZN(W16051));
  INVX1 G48774 (.I(W6688), .ZN(W16054));
  INVX1 G48775 (.I(W5627), .ZN(W34766));
  INVX1 G48776 (.I(W4999), .ZN(W34765));
  INVX1 G48777 (.I(W89), .ZN(W16058));
  INVX1 G48778 (.I(W14298), .ZN(W16060));
  INVX1 G48779 (.I(W20225), .ZN(W34723));
  INVX1 G48780 (.I(W2336), .ZN(W16063));
  INVX1 G48781 (.I(W9988), .ZN(W16064));
  INVX1 G48782 (.I(W11400), .ZN(W16065));
  INVX1 G48783 (.I(W6460), .ZN(W16068));
  INVX1 G48784 (.I(W26080), .ZN(O7432));
  INVX1 G48785 (.I(W1673), .ZN(O7430));
  INVX1 G48786 (.I(W5234), .ZN(W34753));
  INVX1 G48787 (.I(W953), .ZN(O1116));
  INVX1 G48788 (.I(W12997), .ZN(O7429));
  INVX1 G48789 (.I(W889), .ZN(W16132));
  INVX1 G48790 (.I(W9760), .ZN(W34697));
  INVX1 G48791 (.I(I748), .ZN(W16123));
  INVX1 G48792 (.I(W14830), .ZN(O7396));
  INVX1 G48793 (.I(W1865), .ZN(W16126));
  INVX1 G48794 (.I(W6820), .ZN(W16127));
  INVX1 G48795 (.I(W6671), .ZN(W16128));
  INVX1 G48796 (.I(W33927), .ZN(O7395));
  INVX1 G48797 (.I(W14225), .ZN(W34690));
  INVX1 G48798 (.I(I970), .ZN(W16129));
  INVX1 G48799 (.I(W17713), .ZN(O7397));
  INVX1 G48800 (.I(W20054), .ZN(W34686));
  INVX1 G48801 (.I(W11756), .ZN(W34685));
  INVX1 G48802 (.I(W20440), .ZN(O7393));
  INVX1 G48803 (.I(W6307), .ZN(W16135));
  INVX1 G48804 (.I(W9499), .ZN(O7391));
  INVX1 G48805 (.I(W14983), .ZN(O7389));
  INVX1 G48806 (.I(W19963), .ZN(O7387));
  INVX1 G48807 (.I(W9762), .ZN(W16148));
  INVX1 G48808 (.I(W22193), .ZN(O7385));
  INVX1 G48809 (.I(W27003), .ZN(O7405));
  INVX1 G48810 (.I(W6793), .ZN(W34722));
  INVX1 G48811 (.I(W4039), .ZN(W34719));
  INVX1 G48812 (.I(W29094), .ZN(O7409));
  INVX1 G48813 (.I(W13938), .ZN(W16101));
  INVX1 G48814 (.I(W3890), .ZN(W16103));
  INVX1 G48815 (.I(W3295), .ZN(O1120));
  INVX1 G48816 (.I(I1970), .ZN(O1121));
  INVX1 G48817 (.I(W25831), .ZN(W34712));
  INVX1 G48818 (.I(W16254), .ZN(W34710));
  INVX1 G48819 (.I(W8232), .ZN(O7442));
  INVX1 G48820 (.I(W33527), .ZN(W34708));
  INVX1 G48821 (.I(W10561), .ZN(W16110));
  INVX1 G48822 (.I(W3947), .ZN(W16114));
  INVX1 G48823 (.I(W22928), .ZN(O7402));
  INVX1 G48824 (.I(W16019), .ZN(W16115));
  INVX1 G48825 (.I(W3210), .ZN(W16118));
  INVX1 G48826 (.I(W550), .ZN(O1125));
  INVX1 G48827 (.I(W6364), .ZN(W16121));
  INVX1 G48828 (.I(W3549), .ZN(W16122));
  INVX1 G48829 (.I(W2277), .ZN(W15980));
  INVX1 G48830 (.I(W5264), .ZN(W34858));
  INVX1 G48831 (.I(W6487), .ZN(W15968));
  INVX1 G48832 (.I(W29150), .ZN(O7481));
  INVX1 G48833 (.I(I3), .ZN(O1097));
  INVX1 G48834 (.I(W9012), .ZN(W15975));
  INVX1 G48835 (.I(W26674), .ZN(O7479));
  INVX1 G48836 (.I(W7598), .ZN(W15978));
  INVX1 G48837 (.I(W22899), .ZN(O7478));
  INVX1 G48838 (.I(W6194), .ZN(W15979));
  INVX1 G48839 (.I(W6017), .ZN(W15964));
  INVX1 G48840 (.I(W8401), .ZN(W15981));
  INVX1 G48841 (.I(W13321), .ZN(W15983));
  INVX1 G48842 (.I(W21998), .ZN(O7474));
  INVX1 G48843 (.I(I1286), .ZN(O7473));
  INVX1 G48844 (.I(W6655), .ZN(W15986));
  INVX1 G48845 (.I(W15066), .ZN(W15987));
  INVX1 G48846 (.I(W4901), .ZN(W15988));
  INVX1 G48847 (.I(W3918), .ZN(W34835));
  INVX1 G48848 (.I(W4508), .ZN(W15991));
  INVX1 G48849 (.I(W15209), .ZN(O7491));
  INVX1 G48850 (.I(W8653), .ZN(W34886));
  INVX1 G48851 (.I(I261), .ZN(W15947));
  INVX1 G48852 (.I(W7155), .ZN(W15948));
  INVX1 G48853 (.I(W13575), .ZN(W15949));
  INVX1 G48854 (.I(W277), .ZN(O7493));
  INVX1 G48855 (.I(W11159), .ZN(W34880));
  INVX1 G48856 (.I(W21066), .ZN(W34877));
  INVX1 G48857 (.I(W12234), .ZN(W15953));
  INVX1 G48858 (.I(W6913), .ZN(W15955));
  INVX1 G48859 (.I(W33395), .ZN(W34831));
  INVX1 G48860 (.I(W17841), .ZN(W34872));
  INVX1 G48861 (.I(W126), .ZN(W34871));
  INVX1 G48862 (.I(W5130), .ZN(W15957));
  INVX1 G48863 (.I(W25466), .ZN(O7489));
  INVX1 G48864 (.I(W3003), .ZN(W15959));
  INVX1 G48865 (.I(W15717), .ZN(W34866));
  INVX1 G48866 (.I(W1779), .ZN(W15960));
  INVX1 G48867 (.I(W12371), .ZN(O7487));
  INVX1 G48868 (.I(W12571), .ZN(W34861));
  INVX1 G48869 (.I(W1790), .ZN(O1110));
  INVX1 G48870 (.I(I1194), .ZN(W34806));
  INVX1 G48871 (.I(I1447), .ZN(O1104));
  INVX1 G48872 (.I(W10435), .ZN(W34803));
  INVX1 G48873 (.I(W4774), .ZN(O7454));
  INVX1 G48874 (.I(W4639), .ZN(W34799));
  INVX1 G48875 (.I(W4476), .ZN(W16029));
  INVX1 G48876 (.I(W3140), .ZN(W34797));
  INVX1 G48877 (.I(W4312), .ZN(W34796));
  INVX1 G48878 (.I(W32491), .ZN(O7452));
  INVX1 G48879 (.I(I1457), .ZN(W16015));
  INVX1 G48880 (.I(W3814), .ZN(W16031));
  INVX1 G48881 (.I(W25749), .ZN(W34792));
  INVX1 G48882 (.I(W5713), .ZN(W34791));
  INVX1 G48883 (.I(W31327), .ZN(O7448));
  INVX1 G48884 (.I(W33053), .ZN(O7447));
  INVX1 G48885 (.I(W1778), .ZN(W34783));
  INVX1 G48886 (.I(W13845), .ZN(W16040));
  INVX1 G48887 (.I(W11941), .ZN(W16041));
  INVX1 G48888 (.I(W8706), .ZN(O7445));
  INVX1 G48889 (.I(W18813), .ZN(O7462));
  INVX1 G48890 (.I(W7088), .ZN(W34829));
  INVX1 G48891 (.I(W554), .ZN(W15996));
  INVX1 G48892 (.I(W3718), .ZN(O7468));
  INVX1 G48893 (.I(W13253), .ZN(W15998));
  INVX1 G48894 (.I(W15791), .ZN(O7465));
  INVX1 G48895 (.I(W13040), .ZN(W16000));
  INVX1 G48896 (.I(W23639), .ZN(W34821));
  INVX1 G48897 (.I(I1506), .ZN(W16001));
  INVX1 G48898 (.I(W3671), .ZN(W16003));
  INVX1 G48899 (.I(W2114), .ZN(W16149));
  INVX1 G48900 (.I(W14624), .ZN(W16006));
  INVX1 G48901 (.I(W837), .ZN(W34815));
  INVX1 G48902 (.I(W26072), .ZN(O7459));
  INVX1 G48903 (.I(W579), .ZN(W16007));
  INVX1 G48904 (.I(W7090), .ZN(O1103));
  INVX1 G48905 (.I(W15089), .ZN(W16010));
  INVX1 G48906 (.I(W13526), .ZN(W16011));
  INVX1 G48907 (.I(W12486), .ZN(W16014));
  INVX1 G48908 (.I(W1767), .ZN(W34808));
  INVX1 G48909 (.I(W18415), .ZN(O7294));
  INVX1 G48910 (.I(W12532), .ZN(O7303));
  INVX1 G48911 (.I(W22814), .ZN(O7300));
  INVX1 G48912 (.I(W6448), .ZN(W16340));
  INVX1 G48913 (.I(W17101), .ZN(O7299));
  INVX1 G48914 (.I(W7465), .ZN(O7297));
  INVX1 G48915 (.I(W5523), .ZN(W16349));
  INVX1 G48916 (.I(W2362), .ZN(W34504));
  INVX1 G48917 (.I(W4828), .ZN(O7295));
  INVX1 G48918 (.I(W32053), .ZN(W34502));
  INVX1 G48919 (.I(W994), .ZN(O1161));
  INVX1 G48920 (.I(W10242), .ZN(W16334));
  INVX1 G48921 (.I(W381), .ZN(O1163));
  INVX1 G48922 (.I(W6169), .ZN(W34496));
  INVX1 G48923 (.I(W9750), .ZN(W16360));
  INVX1 G48924 (.I(W107), .ZN(W16361));
  INVX1 G48925 (.I(W25505), .ZN(O7287));
  INVX1 G48926 (.I(W16349), .ZN(W16369));
  INVX1 G48927 (.I(W8831), .ZN(O1170));
  INVX1 G48928 (.I(W20848), .ZN(W34486));
  INVX1 G48929 (.I(W15408), .ZN(W16373));
  INVX1 G48930 (.I(W14963), .ZN(W34528));
  INVX1 G48931 (.I(W12688), .ZN(O1157));
  INVX1 G48932 (.I(W2828), .ZN(W16313));
  INVX1 G48933 (.I(W31477), .ZN(O7316));
  INVX1 G48934 (.I(W33051), .ZN(O7315));
  INVX1 G48935 (.I(W4609), .ZN(W16315));
  INVX1 G48936 (.I(W11374), .ZN(W16319));
  INVX1 G48937 (.I(W13516), .ZN(W16322));
  INVX1 G48938 (.I(W4982), .ZN(W16325));
  INVX1 G48939 (.I(W17764), .ZN(W34529));
  INVX1 G48940 (.I(W5366), .ZN(O7283));
  INVX1 G48941 (.I(W15504), .ZN(O7311));
  INVX1 G48942 (.I(W14312), .ZN(W16326));
  INVX1 G48943 (.I(I929), .ZN(W16327));
  INVX1 G48944 (.I(W10487), .ZN(W16330));
  INVX1 G48945 (.I(W19071), .ZN(W34522));
  INVX1 G48946 (.I(W611), .ZN(W16332));
  INVX1 G48947 (.I(W13813), .ZN(W16333));
  INVX1 G48948 (.I(W18779), .ZN(W34519));
  INVX1 G48949 (.I(W16612), .ZN(O7306));
  INVX1 G48950 (.I(W5932), .ZN(O1176));
  INVX1 G48951 (.I(W12932), .ZN(W16409));
  INVX1 G48952 (.I(W28923), .ZN(W34453));
  INVX1 G48953 (.I(W33095), .ZN(O7264));
  INVX1 G48954 (.I(W7884), .ZN(W16412));
  INVX1 G48955 (.I(W1656), .ZN(W16414));
  INVX1 G48956 (.I(W12544), .ZN(O1174));
  INVX1 G48957 (.I(W12027), .ZN(W16421));
  INVX1 G48958 (.I(W1188), .ZN(W34444));
  INVX1 G48959 (.I(W6662), .ZN(W16423));
  INVX1 G48960 (.I(W7205), .ZN(W16407));
  INVX1 G48961 (.I(W12164), .ZN(O1177));
  INVX1 G48962 (.I(W30215), .ZN(O7258));
  INVX1 G48963 (.I(W14931), .ZN(W16430));
  INVX1 G48964 (.I(W6447), .ZN(W16431));
  INVX1 G48965 (.I(I1020), .ZN(W34435));
  INVX1 G48966 (.I(W31801), .ZN(O7255));
  INVX1 G48967 (.I(W7178), .ZN(W34431));
  INVX1 G48968 (.I(W19563), .ZN(W34428));
  INVX1 G48969 (.I(W31139), .ZN(O7251));
  INVX1 G48970 (.I(W32215), .ZN(O7275));
  INVX1 G48971 (.I(W11124), .ZN(W16376));
  INVX1 G48972 (.I(W27455), .ZN(W34480));
  INVX1 G48973 (.I(W348), .ZN(W16377));
  INVX1 G48974 (.I(W5116), .ZN(W16378));
  INVX1 G48975 (.I(W9721), .ZN(W34475));
  INVX1 G48976 (.I(W24355), .ZN(O7279));
  INVX1 G48977 (.I(W2671), .ZN(W16382));
  INVX1 G48978 (.I(W2501), .ZN(W16386));
  INVX1 G48979 (.I(I56), .ZN(O7276));
  INVX1 G48980 (.I(W3315), .ZN(W16307));
  INVX1 G48981 (.I(W14928), .ZN(W16391));
  INVX1 G48982 (.I(W502), .ZN(O1172));
  INVX1 G48983 (.I(W10117), .ZN(W16393));
  INVX1 G48984 (.I(W14433), .ZN(W16397));
  INVX1 G48985 (.I(W10206), .ZN(W16398));
  INVX1 G48986 (.I(W12435), .ZN(W16400));
  INVX1 G48987 (.I(W10153), .ZN(W16402));
  INVX1 G48988 (.I(W3720), .ZN(W16406));
  INVX1 G48989 (.I(W22197), .ZN(O7267));
  INVX1 G48990 (.I(W8377), .ZN(W16228));
  INVX1 G48991 (.I(W6551), .ZN(W16200));
  INVX1 G48992 (.I(W3801), .ZN(O7367));
  INVX1 G48993 (.I(W5022), .ZN(W16202));
  INVX1 G48994 (.I(W20375), .ZN(O7365));
  INVX1 G48995 (.I(W1283), .ZN(W16206));
  INVX1 G48996 (.I(W8448), .ZN(W16208));
  INVX1 G48997 (.I(W13833), .ZN(W16213));
  INVX1 G48998 (.I(W27051), .ZN(O7358));
  INVX1 G48999 (.I(W22800), .ZN(W34615));
  INVX1 G49000 (.I(W712), .ZN(W34636));
  INVX1 G49001 (.I(W1133), .ZN(W16229));
  INVX1 G49002 (.I(W11323), .ZN(W16230));
  INVX1 G49003 (.I(W20850), .ZN(W34610));
  INVX1 G49004 (.I(W27091), .ZN(O7353));
  INVX1 G49005 (.I(W19766), .ZN(O7352));
  INVX1 G49006 (.I(W9742), .ZN(W16234));
  INVX1 G49007 (.I(W26468), .ZN(O7349));
  INVX1 G49008 (.I(W951), .ZN(W34604));
  INVX1 G49009 (.I(W13802), .ZN(W34603));
  INVX1 G49010 (.I(W16059), .ZN(W16186));
  INVX1 G49011 (.I(W2669), .ZN(O1132));
  INVX1 G49012 (.I(W8466), .ZN(O7381));
  INVX1 G49013 (.I(W2318), .ZN(O7379));
  INVX1 G49014 (.I(W6667), .ZN(W16165));
  INVX1 G49015 (.I(W7800), .ZN(W34659));
  INVX1 G49016 (.I(W10801), .ZN(W16176));
  INVX1 G49017 (.I(I916), .ZN(O7374));
  INVX1 G49018 (.I(I1006), .ZN(O1136));
  INVX1 G49019 (.I(W15118), .ZN(W16184));
  INVX1 G49020 (.I(W6331), .ZN(W16236));
  INVX1 G49021 (.I(W9568), .ZN(W16190));
  INVX1 G49022 (.I(W13142), .ZN(W16191));
  INVX1 G49023 (.I(W15846), .ZN(W16192));
  INVX1 G49024 (.I(W13795), .ZN(W16193));
  INVX1 G49025 (.I(W24991), .ZN(W34643));
  INVX1 G49026 (.I(W6619), .ZN(W16194));
  INVX1 G49027 (.I(W4386), .ZN(W34641));
  INVX1 G49028 (.I(W2297), .ZN(W34639));
  INVX1 G49029 (.I(W30487), .ZN(W34638));
  INVX1 G49030 (.I(W13879), .ZN(W16290));
  INVX1 G49031 (.I(W1707), .ZN(W16276));
  INVX1 G49032 (.I(W9595), .ZN(W16280));
  INVX1 G49033 (.I(W6704), .ZN(W16281));
  INVX1 G49034 (.I(W2917), .ZN(W16282));
  INVX1 G49035 (.I(W26216), .ZN(O7329));
  INVX1 G49036 (.I(W8768), .ZN(O1154));
  INVX1 G49037 (.I(W12734), .ZN(W16286));
  INVX1 G49038 (.I(W10291), .ZN(W16287));
  INVX1 G49039 (.I(I1970), .ZN(W16289));
  INVX1 G49040 (.I(W7343), .ZN(O1152));
  INVX1 G49041 (.I(W32534), .ZN(O7327));
  INVX1 G49042 (.I(W4224), .ZN(O7325));
  INVX1 G49043 (.I(W7114), .ZN(W16293));
  INVX1 G49044 (.I(I1243), .ZN(W16294));
  INVX1 G49045 (.I(W10205), .ZN(O7323));
  INVX1 G49046 (.I(W22162), .ZN(W34548));
  INVX1 G49047 (.I(W11374), .ZN(O7321));
  INVX1 G49048 (.I(W9017), .ZN(W16300));
  INVX1 G49049 (.I(W12931), .ZN(W16306));
  INVX1 G49050 (.I(W20439), .ZN(O7340));
  INVX1 G49051 (.I(W17960), .ZN(O7347));
  INVX1 G49052 (.I(I1590), .ZN(W16244));
  INVX1 G49053 (.I(W15698), .ZN(W34597));
  INVX1 G49054 (.I(W16046), .ZN(W16250));
  INVX1 G49055 (.I(W9814), .ZN(W16251));
  INVX1 G49056 (.I(W9033), .ZN(O1146));
  INVX1 G49057 (.I(W2235), .ZN(W16256));
  INVX1 G49058 (.I(W15077), .ZN(O1147));
  INVX1 G49059 (.I(W6176), .ZN(O7341));
  INVX1 G49060 (.I(W8799), .ZN(O1294));
  INVX1 G49061 (.I(W12314), .ZN(W16263));
  INVX1 G49062 (.I(W6737), .ZN(W16264));
  INVX1 G49063 (.I(W29012), .ZN(O7337));
  INVX1 G49064 (.I(W9007), .ZN(W16265));
  INVX1 G49065 (.I(W30682), .ZN(W34579));
  INVX1 G49066 (.I(W11210), .ZN(W16266));
  INVX1 G49067 (.I(W14618), .ZN(W16269));
  INVX1 G49068 (.I(W22215), .ZN(O7334));
  INVX1 G49069 (.I(W12658), .ZN(W16270));
  INVX1 G49070 (.I(W4903), .ZN(W17627));
  INVX1 G49071 (.I(W17596), .ZN(W33284));
  INVX1 G49072 (.I(W13228), .ZN(W17603));
  INVX1 G49073 (.I(W269), .ZN(O1416));
  INVX1 G49074 (.I(W16876), .ZN(W33279));
  INVX1 G49075 (.I(I297), .ZN(W17608));
  INVX1 G49076 (.I(W8905), .ZN(W17616));
  INVX1 G49077 (.I(W11763), .ZN(W17618));
  INVX1 G49078 (.I(W4657), .ZN(W17623));
  INVX1 G49079 (.I(W16940), .ZN(O1417));
  INVX1 G49080 (.I(W29943), .ZN(O6628));
  INVX1 G49081 (.I(W10964), .ZN(O1415));
  INVX1 G49082 (.I(W17047), .ZN(W33266));
  INVX1 G49083 (.I(W11836), .ZN(O1418));
  INVX1 G49084 (.I(W2205), .ZN(W17630));
  INVX1 G49085 (.I(W5850), .ZN(W17633));
  INVX1 G49086 (.I(I896), .ZN(W17635));
  INVX1 G49087 (.I(W10756), .ZN(O6624));
  INVX1 G49088 (.I(W16972), .ZN(W33257));
  INVX1 G49089 (.I(W15899), .ZN(O1419));
  INVX1 G49090 (.I(W15209), .ZN(W17639));
  INVX1 G49091 (.I(W987), .ZN(W17588));
  INVX1 G49092 (.I(W4682), .ZN(O6645));
  INVX1 G49093 (.I(W13614), .ZN(W33319));
  INVX1 G49094 (.I(W7836), .ZN(O6644));
  INVX1 G49095 (.I(I1577), .ZN(W33315));
  INVX1 G49096 (.I(I1913), .ZN(W17567));
  INVX1 G49097 (.I(W12156), .ZN(W17574));
  INVX1 G49098 (.I(W15819), .ZN(W17576));
  INVX1 G49099 (.I(W5750), .ZN(W33304));
  INVX1 G49100 (.I(W3673), .ZN(W17586));
  INVX1 G49101 (.I(W21873), .ZN(W33253));
  INVX1 G49102 (.I(W33262), .ZN(W33298));
  INVX1 G49103 (.I(W8478), .ZN(W17591));
  INVX1 G49104 (.I(W17564), .ZN(W17592));
  INVX1 G49105 (.I(W9855), .ZN(O6636));
  INVX1 G49106 (.I(W3351), .ZN(O6635));
  INVX1 G49107 (.I(W4513), .ZN(W17594));
  INVX1 G49108 (.I(W16817), .ZN(W17597));
  INVX1 G49109 (.I(I1416), .ZN(O1412));
  INVX1 G49110 (.I(I1221), .ZN(O1413));
  INVX1 G49111 (.I(W8491), .ZN(W17666));
  INVX1 G49112 (.I(W8177), .ZN(W17655));
  INVX1 G49113 (.I(W22097), .ZN(W33227));
  INVX1 G49114 (.I(W17562), .ZN(O1424));
  INVX1 G49115 (.I(W23783), .ZN(W33225));
  INVX1 G49116 (.I(W7790), .ZN(W17660));
  INVX1 G49117 (.I(I1366), .ZN(O6603));
  INVX1 G49118 (.I(W12320), .ZN(O6601));
  INVX1 G49119 (.I(W7769), .ZN(W17664));
  INVX1 G49120 (.I(W28177), .ZN(O6599));
  INVX1 G49121 (.I(W8390), .ZN(W17652));
  INVX1 G49122 (.I(W7238), .ZN(W33215));
  INVX1 G49123 (.I(W4613), .ZN(O1426));
  INVX1 G49124 (.I(W12418), .ZN(W17669));
  INVX1 G49125 (.I(W12778), .ZN(O6595));
  INVX1 G49126 (.I(W20179), .ZN(O6594));
  INVX1 G49127 (.I(W21144), .ZN(W33206));
  INVX1 G49128 (.I(W9166), .ZN(W17673));
  INVX1 G49129 (.I(W28284), .ZN(O6593));
  INVX1 G49130 (.I(W28088), .ZN(W33203));
  INVX1 G49131 (.I(W7833), .ZN(W17644));
  INVX1 G49132 (.I(W9459), .ZN(O1420));
  INVX1 G49133 (.I(W31545), .ZN(O6620));
  INVX1 G49134 (.I(W11916), .ZN(O6619));
  INVX1 G49135 (.I(W21184), .ZN(O6618));
  INVX1 G49136 (.I(W5559), .ZN(O6617));
  INVX1 G49137 (.I(W14770), .ZN(W33246));
  INVX1 G49138 (.I(W25015), .ZN(O6616));
  INVX1 G49139 (.I(W29575), .ZN(W33244));
  INVX1 G49140 (.I(W2186), .ZN(O6615));
  INVX1 G49141 (.I(W18446), .ZN(O6646));
  INVX1 G49142 (.I(W6222), .ZN(W17646));
  INVX1 G49143 (.I(W30159), .ZN(O6613));
  INVX1 G49144 (.I(W32765), .ZN(O6612));
  INVX1 G49145 (.I(W17347), .ZN(O1422));
  INVX1 G49146 (.I(W26444), .ZN(O6611));
  INVX1 G49147 (.I(W31), .ZN(O6610));
  INVX1 G49148 (.I(W12886), .ZN(W17650));
  INVX1 G49149 (.I(W32162), .ZN(W33234));
  INVX1 G49150 (.I(W20074), .ZN(O6607));
  INVX1 G49151 (.I(W31871), .ZN(W33391));
  INVX1 G49152 (.I(W12228), .ZN(W17495));
  INVX1 G49153 (.I(W17753), .ZN(O6685));
  INVX1 G49154 (.I(W32528), .ZN(W33402));
  INVX1 G49155 (.I(W2096), .ZN(W33400));
  INVX1 G49156 (.I(W7409), .ZN(W33396));
  INVX1 G49157 (.I(W21866), .ZN(W33395));
  INVX1 G49158 (.I(W15777), .ZN(W17502));
  INVX1 G49159 (.I(W31987), .ZN(O6683));
  INVX1 G49160 (.I(I39), .ZN(O6682));
  INVX1 G49161 (.I(W11867), .ZN(W17493));
  INVX1 G49162 (.I(W21699), .ZN(O6681));
  INVX1 G49163 (.I(W647), .ZN(W17503));
  INVX1 G49164 (.I(W1931), .ZN(O6680));
  INVX1 G49165 (.I(W5828), .ZN(W33386));
  INVX1 G49166 (.I(W30803), .ZN(W33385));
  INVX1 G49167 (.I(W26811), .ZN(W33383));
  INVX1 G49168 (.I(W13797), .ZN(O6679));
  INVX1 G49169 (.I(W10393), .ZN(W17509));
  INVX1 G49170 (.I(W6769), .ZN(W17510));
  INVX1 G49171 (.I(W13341), .ZN(W33423));
  INVX1 G49172 (.I(W6435), .ZN(O1394));
  INVX1 G49173 (.I(W19438), .ZN(W33434));
  INVX1 G49174 (.I(W4473), .ZN(W33433));
  INVX1 G49175 (.I(W2798), .ZN(O1395));
  INVX1 G49176 (.I(I759), .ZN(O6696));
  INVX1 G49177 (.I(W13488), .ZN(W33430));
  INVX1 G49178 (.I(W23543), .ZN(O6694));
  INVX1 G49179 (.I(I184), .ZN(O6693));
  INVX1 G49180 (.I(W3114), .ZN(W17477));
  INVX1 G49181 (.I(W6238), .ZN(W17511));
  INVX1 G49182 (.I(W5825), .ZN(W17480));
  INVX1 G49183 (.I(W402), .ZN(O6692));
  INVX1 G49184 (.I(W28859), .ZN(W33418));
  INVX1 G49185 (.I(W3577), .ZN(O6689));
  INVX1 G49186 (.I(W2132), .ZN(W33415));
  INVX1 G49187 (.I(W5419), .ZN(O6687));
  INVX1 G49188 (.I(W13137), .ZN(W17488));
  INVX1 G49189 (.I(W7542), .ZN(O1401));
  INVX1 G49190 (.I(W18492), .ZN(W33408));
  INVX1 G49191 (.I(W10644), .ZN(W17551));
  INVX1 G49192 (.I(W8780), .ZN(W17538));
  INVX1 G49193 (.I(W1195), .ZN(W17541));
  INVX1 G49194 (.I(W15803), .ZN(W33344));
  INVX1 G49195 (.I(W16135), .ZN(O6660));
  INVX1 G49196 (.I(W9600), .ZN(O1409));
  INVX1 G49197 (.I(W3074), .ZN(O1410));
  INVX1 G49198 (.I(W3520), .ZN(O6657));
  INVX1 G49199 (.I(W658), .ZN(W17550));
  INVX1 G49200 (.I(W5916), .ZN(O6656));
  INVX1 G49201 (.I(W16246), .ZN(W17537));
  INVX1 G49202 (.I(W9142), .ZN(W33335));
  INVX1 G49203 (.I(W14859), .ZN(O6653));
  INVX1 G49204 (.I(W14266), .ZN(W17556));
  INVX1 G49205 (.I(W19715), .ZN(O6651));
  INVX1 G49206 (.I(W16850), .ZN(W17559));
  INVX1 G49207 (.I(I1944), .ZN(O6649));
  INVX1 G49208 (.I(W15959), .ZN(O6648));
  INVX1 G49209 (.I(W3544), .ZN(W17562));
  INVX1 G49210 (.I(W17198), .ZN(O6647));
  INVX1 G49211 (.I(W14582), .ZN(W33362));
  INVX1 G49212 (.I(W8689), .ZN(W33376));
  INVX1 G49213 (.I(W11206), .ZN(W17515));
  INVX1 G49214 (.I(W28556), .ZN(W33372));
  INVX1 G49215 (.I(W12991), .ZN(W17517));
  INVX1 G49216 (.I(W88), .ZN(W17518));
  INVX1 G49217 (.I(I222), .ZN(W17521));
  INVX1 G49218 (.I(W15032), .ZN(W17523));
  INVX1 G49219 (.I(W648), .ZN(W33366));
  INVX1 G49220 (.I(W23668), .ZN(O6672));
  INVX1 G49221 (.I(W22717), .ZN(O6591));
  INVX1 G49222 (.I(W9057), .ZN(W17526));
  INVX1 G49223 (.I(W11762), .ZN(W17527));
  INVX1 G49224 (.I(W16664), .ZN(O6669));
  INVX1 G49225 (.I(W6532), .ZN(W17529));
  INVX1 G49226 (.I(W23302), .ZN(W33357));
  INVX1 G49227 (.I(W1398), .ZN(W17532));
  INVX1 G49228 (.I(W3435), .ZN(W17533));
  INVX1 G49229 (.I(W27320), .ZN(W33352));
  INVX1 G49230 (.I(I622), .ZN(O6664));
  INVX1 G49231 (.I(W8849), .ZN(W17833));
  INVX1 G49232 (.I(W15224), .ZN(O1451));
  INVX1 G49233 (.I(W10521), .ZN(O6521));
  INVX1 G49234 (.I(W29845), .ZN(W33053));
  INVX1 G49235 (.I(W14348), .ZN(W33052));
  INVX1 G49236 (.I(W16239), .ZN(W17826));
  INVX1 G49237 (.I(W13873), .ZN(O6520));
  INVX1 G49238 (.I(W1477), .ZN(W17830));
  INVX1 G49239 (.I(W2169), .ZN(O6519));
  INVX1 G49240 (.I(W21691), .ZN(W33045));
  INVX1 G49241 (.I(W11065), .ZN(O6517));
  INVX1 G49242 (.I(W14746), .ZN(W17821));
  INVX1 G49243 (.I(W1642), .ZN(W17834));
  INVX1 G49244 (.I(W2298), .ZN(W17836));
  INVX1 G49245 (.I(W3348), .ZN(W33035));
  INVX1 G49246 (.I(W385), .ZN(O6513));
  INVX1 G49247 (.I(W1799), .ZN(W33033));
  INVX1 G49248 (.I(W5192), .ZN(W33032));
  INVX1 G49249 (.I(W16001), .ZN(W33031));
  INVX1 G49250 (.I(W23289), .ZN(O6512));
  INVX1 G49251 (.I(W8848), .ZN(O6510));
  INVX1 G49252 (.I(W15191), .ZN(O6527));
  INVX1 G49253 (.I(W24355), .ZN(W33080));
  INVX1 G49254 (.I(W9188), .ZN(W33079));
  INVX1 G49255 (.I(W7680), .ZN(O1445));
  INVX1 G49256 (.I(W27233), .ZN(W33075));
  INVX1 G49257 (.I(W17731), .ZN(W33074));
  INVX1 G49258 (.I(W11735), .ZN(O1447));
  INVX1 G49259 (.I(W6094), .ZN(W17803));
  INVX1 G49260 (.I(W13327), .ZN(W17804));
  INVX1 G49261 (.I(W13662), .ZN(O1449));
  INVX1 G49262 (.I(W1033), .ZN(W33024));
  INVX1 G49263 (.I(W923), .ZN(W17810));
  INVX1 G49264 (.I(W28052), .ZN(O6526));
  INVX1 G49265 (.I(W2061), .ZN(W17813));
  INVX1 G49266 (.I(W24701), .ZN(W33063));
  INVX1 G49267 (.I(W16957), .ZN(O6525));
  INVX1 G49268 (.I(W8346), .ZN(W17817));
  INVX1 G49269 (.I(W13851), .ZN(W17818));
  INVX1 G49270 (.I(W2638), .ZN(W17819));
  INVX1 G49271 (.I(W4906), .ZN(W33057));
  INVX1 G49272 (.I(W6695), .ZN(W17897));
  INVX1 G49273 (.I(W4977), .ZN(W17878));
  INVX1 G49274 (.I(W3983), .ZN(O1461));
  INVX1 G49275 (.I(W31489), .ZN(W32984));
  INVX1 G49276 (.I(W27999), .ZN(W32983));
  INVX1 G49277 (.I(W10854), .ZN(O6485));
  INVX1 G49278 (.I(W12046), .ZN(W17892));
  INVX1 G49279 (.I(W9789), .ZN(W32975));
  INVX1 G49280 (.I(W13784), .ZN(W17895));
  INVX1 G49281 (.I(W32208), .ZN(O6481));
  INVX1 G49282 (.I(W18455), .ZN(W32989));
  INVX1 G49283 (.I(W13604), .ZN(O1466));
  INVX1 G49284 (.I(W8660), .ZN(W17901));
  INVX1 G49285 (.I(W15485), .ZN(O6479));
  INVX1 G49286 (.I(W13817), .ZN(O6478));
  INVX1 G49287 (.I(W17511), .ZN(W32966));
  INVX1 G49288 (.I(W30357), .ZN(O6477));
  INVX1 G49289 (.I(W9722), .ZN(O6475));
  INVX1 G49290 (.I(W1098), .ZN(W17905));
  INVX1 G49291 (.I(W15843), .ZN(W17908));
  INVX1 G49292 (.I(W15688), .ZN(O6502));
  INVX1 G49293 (.I(W16898), .ZN(W33021));
  INVX1 G49294 (.I(W4282), .ZN(W17852));
  INVX1 G49295 (.I(W29912), .ZN(O6506));
  INVX1 G49296 (.I(W15306), .ZN(W17854));
  INVX1 G49297 (.I(W24652), .ZN(W33014));
  INVX1 G49298 (.I(W13365), .ZN(W33013));
  INVX1 G49299 (.I(W11619), .ZN(W17856));
  INVX1 G49300 (.I(I1900), .ZN(W33010));
  INVX1 G49301 (.I(W15893), .ZN(W33009));
  INVX1 G49302 (.I(I1162), .ZN(W17787));
  INVX1 G49303 (.I(W3694), .ZN(W17859));
  INVX1 G49304 (.I(W6272), .ZN(W17862));
  INVX1 G49305 (.I(W480), .ZN(W33001));
  INVX1 G49306 (.I(W4522), .ZN(O6496));
  INVX1 G49307 (.I(W13621), .ZN(W17871));
  INVX1 G49308 (.I(W23663), .ZN(W32995));
  INVX1 G49309 (.I(W16699), .ZN(O6493));
  INVX1 G49310 (.I(W17048), .ZN(O1459));
  INVX1 G49311 (.I(W1688), .ZN(W32990));
  INVX1 G49312 (.I(W23999), .ZN(O6569));
  INVX1 G49313 (.I(W16570), .ZN(W17702));
  INVX1 G49314 (.I(W8580), .ZN(W17704));
  INVX1 G49315 (.I(W13426), .ZN(O6574));
  INVX1 G49316 (.I(W17896), .ZN(O6573));
  INVX1 G49317 (.I(W3470), .ZN(O6572));
  INVX1 G49318 (.I(W16040), .ZN(W17705));
  INVX1 G49319 (.I(W21625), .ZN(O6571));
  INVX1 G49320 (.I(W4756), .ZN(W33158));
  INVX1 G49321 (.I(W9743), .ZN(W17711));
  INVX1 G49322 (.I(W31105), .ZN(W33167));
  INVX1 G49323 (.I(W9135), .ZN(W17713));
  INVX1 G49324 (.I(W6365), .ZN(W17714));
  INVX1 G49325 (.I(W2213), .ZN(W33151));
  INVX1 G49326 (.I(W6787), .ZN(W17718));
  INVX1 G49327 (.I(W2669), .ZN(W17721));
  INVX1 G49328 (.I(W9270), .ZN(W17722));
  INVX1 G49329 (.I(W7072), .ZN(W17723));
  INVX1 G49330 (.I(W4436), .ZN(O6566));
  INVX1 G49331 (.I(W28335), .ZN(W33144));
  INVX1 G49332 (.I(W25421), .ZN(W33185));
  INVX1 G49333 (.I(W6872), .ZN(W33198));
  INVX1 G49334 (.I(W21685), .ZN(O6590));
  INVX1 G49335 (.I(W5004), .ZN(W17678));
  INVX1 G49336 (.I(W14235), .ZN(O6587));
  INVX1 G49337 (.I(W7521), .ZN(W33193));
  INVX1 G49338 (.I(W14550), .ZN(W33191));
  INVX1 G49339 (.I(W2238), .ZN(W33190));
  INVX1 G49340 (.I(W5704), .ZN(O1430));
  INVX1 G49341 (.I(W15496), .ZN(O1431));
  INVX1 G49342 (.I(W17059), .ZN(O1436));
  INVX1 G49343 (.I(W11013), .ZN(O1432));
  INVX1 G49344 (.I(W16393), .ZN(W17689));
  INVX1 G49345 (.I(W32216), .ZN(W33177));
  INVX1 G49346 (.I(W11898), .ZN(W17698));
  INVX1 G49347 (.I(W12125), .ZN(W33173));
  INVX1 G49348 (.I(W8587), .ZN(W17699));
  INVX1 G49349 (.I(W7429), .ZN(W17700));
  INVX1 G49350 (.I(W17884), .ZN(W33170));
  INVX1 G49351 (.I(W14109), .ZN(W33168));
  INVX1 G49352 (.I(W32850), .ZN(W33099));
  INVX1 G49353 (.I(W17066), .ZN(W17761));
  INVX1 G49354 (.I(W10183), .ZN(W17764));
  INVX1 G49355 (.I(W14881), .ZN(O6546));
  INVX1 G49356 (.I(W26545), .ZN(O6544));
  INVX1 G49357 (.I(W12447), .ZN(W17768));
  INVX1 G49358 (.I(W13338), .ZN(O1441));
  INVX1 G49359 (.I(W21494), .ZN(W33103));
  INVX1 G49360 (.I(W7033), .ZN(O6542));
  INVX1 G49361 (.I(I46), .ZN(W33100));
  INVX1 G49362 (.I(W11860), .ZN(O1439));
  INVX1 G49363 (.I(I1030), .ZN(W17773));
  INVX1 G49364 (.I(W2947), .ZN(W33095));
  INVX1 G49365 (.I(W17706), .ZN(W17776));
  INVX1 G49366 (.I(W15701), .ZN(O1442));
  INVX1 G49367 (.I(W10230), .ZN(O6536));
  INVX1 G49368 (.I(I1215), .ZN(O6535));
  INVX1 G49369 (.I(W19966), .ZN(O6534));
  INVX1 G49370 (.I(W3771), .ZN(W17786));
  INVX1 G49371 (.I(I1224), .ZN(O6533));
  INVX1 G49372 (.I(W6358), .ZN(W33127));
  INVX1 G49373 (.I(W8424), .ZN(W33142));
  INVX1 G49374 (.I(W3471), .ZN(W33141));
  INVX1 G49375 (.I(W2128), .ZN(O1437));
  INVX1 G49376 (.I(W30135), .ZN(W33139));
  INVX1 G49377 (.I(W9513), .ZN(W17733));
  INVX1 G49378 (.I(W16157), .ZN(W17737));
  INVX1 G49379 (.I(W1382), .ZN(W17741));
  INVX1 G49380 (.I(W28228), .ZN(O6558));
  INVX1 G49381 (.I(I1201), .ZN(W17742));
  INVX1 G49382 (.I(I1263), .ZN(W17467));
  INVX1 G49383 (.I(W10441), .ZN(W17743));
  INVX1 G49384 (.I(W3396), .ZN(W17744));
  INVX1 G49385 (.I(I225), .ZN(W33124));
  INVX1 G49386 (.I(W13109), .ZN(O6556));
  INVX1 G49387 (.I(W15673), .ZN(W17745));
  INVX1 G49388 (.I(W835), .ZN(W17748));
  INVX1 G49389 (.I(W13524), .ZN(O1438));
  INVX1 G49390 (.I(W648), .ZN(O6554));
  INVX1 G49391 (.I(W16524), .ZN(W17753));
  INVX1 G49392 (.I(W14737), .ZN(O6867));
  INVX1 G49393 (.I(W7419), .ZN(O1326));
  INVX1 G49394 (.I(W13017), .ZN(W17133));
  INVX1 G49395 (.I(W1777), .ZN(W33771));
  INVX1 G49396 (.I(W4189), .ZN(O6871));
  INVX1 G49397 (.I(W15981), .ZN(O6870));
  INVX1 G49398 (.I(W11066), .ZN(W17137));
  INVX1 G49399 (.I(W5877), .ZN(W33762));
  INVX1 G49400 (.I(W16706), .ZN(W17143));
  INVX1 G49401 (.I(W13962), .ZN(O1332));
  INVX1 G49402 (.I(W14272), .ZN(W33759));
  INVX1 G49403 (.I(W12504), .ZN(W17123));
  INVX1 G49404 (.I(W18279), .ZN(W33757));
  INVX1 G49405 (.I(W2546), .ZN(W17145));
  INVX1 G49406 (.I(W13214), .ZN(W17147));
  INVX1 G49407 (.I(W11862), .ZN(W17148));
  INVX1 G49408 (.I(I1292), .ZN(O6866));
  INVX1 G49409 (.I(W28408), .ZN(W33752));
  INVX1 G49410 (.I(W25676), .ZN(W33751));
  INVX1 G49411 (.I(W26281), .ZN(W33750));
  INVX1 G49412 (.I(W15493), .ZN(W17149));
  INVX1 G49413 (.I(W4141), .ZN(O1320));
  INVX1 G49414 (.I(W3045), .ZN(O6896));
  INVX1 G49415 (.I(W13219), .ZN(W17099));
  INVX1 G49416 (.I(W5106), .ZN(W17102));
  INVX1 G49417 (.I(I48), .ZN(W33803));
  INVX1 G49418 (.I(W16031), .ZN(W17104));
  INVX1 G49419 (.I(I1076), .ZN(O1319));
  INVX1 G49420 (.I(W20141), .ZN(W33799));
  INVX1 G49421 (.I(W17008), .ZN(O6887));
  INVX1 G49422 (.I(W14246), .ZN(W17109));
  INVX1 G49423 (.I(W2312), .ZN(O1334));
  INVX1 G49424 (.I(W8089), .ZN(O6884));
  INVX1 G49425 (.I(W7988), .ZN(W17113));
  INVX1 G49426 (.I(W27010), .ZN(W33791));
  INVX1 G49427 (.I(W4230), .ZN(W17115));
  INVX1 G49428 (.I(W3312), .ZN(O6880));
  INVX1 G49429 (.I(W7450), .ZN(O6878));
  INVX1 G49430 (.I(W2082), .ZN(W17120));
  INVX1 G49431 (.I(W1371), .ZN(W33782));
  INVX1 G49432 (.I(W19979), .ZN(W33779));
  INVX1 G49433 (.I(W8604), .ZN(W17211));
  INVX1 G49434 (.I(W10846), .ZN(W17181));
  INVX1 G49435 (.I(W12963), .ZN(W17186));
  INVX1 G49436 (.I(W27531), .ZN(W33716));
  INVX1 G49437 (.I(I1462), .ZN(O6846));
  INVX1 G49438 (.I(W13257), .ZN(W33710));
  INVX1 G49439 (.I(W5613), .ZN(O6843));
  INVX1 G49440 (.I(W1699), .ZN(O1343));
  INVX1 G49441 (.I(W11468), .ZN(W33703));
  INVX1 G49442 (.I(W8759), .ZN(O1345));
  INVX1 G49443 (.I(W11370), .ZN(O6850));
  INVX1 G49444 (.I(W17916), .ZN(O6838));
  INVX1 G49445 (.I(I1126), .ZN(W33696));
  INVX1 G49446 (.I(W1593), .ZN(W17215));
  INVX1 G49447 (.I(W14987), .ZN(W17217));
  INVX1 G49448 (.I(W4985), .ZN(O6837));
  INVX1 G49449 (.I(I153), .ZN(O6836));
  INVX1 G49450 (.I(W13861), .ZN(O6835));
  INVX1 G49451 (.I(W31470), .ZN(O6834));
  INVX1 G49452 (.I(W29895), .ZN(W33687));
  INVX1 G49453 (.I(W13391), .ZN(O6858));
  INVX1 G49454 (.I(W4613), .ZN(W33746));
  INVX1 G49455 (.I(W26491), .ZN(W33745));
  INVX1 G49456 (.I(W11840), .ZN(O1335));
  INVX1 G49457 (.I(W4798), .ZN(W17157));
  INVX1 G49458 (.I(W19140), .ZN(W33739));
  INVX1 G49459 (.I(W9031), .ZN(O6861));
  INVX1 G49460 (.I(W27723), .ZN(W33737));
  INVX1 G49461 (.I(W7931), .ZN(O1337));
  INVX1 G49462 (.I(W24503), .ZN(O6859));
  INVX1 G49463 (.I(W5471), .ZN(O1317));
  INVX1 G49464 (.I(W26897), .ZN(O6857));
  INVX1 G49465 (.I(W14536), .ZN(W17162));
  INVX1 G49466 (.I(W26592), .ZN(W33729));
  INVX1 G49467 (.I(W27908), .ZN(O6854));
  INVX1 G49468 (.I(W6602), .ZN(W17167));
  INVX1 G49469 (.I(W13044), .ZN(O6853));
  INVX1 G49470 (.I(W9358), .ZN(O1339));
  INVX1 G49471 (.I(W2850), .ZN(W17175));
  INVX1 G49472 (.I(W15157), .ZN(W17178));
  INVX1 G49473 (.I(W4663), .ZN(W17036));
  INVX1 G49474 (.I(W10729), .ZN(W17018));
  INVX1 G49475 (.I(W649), .ZN(O1301));
  INVX1 G49476 (.I(W1184), .ZN(W17021));
  INVX1 G49477 (.I(W10427), .ZN(W17028));
  INVX1 G49478 (.I(W2863), .ZN(O6936));
  INVX1 G49479 (.I(W13448), .ZN(O1302));
  INVX1 G49480 (.I(W31475), .ZN(W33884));
  INVX1 G49481 (.I(I1848), .ZN(O1303));
  INVX1 G49482 (.I(W14763), .ZN(W33878));
  INVX1 G49483 (.I(W29894), .ZN(O6941));
  INVX1 G49484 (.I(W11296), .ZN(W33876));
  INVX1 G49485 (.I(W13816), .ZN(O6928));
  INVX1 G49486 (.I(W13399), .ZN(W17038));
  INVX1 G49487 (.I(W1117), .ZN(W17041));
  INVX1 G49488 (.I(W8136), .ZN(W17042));
  INVX1 G49489 (.I(W6327), .ZN(W33870));
  INVX1 G49490 (.I(W20575), .ZN(W33868));
  INVX1 G49491 (.I(W5396), .ZN(W17045));
  INVX1 G49492 (.I(W31474), .ZN(W33865));
  INVX1 G49493 (.I(W15955), .ZN(W17004));
  INVX1 G49494 (.I(W32480), .ZN(O6959));
  INVX1 G49495 (.I(W26816), .ZN(O6957));
  INVX1 G49496 (.I(W7129), .ZN(W33920));
  INVX1 G49497 (.I(W33376), .ZN(O6956));
  INVX1 G49498 (.I(W16982), .ZN(O1296));
  INVX1 G49499 (.I(W1962), .ZN(O1297));
  INVX1 G49500 (.I(W6834), .ZN(O6951));
  INVX1 G49501 (.I(W17415), .ZN(W33912));
  INVX1 G49502 (.I(W33307), .ZN(W33910));
  INVX1 G49503 (.I(W14285), .ZN(W33863));
  INVX1 G49504 (.I(W3241), .ZN(W17005));
  INVX1 G49505 (.I(W191), .ZN(W33907));
  INVX1 G49506 (.I(W2008), .ZN(O1299));
  INVX1 G49507 (.I(W14553), .ZN(W17007));
  INVX1 G49508 (.I(W1543), .ZN(W17011));
  INVX1 G49509 (.I(W6632), .ZN(W17013));
  INVX1 G49510 (.I(W15630), .ZN(O6944));
  INVX1 G49511 (.I(I898), .ZN(W17014));
  INVX1 G49512 (.I(W21101), .ZN(W33896));
  INVX1 G49513 (.I(W5240), .ZN(O6905));
  INVX1 G49514 (.I(W2368), .ZN(O1313));
  INVX1 G49515 (.I(W18376), .ZN(O6911));
  INVX1 G49516 (.I(W20862), .ZN(O6910));
  INVX1 G49517 (.I(W24306), .ZN(O6909));
  INVX1 G49518 (.I(W13313), .ZN(W17085));
  INVX1 G49519 (.I(W15989), .ZN(W33827));
  INVX1 G49520 (.I(I1426), .ZN(W17086));
  INVX1 G49521 (.I(W33466), .ZN(O6907));
  INVX1 G49522 (.I(W26835), .ZN(O6906));
  INVX1 G49523 (.I(W14072), .ZN(W17078));
  INVX1 G49524 (.I(W9769), .ZN(O6904));
  INVX1 G49525 (.I(W14272), .ZN(O6903));
  INVX1 G49526 (.I(W15049), .ZN(W17090));
  INVX1 G49527 (.I(W18002), .ZN(W33817));
  INVX1 G49528 (.I(W21413), .ZN(O6901));
  INVX1 G49529 (.I(W4314), .ZN(O6900));
  INVX1 G49530 (.I(W806), .ZN(W17091));
  INVX1 G49531 (.I(W14308), .ZN(O1316));
  INVX1 G49532 (.I(W15182), .ZN(W17094));
  INVX1 G49533 (.I(W1645), .ZN(W17061));
  INVX1 G49534 (.I(W7802), .ZN(W17048));
  INVX1 G49535 (.I(W7669), .ZN(W17050));
  INVX1 G49536 (.I(W1854), .ZN(W33860));
  INVX1 G49537 (.I(W435), .ZN(O1305));
  INVX1 G49538 (.I(W13494), .ZN(W33858));
  INVX1 G49539 (.I(W6435), .ZN(W17053));
  INVX1 G49540 (.I(W16971), .ZN(W17058));
  INVX1 G49541 (.I(W12114), .ZN(O6919));
  INVX1 G49542 (.I(W22631), .ZN(O6918));
  INVX1 G49543 (.I(W21855), .ZN(W33686));
  INVX1 G49544 (.I(W4167), .ZN(O1307));
  INVX1 G49545 (.I(W12721), .ZN(O1308));
  INVX1 G49546 (.I(W9733), .ZN(W33845));
  INVX1 G49547 (.I(W28942), .ZN(O6915));
  INVX1 G49548 (.I(W15193), .ZN(W17067));
  INVX1 G49549 (.I(W7316), .ZN(O1310));
  INVX1 G49550 (.I(W1611), .ZN(W17074));
  INVX1 G49551 (.I(W6721), .ZN(W33840));
  INVX1 G49552 (.I(W15551), .ZN(W17075));
  INVX1 G49553 (.I(W9734), .ZN(O1380));
  INVX1 G49554 (.I(W1213), .ZN(O1377));
  INVX1 G49555 (.I(W4055), .ZN(W33531));
  INVX1 G49556 (.I(W9568), .ZN(O1378));
  INVX1 G49557 (.I(W4686), .ZN(W33529));
  INVX1 G49558 (.I(W22191), .ZN(W33528));
  INVX1 G49559 (.I(W6030), .ZN(W17368));
  INVX1 G49560 (.I(W12935), .ZN(W17376));
  INVX1 G49561 (.I(W13438), .ZN(O6741));
  INVX1 G49562 (.I(W9042), .ZN(W33517));
  INVX1 G49563 (.I(W24634), .ZN(W33516));
  INVX1 G49564 (.I(W10332), .ZN(O6746));
  INVX1 G49565 (.I(W20259), .ZN(W33514));
  INVX1 G49566 (.I(W26775), .ZN(O6739));
  INVX1 G49567 (.I(W1527), .ZN(W33511));
  INVX1 G49568 (.I(W16066), .ZN(W17383));
  INVX1 G49569 (.I(W1719), .ZN(W17386));
  INVX1 G49570 (.I(W11787), .ZN(O6736));
  INVX1 G49571 (.I(W27150), .ZN(O6735));
  INVX1 G49572 (.I(W887), .ZN(W33506));
  INVX1 G49573 (.I(I1006), .ZN(W17387));
  INVX1 G49574 (.I(W11016), .ZN(O1375));
  INVX1 G49575 (.I(W16390), .ZN(W33564));
  INVX1 G49576 (.I(W4384), .ZN(W17331));
  INVX1 G49577 (.I(W3154), .ZN(O1373));
  INVX1 G49578 (.I(W25290), .ZN(W33559));
  INVX1 G49579 (.I(W9048), .ZN(W17337));
  INVX1 G49580 (.I(W12693), .ZN(W17338));
  INVX1 G49581 (.I(W11057), .ZN(W33555));
  INVX1 G49582 (.I(W10322), .ZN(W17341));
  INVX1 G49583 (.I(W5699), .ZN(W17342));
  INVX1 G49584 (.I(W16578), .ZN(O1381));
  INVX1 G49585 (.I(W13152), .ZN(W17345));
  INVX1 G49586 (.I(W33057), .ZN(O6755));
  INVX1 G49587 (.I(W11510), .ZN(W17346));
  INVX1 G49588 (.I(W7476), .ZN(W17347));
  INVX1 G49589 (.I(W11649), .ZN(O6753));
  INVX1 G49590 (.I(W6113), .ZN(W33542));
  INVX1 G49591 (.I(W31613), .ZN(O6750));
  INVX1 G49592 (.I(W1728), .ZN(W17355));
  INVX1 G49593 (.I(W117), .ZN(W17360));
  INVX1 G49594 (.I(W18944), .ZN(W33449));
  INVX1 G49595 (.I(W2336), .ZN(O1386));
  INVX1 G49596 (.I(W6236), .ZN(W17437));
  INVX1 G49597 (.I(W4985), .ZN(W17438));
  INVX1 G49598 (.I(I943), .ZN(O6713));
  INVX1 G49599 (.I(W19690), .ZN(O6710));
  INVX1 G49600 (.I(W2715), .ZN(O1391));
  INVX1 G49601 (.I(W12476), .ZN(O1392));
  INVX1 G49602 (.I(W13426), .ZN(O6705));
  INVX1 G49603 (.I(W14115), .ZN(W17456));
  INVX1 G49604 (.I(W12589), .ZN(W17421));
  INVX1 G49605 (.I(W11524), .ZN(W17457));
  INVX1 G49606 (.I(W11989), .ZN(W33446));
  INVX1 G49607 (.I(W3451), .ZN(O1393));
  INVX1 G49608 (.I(I893), .ZN(W17462));
  INVX1 G49609 (.I(W14382), .ZN(W17463));
  INVX1 G49610 (.I(W11397), .ZN(W33440));
  INVX1 G49611 (.I(W13084), .ZN(W17465));
  INVX1 G49612 (.I(W3704), .ZN(O6699));
  INVX1 G49613 (.I(W7000), .ZN(W17466));
  INVX1 G49614 (.I(W798), .ZN(W33489));
  INVX1 G49615 (.I(W8477), .ZN(W33503));
  INVX1 G49616 (.I(W1086), .ZN(W33501));
  INVX1 G49617 (.I(W2235), .ZN(W17394));
  INVX1 G49618 (.I(W12656), .ZN(W17396));
  INVX1 G49619 (.I(W136), .ZN(W17397));
  INVX1 G49620 (.I(W14984), .ZN(W17401));
  INVX1 G49621 (.I(W8329), .ZN(W33494));
  INVX1 G49622 (.I(W4255), .ZN(W33491));
  INVX1 G49623 (.I(W29562), .ZN(O6729));
  INVX1 G49624 (.I(W28585), .ZN(W33565));
  INVX1 G49625 (.I(W3162), .ZN(W17406));
  INVX1 G49626 (.I(W2658), .ZN(W17407));
  INVX1 G49627 (.I(W9059), .ZN(W17408));
  INVX1 G49628 (.I(W9717), .ZN(O6727));
  INVX1 G49629 (.I(W28572), .ZN(W33482));
  INVX1 G49630 (.I(W29805), .ZN(O6725));
  INVX1 G49631 (.I(I636), .ZN(W17415));
  INVX1 G49632 (.I(W16510), .ZN(O6722));
  INVX1 G49633 (.I(W5074), .ZN(W17420));
  INVX1 G49634 (.I(I1675), .ZN(W33641));
  INVX1 G49635 (.I(W105), .ZN(O1355));
  INVX1 G49636 (.I(W8741), .ZN(O1356));
  INVX1 G49637 (.I(W1085), .ZN(W17252));
  INVX1 G49638 (.I(W24006), .ZN(W33652));
  INVX1 G49639 (.I(W8197), .ZN(O6809));
  INVX1 G49640 (.I(W1899), .ZN(W17255));
  INVX1 G49641 (.I(W3109), .ZN(O6807));
  INVX1 G49642 (.I(W14722), .ZN(W17257));
  INVX1 G49643 (.I(W29734), .ZN(W33642));
  INVX1 G49644 (.I(W10705), .ZN(W33656));
  INVX1 G49645 (.I(I478), .ZN(W17264));
  INVX1 G49646 (.I(W22144), .ZN(O6802));
  INVX1 G49647 (.I(W25723), .ZN(O6801));
  INVX1 G49648 (.I(W15165), .ZN(W17267));
  INVX1 G49649 (.I(W2919), .ZN(W33634));
  INVX1 G49650 (.I(W5115), .ZN(O6800));
  INVX1 G49651 (.I(W1696), .ZN(O6799));
  INVX1 G49652 (.I(W30491), .ZN(O6796));
  INVX1 G49653 (.I(W24491), .ZN(O6794));
  INVX1 G49654 (.I(W14293), .ZN(O1351));
  INVX1 G49655 (.I(W3745), .ZN(W17223));
  INVX1 G49656 (.I(W7881), .ZN(O6832));
  INVX1 G49657 (.I(W8499), .ZN(W17224));
  INVX1 G49658 (.I(W28985), .ZN(O6830));
  INVX1 G49659 (.I(W5076), .ZN(W17225));
  INVX1 G49660 (.I(W4959), .ZN(W33678));
  INVX1 G49661 (.I(W1432), .ZN(O6827));
  INVX1 G49662 (.I(W5646), .ZN(W17232));
  INVX1 G49663 (.I(W26733), .ZN(O6825));
  INVX1 G49664 (.I(W2114), .ZN(W17272));
  INVX1 G49665 (.I(I1399), .ZN(O6822));
  INVX1 G49666 (.I(W2912), .ZN(W17238));
  INVX1 G49667 (.I(W1909), .ZN(W33668));
  INVX1 G49668 (.I(W5206), .ZN(W17239));
  INVX1 G49669 (.I(W32439), .ZN(O6820));
  INVX1 G49670 (.I(W4270), .ZN(W17244));
  INVX1 G49671 (.I(W13083), .ZN(W17246));
  INVX1 G49672 (.I(W27854), .ZN(O6814));
  INVX1 G49673 (.I(W2941), .ZN(W33657));
  INVX1 G49674 (.I(W6325), .ZN(O1371));
  INVX1 G49675 (.I(W33559), .ZN(W33590));
  INVX1 G49676 (.I(W15568), .ZN(O6772));
  INVX1 G49677 (.I(W3589), .ZN(W33588));
  INVX1 G49678 (.I(W4037), .ZN(W17311));
  INVX1 G49679 (.I(W30627), .ZN(W33586));
  INVX1 G49680 (.I(W16980), .ZN(O1369));
  INVX1 G49681 (.I(W2755), .ZN(W17314));
  INVX1 G49682 (.I(W11832), .ZN(O1370));
  INVX1 G49683 (.I(W8982), .ZN(W17317));
  INVX1 G49684 (.I(W8416), .ZN(W17308));
  INVX1 G49685 (.I(W10204), .ZN(W17323));
  INVX1 G49686 (.I(W16981), .ZN(W17325));
  INVX1 G49687 (.I(W11768), .ZN(O6766));
  INVX1 G49688 (.I(W15890), .ZN(W17328));
  INVX1 G49689 (.I(W32344), .ZN(W33571));
  INVX1 G49690 (.I(W17184), .ZN(O6765));
  INVX1 G49691 (.I(W28228), .ZN(W33568));
  INVX1 G49692 (.I(W4656), .ZN(O6764));
  INVX1 G49693 (.I(W5487), .ZN(O1372));
  INVX1 G49694 (.I(W14967), .ZN(W17288));
  INVX1 G49695 (.I(W32731), .ZN(O6792));
  INVX1 G49696 (.I(W10020), .ZN(W17275));
  INVX1 G49697 (.I(W3498), .ZN(W17276));
  INVX1 G49698 (.I(W9263), .ZN(W17278));
  INVX1 G49699 (.I(W1506), .ZN(W17280));
  INVX1 G49700 (.I(W4667), .ZN(W33617));
  INVX1 G49701 (.I(W6917), .ZN(W17285));
  INVX1 G49702 (.I(W18857), .ZN(O6786));
  INVX1 G49703 (.I(W17021), .ZN(W17287));
  INVX1 G49704 (.I(W12271), .ZN(W15945));
  INVX1 G49705 (.I(W11340), .ZN(O6784));
  INVX1 G49706 (.I(W24474), .ZN(W33605));
  INVX1 G49707 (.I(W14973), .ZN(W33603));
  INVX1 G49708 (.I(W102), .ZN(O1363));
  INVX1 G49709 (.I(W18396), .ZN(O6779));
  INVX1 G49710 (.I(W676), .ZN(O6778));
  INVX1 G49711 (.I(W5600), .ZN(W33598));
  INVX1 G49712 (.I(W7029), .ZN(O6773));
  INVX1 G49713 (.I(I164), .ZN(W33592));
  INVX1 G49714 (.I(W7416), .ZN(W14617));
  INVX1 G49715 (.I(W965), .ZN(O8263));
  INVX1 G49716 (.I(W9281), .ZN(W36216));
  INVX1 G49717 (.I(W12167), .ZN(O888));
  INVX1 G49718 (.I(W8967), .ZN(W14602));
  INVX1 G49719 (.I(W12819), .ZN(W14604));
  INVX1 G49720 (.I(W5943), .ZN(W14606));
  INVX1 G49721 (.I(W12052), .ZN(W14607));
  INVX1 G49722 (.I(W4874), .ZN(W36208));
  INVX1 G49723 (.I(W1426), .ZN(W36205));
  INVX1 G49724 (.I(W10975), .ZN(O8257));
  INVX1 G49725 (.I(W11828), .ZN(W14595));
  INVX1 G49726 (.I(W36065), .ZN(O8255));
  INVX1 G49727 (.I(W9325), .ZN(W14619));
  INVX1 G49728 (.I(W2878), .ZN(W14622));
  INVX1 G49729 (.I(W2776), .ZN(W14623));
  INVX1 G49730 (.I(I532), .ZN(O8253));
  INVX1 G49731 (.I(W7312), .ZN(W14624));
  INVX1 G49732 (.I(W7996), .ZN(W14626));
  INVX1 G49733 (.I(W9928), .ZN(W14627));
  INVX1 G49734 (.I(W4229), .ZN(W36191));
  INVX1 G49735 (.I(W11197), .ZN(W14585));
  INVX1 G49736 (.I(W33409), .ZN(O8279));
  INVX1 G49737 (.I(W24205), .ZN(W36243));
  INVX1 G49738 (.I(W15362), .ZN(O8278));
  INVX1 G49739 (.I(W13272), .ZN(W14570));
  INVX1 G49740 (.I(W4842), .ZN(W14577));
  INVX1 G49741 (.I(W8365), .ZN(W36237));
  INVX1 G49742 (.I(W13110), .ZN(W14582));
  INVX1 G49743 (.I(W13240), .ZN(W14583));
  INVX1 G49744 (.I(W11802), .ZN(W14584));
  INVX1 G49745 (.I(W28182), .ZN(O8249));
  INVX1 G49746 (.I(W8372), .ZN(O8273));
  INVX1 G49747 (.I(W5643), .ZN(W14586));
  INVX1 G49748 (.I(W35432), .ZN(O8271));
  INVX1 G49749 (.I(W5838), .ZN(W14588));
  INVX1 G49750 (.I(W7282), .ZN(W14589));
  INVX1 G49751 (.I(W16382), .ZN(O8269));
  INVX1 G49752 (.I(W8217), .ZN(O8268));
  INVX1 G49753 (.I(W6274), .ZN(O8267));
  INVX1 G49754 (.I(W352), .ZN(W14593));
  INVX1 G49755 (.I(W19232), .ZN(W36140));
  INVX1 G49756 (.I(W30874), .ZN(W36154));
  INVX1 G49757 (.I(W6560), .ZN(W14668));
  INVX1 G49758 (.I(W27534), .ZN(O8229));
  INVX1 G49759 (.I(W8504), .ZN(W14669));
  INVX1 G49760 (.I(W13225), .ZN(W36148));
  INVX1 G49761 (.I(W12458), .ZN(W14675));
  INVX1 G49762 (.I(W13246), .ZN(W36144));
  INVX1 G49763 (.I(W948), .ZN(W36142));
  INVX1 G49764 (.I(W30690), .ZN(O8225));
  INVX1 G49765 (.I(W12684), .ZN(O8232));
  INVX1 G49766 (.I(W9540), .ZN(O900));
  INVX1 G49767 (.I(W30844), .ZN(O8224));
  INVX1 G49768 (.I(W23781), .ZN(O8222));
  INVX1 G49769 (.I(W15768), .ZN(W36135));
  INVX1 G49770 (.I(W16115), .ZN(O8221));
  INVX1 G49771 (.I(W14463), .ZN(W14684));
  INVX1 G49772 (.I(W9237), .ZN(W36132));
  INVX1 G49773 (.I(W362), .ZN(W14685));
  INVX1 G49774 (.I(W8657), .ZN(W36130));
  INVX1 G49775 (.I(W7459), .ZN(W14641));
  INVX1 G49776 (.I(I329), .ZN(W14630));
  INVX1 G49777 (.I(W29978), .ZN(O8248));
  INVX1 G49778 (.I(W35851), .ZN(O8247));
  INVX1 G49779 (.I(W7491), .ZN(W36181));
  INVX1 G49780 (.I(W4586), .ZN(O893));
  INVX1 G49781 (.I(W7769), .ZN(W14637));
  INVX1 G49782 (.I(W3682), .ZN(W36177));
  INVX1 G49783 (.I(W17650), .ZN(W36175));
  INVX1 G49784 (.I(W32288), .ZN(O8242));
  INVX1 G49785 (.I(W5481), .ZN(W36245));
  INVX1 G49786 (.I(W4707), .ZN(O894));
  INVX1 G49787 (.I(W8531), .ZN(W14644));
  INVX1 G49788 (.I(W10805), .ZN(W14647));
  INVX1 G49789 (.I(W7089), .ZN(W14648));
  INVX1 G49790 (.I(W2631), .ZN(W14651));
  INVX1 G49791 (.I(W11525), .ZN(W14656));
  INVX1 G49792 (.I(W6631), .ZN(W14657));
  INVX1 G49793 (.I(W17924), .ZN(W36160));
  INVX1 G49794 (.I(W125), .ZN(W14661));
  INVX1 G49795 (.I(W17572), .ZN(O8330));
  INVX1 G49796 (.I(I1748), .ZN(W14468));
  INVX1 G49797 (.I(W17515), .ZN(W36339));
  INVX1 G49798 (.I(W15911), .ZN(W36337));
  INVX1 G49799 (.I(W370), .ZN(W36336));
  INVX1 G49800 (.I(W14096), .ZN(W14475));
  INVX1 G49801 (.I(W11503), .ZN(O8333));
  INVX1 G49802 (.I(W4468), .ZN(W14481));
  INVX1 G49803 (.I(W634), .ZN(W36326));
  INVX1 G49804 (.I(W11710), .ZN(W14486));
  INVX1 G49805 (.I(W5556), .ZN(W14467));
  INVX1 G49806 (.I(W23881), .ZN(O8328));
  INVX1 G49807 (.I(W11997), .ZN(W36319));
  INVX1 G49808 (.I(W8081), .ZN(W36318));
  INVX1 G49809 (.I(W13142), .ZN(W36317));
  INVX1 G49810 (.I(W12859), .ZN(W14491));
  INVX1 G49811 (.I(W10054), .ZN(W14492));
  INVX1 G49812 (.I(W938), .ZN(W14495));
  INVX1 G49813 (.I(W10648), .ZN(O877));
  INVX1 G49814 (.I(W27359), .ZN(O8321));
  INVX1 G49815 (.I(W5727), .ZN(W36358));
  INVX1 G49816 (.I(W10456), .ZN(W14443));
  INVX1 G49817 (.I(W7887), .ZN(O8352));
  INVX1 G49818 (.I(W2040), .ZN(O8351));
  INVX1 G49819 (.I(W12368), .ZN(W14446));
  INVX1 G49820 (.I(W18922), .ZN(O8349));
  INVX1 G49821 (.I(W10128), .ZN(W14449));
  INVX1 G49822 (.I(W14703), .ZN(O8347));
  INVX1 G49823 (.I(W25065), .ZN(W36362));
  INVX1 G49824 (.I(W10359), .ZN(W14451));
  INVX1 G49825 (.I(W13442), .ZN(W14497));
  INVX1 G49826 (.I(W9914), .ZN(O873));
  INVX1 G49827 (.I(W3428), .ZN(W36353));
  INVX1 G49828 (.I(W11355), .ZN(O874));
  INVX1 G49829 (.I(W20471), .ZN(W36350));
  INVX1 G49830 (.I(W18856), .ZN(W36348));
  INVX1 G49831 (.I(W6577), .ZN(W14463));
  INVX1 G49832 (.I(W11915), .ZN(W14464));
  INVX1 G49833 (.I(W4684), .ZN(W14465));
  INVX1 G49834 (.I(W14192), .ZN(O875));
  INVX1 G49835 (.I(W2109), .ZN(O8291));
  INVX1 G49836 (.I(W4913), .ZN(W14534));
  INVX1 G49837 (.I(W11863), .ZN(W14535));
  INVX1 G49838 (.I(W16644), .ZN(W36277));
  INVX1 G49839 (.I(W3282), .ZN(O8297));
  INVX1 G49840 (.I(W11265), .ZN(O8296));
  INVX1 G49841 (.I(W31111), .ZN(O8295));
  INVX1 G49842 (.I(W23385), .ZN(O8294));
  INVX1 G49843 (.I(W4894), .ZN(W36270));
  INVX1 G49844 (.I(W6303), .ZN(O881));
  INVX1 G49845 (.I(W1433), .ZN(W14532));
  INVX1 G49846 (.I(W30291), .ZN(O8290));
  INVX1 G49847 (.I(W9609), .ZN(O8289));
  INVX1 G49848 (.I(W9213), .ZN(W14547));
  INVX1 G49849 (.I(W22422), .ZN(O8283));
  INVX1 G49850 (.I(W260), .ZN(O883));
  INVX1 G49851 (.I(W4773), .ZN(O884));
  INVX1 G49852 (.I(W20896), .ZN(O8281));
  INVX1 G49853 (.I(W14526), .ZN(W14561));
  INVX1 G49854 (.I(W9171), .ZN(W14565));
  INVX1 G49855 (.I(W9363), .ZN(W14519));
  INVX1 G49856 (.I(W33936), .ZN(O8319));
  INVX1 G49857 (.I(W5555), .ZN(W14504));
  INVX1 G49858 (.I(W538), .ZN(O8316));
  INVX1 G49859 (.I(W10215), .ZN(W14505));
  INVX1 G49860 (.I(W9807), .ZN(W14507));
  INVX1 G49861 (.I(W1052), .ZN(W14515));
  INVX1 G49862 (.I(W18308), .ZN(W36298));
  INVX1 G49863 (.I(W11518), .ZN(O880));
  INVX1 G49864 (.I(W34383), .ZN(W36295));
  INVX1 G49865 (.I(W14420), .ZN(W14688));
  INVX1 G49866 (.I(W5554), .ZN(O8309));
  INVX1 G49867 (.I(W9026), .ZN(W14521));
  INVX1 G49868 (.I(W965), .ZN(O8307));
  INVX1 G49869 (.I(W31719), .ZN(O8305));
  INVX1 G49870 (.I(W16630), .ZN(O8304));
  INVX1 G49871 (.I(I634), .ZN(W14526));
  INVX1 G49872 (.I(W8101), .ZN(W14527));
  INVX1 G49873 (.I(W6871), .ZN(W14529));
  INVX1 G49874 (.I(W1791), .ZN(W14531));
  INVX1 G49875 (.I(W22244), .ZN(O8118));
  INVX1 G49876 (.I(W8534), .ZN(W35987));
  INVX1 G49877 (.I(W17293), .ZN(W35986));
  INVX1 G49878 (.I(W7775), .ZN(W35984));
  INVX1 G49879 (.I(W9992), .ZN(O8126));
  INVX1 G49880 (.I(W2618), .ZN(W35982));
  INVX1 G49881 (.I(W12520), .ZN(W14820));
  INVX1 G49882 (.I(W33521), .ZN(O8125));
  INVX1 G49883 (.I(I1421), .ZN(W35978));
  INVX1 G49884 (.I(W21653), .ZN(O8122));
  INVX1 G49885 (.I(W5968), .ZN(W14827));
  INVX1 G49886 (.I(W9516), .ZN(W35988));
  INVX1 G49887 (.I(W10183), .ZN(W14834));
  INVX1 G49888 (.I(W8461), .ZN(W14838));
  INVX1 G49889 (.I(W13386), .ZN(O8114));
  INVX1 G49890 (.I(W28420), .ZN(O8113));
  INVX1 G49891 (.I(W30230), .ZN(W35962));
  INVX1 G49892 (.I(W26027), .ZN(W35961));
  INVX1 G49893 (.I(W35548), .ZN(O8111));
  INVX1 G49894 (.I(W12563), .ZN(O925));
  INVX1 G49895 (.I(W12891), .ZN(O8110));
  INVX1 G49896 (.I(W14125), .ZN(W14808));
  INVX1 G49897 (.I(W24818), .ZN(W36011));
  INVX1 G49898 (.I(W8948), .ZN(W14799));
  INVX1 G49899 (.I(W9034), .ZN(W14800));
  INVX1 G49900 (.I(W27592), .ZN(O8140));
  INVX1 G49901 (.I(W2115), .ZN(W14801));
  INVX1 G49902 (.I(W6664), .ZN(W14802));
  INVX1 G49903 (.I(W15495), .ZN(O8137));
  INVX1 G49904 (.I(W8988), .ZN(W14807));
  INVX1 G49905 (.I(W19005), .ZN(O8135));
  INVX1 G49906 (.I(W13103), .ZN(O8108));
  INVX1 G49907 (.I(W3685), .ZN(W14809));
  INVX1 G49908 (.I(W13845), .ZN(O8133));
  INVX1 G49909 (.I(W23362), .ZN(O8131));
  INVX1 G49910 (.I(W6872), .ZN(W14811));
  INVX1 G49911 (.I(W34157), .ZN(W35994));
  INVX1 G49912 (.I(W33133), .ZN(O8130));
  INVX1 G49913 (.I(W5585), .ZN(W14817));
  INVX1 G49914 (.I(I409), .ZN(O8128));
  INVX1 G49915 (.I(I661), .ZN(O922));
  INVX1 G49916 (.I(I1608), .ZN(W14882));
  INVX1 G49917 (.I(W33506), .ZN(O8091));
  INVX1 G49918 (.I(I1660), .ZN(W14870));
  INVX1 G49919 (.I(W33773), .ZN(O8088));
  INVX1 G49920 (.I(W6061), .ZN(W14875));
  INVX1 G49921 (.I(I1760), .ZN(W14878));
  INVX1 G49922 (.I(W28936), .ZN(O8086));
  INVX1 G49923 (.I(W11093), .ZN(W14879));
  INVX1 G49924 (.I(I1636), .ZN(O8084));
  INVX1 G49925 (.I(W29976), .ZN(O8083));
  INVX1 G49926 (.I(W30690), .ZN(O8092));
  INVX1 G49927 (.I(W2170), .ZN(O8081));
  INVX1 G49928 (.I(W549), .ZN(W14886));
  INVX1 G49929 (.I(W1468), .ZN(W14888));
  INVX1 G49930 (.I(W8906), .ZN(W35907));
  INVX1 G49931 (.I(W1891), .ZN(O8077));
  INVX1 G49932 (.I(W26399), .ZN(W35899));
  INVX1 G49933 (.I(W16969), .ZN(O8071));
  INVX1 G49934 (.I(W5382), .ZN(O8070));
  INVX1 G49935 (.I(W14096), .ZN(O8069));
  INVX1 G49936 (.I(W9656), .ZN(W35939));
  INVX1 G49937 (.I(W11942), .ZN(W14851));
  INVX1 G49938 (.I(W6938), .ZN(W14854));
  INVX1 G49939 (.I(W15430), .ZN(O8105));
  INVX1 G49940 (.I(W14985), .ZN(O8104));
  INVX1 G49941 (.I(W8443), .ZN(W35947));
  INVX1 G49942 (.I(W16867), .ZN(W35944));
  INVX1 G49943 (.I(W1706), .ZN(O8102));
  INVX1 G49944 (.I(W34133), .ZN(W35941));
  INVX1 G49945 (.I(W12903), .ZN(W14859));
  INVX1 G49946 (.I(W19907), .ZN(O8143));
  INVX1 G49947 (.I(W7242), .ZN(W14861));
  INVX1 G49948 (.I(W14851), .ZN(W14862));
  INVX1 G49949 (.I(W10488), .ZN(O8096));
  INVX1 G49950 (.I(W14500), .ZN(W14863));
  INVX1 G49951 (.I(W20806), .ZN(O8095));
  INVX1 G49952 (.I(W5496), .ZN(W14864));
  INVX1 G49953 (.I(W7042), .ZN(O8094));
  INVX1 G49954 (.I(I1748), .ZN(W14865));
  INVX1 G49955 (.I(W4606), .ZN(W14867));
  INVX1 G49956 (.I(W26194), .ZN(O8195));
  INVX1 G49957 (.I(I1714), .ZN(O8200));
  INVX1 G49958 (.I(W27139), .ZN(W36099));
  INVX1 G49959 (.I(W14297), .ZN(W14714));
  INVX1 G49960 (.I(W2984), .ZN(O8198));
  INVX1 G49961 (.I(W7605), .ZN(W14716));
  INVX1 G49962 (.I(W3291), .ZN(O907));
  INVX1 G49963 (.I(W11243), .ZN(W14719));
  INVX1 G49964 (.I(W34848), .ZN(W36093));
  INVX1 G49965 (.I(W14669), .ZN(W36091));
  INVX1 G49966 (.I(W7446), .ZN(O8202));
  INVX1 G49967 (.I(W165), .ZN(O8193));
  INVX1 G49968 (.I(W10925), .ZN(W14724));
  INVX1 G49969 (.I(W28457), .ZN(O8191));
  INVX1 G49970 (.I(W1345), .ZN(W14726));
  INVX1 G49971 (.I(W27828), .ZN(O8190));
  INVX1 G49972 (.I(W11610), .ZN(W14728));
  INVX1 G49973 (.I(W2382), .ZN(W14729));
  INVX1 G49974 (.I(W34947), .ZN(W36080));
  INVX1 G49975 (.I(W5062), .ZN(W14730));
  INVX1 G49976 (.I(W12577), .ZN(W14696));
  INVX1 G49977 (.I(W20218), .ZN(O8219));
  INVX1 G49978 (.I(I410), .ZN(W14689));
  INVX1 G49979 (.I(W6923), .ZN(W14691));
  INVX1 G49980 (.I(W29587), .ZN(W36125));
  INVX1 G49981 (.I(I1357), .ZN(O8216));
  INVX1 G49982 (.I(W9966), .ZN(W36123));
  INVX1 G49983 (.I(W14553), .ZN(W14692));
  INVX1 G49984 (.I(I1189), .ZN(W14694));
  INVX1 G49985 (.I(W7462), .ZN(W36118));
  INVX1 G49986 (.I(W13977), .ZN(W14731));
  INVX1 G49987 (.I(I1808), .ZN(W14698));
  INVX1 G49988 (.I(W8333), .ZN(W14701));
  INVX1 G49989 (.I(W10070), .ZN(W14702));
  INVX1 G49990 (.I(W5811), .ZN(W14703));
  INVX1 G49991 (.I(W2141), .ZN(W14705));
  INVX1 G49992 (.I(I1557), .ZN(O8204));
  INVX1 G49993 (.I(W30917), .ZN(W36107));
  INVX1 G49994 (.I(W13099), .ZN(W14710));
  INVX1 G49995 (.I(W4943), .ZN(W14712));
  INVX1 G49996 (.I(W17162), .ZN(O8154));
  INVX1 G49997 (.I(W11310), .ZN(W14761));
  INVX1 G49998 (.I(W546), .ZN(W14764));
  INVX1 G49999 (.I(W24880), .ZN(W36041));
  INVX1 G50000 (.I(W4875), .ZN(W14769));
  INVX1 G50001 (.I(W7277), .ZN(W14775));
  INVX1 G50002 (.I(W12221), .ZN(W14778));
  INVX1 G50003 (.I(W13464), .ZN(W14780));
  INVX1 G50004 (.I(I260), .ZN(O8156));
  INVX1 G50005 (.I(W861), .ZN(O8155));
  INVX1 G50006 (.I(W11169), .ZN(W14758));
  INVX1 G50007 (.I(W8101), .ZN(O915));
  INVX1 G50008 (.I(W12943), .ZN(O8152));
  INVX1 G50009 (.I(W7526), .ZN(W14788));
  INVX1 G50010 (.I(W11758), .ZN(W14789));
  INVX1 G50011 (.I(W13160), .ZN(O8146));
  INVX1 G50012 (.I(W5236), .ZN(W14794));
  INVX1 G50013 (.I(W14048), .ZN(W36015));
  INVX1 G50014 (.I(W31564), .ZN(O8145));
  INVX1 G50015 (.I(W8556), .ZN(O918));
  INVX1 G50016 (.I(W3254), .ZN(O910));
  INVX1 G50017 (.I(W789), .ZN(W36077));
  INVX1 G50018 (.I(W3768), .ZN(W36076));
  INVX1 G50019 (.I(I362), .ZN(O8186));
  INVX1 G50020 (.I(W33863), .ZN(O8185));
  INVX1 G50021 (.I(W2850), .ZN(W14735));
  INVX1 G50022 (.I(W18198), .ZN(O8183));
  INVX1 G50023 (.I(W11685), .ZN(W14737));
  INVX1 G50024 (.I(W8389), .ZN(W14738));
  INVX1 G50025 (.I(W31194), .ZN(O8181));
  INVX1 G50026 (.I(W32583), .ZN(O8355));
  INVX1 G50027 (.I(W1112), .ZN(W14740));
  INVX1 G50028 (.I(W5682), .ZN(W14743));
  INVX1 G50029 (.I(W1924), .ZN(W36060));
  INVX1 G50030 (.I(W13418), .ZN(O8178));
  INVX1 G50031 (.I(W23810), .ZN(O8177));
  INVX1 G50032 (.I(W4471), .ZN(W14748));
  INVX1 G50033 (.I(W12042), .ZN(W14751));
  INVX1 G50034 (.I(W23468), .ZN(O8172));
  INVX1 G50035 (.I(W4519), .ZN(O8171));
  INVX1 G50036 (.I(W1116), .ZN(W14129));
  INVX1 G50037 (.I(W7213), .ZN(W14116));
  INVX1 G50038 (.I(W7093), .ZN(W14118));
  INVX1 G50039 (.I(W26923), .ZN(W36709));
  INVX1 G50040 (.I(W11966), .ZN(W36708));
  INVX1 G50041 (.I(W1415), .ZN(W14119));
  INVX1 G50042 (.I(W2363), .ZN(W14120));
  INVX1 G50043 (.I(W8639), .ZN(O827));
  INVX1 G50044 (.I(W32106), .ZN(W36703));
  INVX1 G50045 (.I(W9436), .ZN(O8552));
  INVX1 G50046 (.I(I831), .ZN(O8551));
  INVX1 G50047 (.I(W7226), .ZN(W14115));
  INVX1 G50048 (.I(W22395), .ZN(W36696));
  INVX1 G50049 (.I(I1533), .ZN(W14130));
  INVX1 G50050 (.I(W4880), .ZN(W14132));
  INVX1 G50051 (.I(I1215), .ZN(W14139));
  INVX1 G50052 (.I(W3870), .ZN(W14140));
  INVX1 G50053 (.I(W10552), .ZN(W14142));
  INVX1 G50054 (.I(W31711), .ZN(O8542));
  INVX1 G50055 (.I(W29074), .ZN(W36687));
  INVX1 G50056 (.I(W13494), .ZN(O8538));
  INVX1 G50057 (.I(W5936), .ZN(W36729));
  INVX1 G50058 (.I(W7976), .ZN(W14085));
  INVX1 G50059 (.I(W4569), .ZN(O8570));
  INVX1 G50060 (.I(W28587), .ZN(O8569));
  INVX1 G50061 (.I(W10390), .ZN(W14086));
  INVX1 G50062 (.I(W26740), .ZN(W36734));
  INVX1 G50063 (.I(I1790), .ZN(W14092));
  INVX1 G50064 (.I(W18949), .ZN(O8567));
  INVX1 G50065 (.I(W8484), .ZN(W36731));
  INVX1 G50066 (.I(I1575), .ZN(W14093));
  INVX1 G50067 (.I(W14960), .ZN(W36678));
  INVX1 G50068 (.I(W29511), .ZN(O8565));
  INVX1 G50069 (.I(W9746), .ZN(W14098));
  INVX1 G50070 (.I(W8096), .ZN(W36725));
  INVX1 G50071 (.I(W1000), .ZN(W14103));
  INVX1 G50072 (.I(W33430), .ZN(O8562));
  INVX1 G50073 (.I(W30165), .ZN(W36720));
  INVX1 G50074 (.I(W5965), .ZN(W14107));
  INVX1 G50075 (.I(W29530), .ZN(W36718));
  INVX1 G50076 (.I(W7212), .ZN(W14109));
  INVX1 G50077 (.I(W6567), .ZN(W14182));
  INVX1 G50078 (.I(W7317), .ZN(W14173));
  INVX1 G50079 (.I(W30370), .ZN(W36649));
  INVX1 G50080 (.I(W13996), .ZN(W14174));
  INVX1 G50081 (.I(W4829), .ZN(W14176));
  INVX1 G50082 (.I(W3048), .ZN(O8522));
  INVX1 G50083 (.I(W25977), .ZN(W36644));
  INVX1 G50084 (.I(W1724), .ZN(W14178));
  INVX1 G50085 (.I(W13897), .ZN(W14179));
  INVX1 G50086 (.I(W32085), .ZN(O8520));
  INVX1 G50087 (.I(W23205), .ZN(O8523));
  INVX1 G50088 (.I(W8760), .ZN(W14183));
  INVX1 G50089 (.I(W8605), .ZN(W14190));
  INVX1 G50090 (.I(W10087), .ZN(O8515));
  INVX1 G50091 (.I(W6366), .ZN(W14194));
  INVX1 G50092 (.I(W4579), .ZN(O840));
  INVX1 G50093 (.I(W7807), .ZN(W14198));
  INVX1 G50094 (.I(W363), .ZN(O841));
  INVX1 G50095 (.I(W26777), .ZN(O8511));
  INVX1 G50096 (.I(W12221), .ZN(O8508));
  INVX1 G50097 (.I(W4614), .ZN(W14160));
  INVX1 G50098 (.I(W3532), .ZN(O832));
  INVX1 G50099 (.I(W19569), .ZN(O8534));
  INVX1 G50100 (.I(W15355), .ZN(W36674));
  INVX1 G50101 (.I(W13352), .ZN(W36672));
  INVX1 G50102 (.I(W10981), .ZN(W14156));
  INVX1 G50103 (.I(W11895), .ZN(W14158));
  INVX1 G50104 (.I(W21759), .ZN(O8532));
  INVX1 G50105 (.I(W11468), .ZN(W14159));
  INVX1 G50106 (.I(W11159), .ZN(W36667));
  INVX1 G50107 (.I(W3050), .ZN(O8572));
  INVX1 G50108 (.I(W2384), .ZN(W14163));
  INVX1 G50109 (.I(W23109), .ZN(W36663));
  INVX1 G50110 (.I(W12503), .ZN(W14164));
  INVX1 G50111 (.I(W5083), .ZN(W14166));
  INVX1 G50112 (.I(W11469), .ZN(O8527));
  INVX1 G50113 (.I(W9573), .ZN(O8526));
  INVX1 G50114 (.I(I290), .ZN(W14169));
  INVX1 G50115 (.I(W7881), .ZN(O8524));
  INVX1 G50116 (.I(W6545), .ZN(W14171));
  INVX1 G50117 (.I(W19883), .ZN(W36821));
  INVX1 G50118 (.I(W8642), .ZN(O813));
  INVX1 G50119 (.I(W1078), .ZN(W13992));
  INVX1 G50120 (.I(W6286), .ZN(O8618));
  INVX1 G50121 (.I(W16766), .ZN(O8617));
  INVX1 G50122 (.I(W33743), .ZN(W36827));
  INVX1 G50123 (.I(W30561), .ZN(O8616));
  INVX1 G50124 (.I(W1072), .ZN(O814));
  INVX1 G50125 (.I(W5381), .ZN(W13998));
  INVX1 G50126 (.I(W33751), .ZN(O8614));
  INVX1 G50127 (.I(W2856), .ZN(W13990));
  INVX1 G50128 (.I(W11663), .ZN(W13999));
  INVX1 G50129 (.I(W7628), .ZN(W14001));
  INVX1 G50130 (.I(W35636), .ZN(O8611));
  INVX1 G50131 (.I(W9441), .ZN(W14003));
  INVX1 G50132 (.I(W21413), .ZN(O8609));
  INVX1 G50133 (.I(W1910), .ZN(W14005));
  INVX1 G50134 (.I(W13955), .ZN(W36813));
  INVX1 G50135 (.I(W7411), .ZN(O8608));
  INVX1 G50136 (.I(W16233), .ZN(W36811));
  INVX1 G50137 (.I(W33167), .ZN(W36843));
  INVX1 G50138 (.I(W9853), .ZN(W36859));
  INVX1 G50139 (.I(W7252), .ZN(W13955));
  INVX1 G50140 (.I(W1704), .ZN(O8638));
  INVX1 G50141 (.I(W9918), .ZN(W13959));
  INVX1 G50142 (.I(W4304), .ZN(W13962));
  INVX1 G50143 (.I(W3709), .ZN(W13963));
  INVX1 G50144 (.I(I412), .ZN(W13969));
  INVX1 G50145 (.I(W11497), .ZN(W13971));
  INVX1 G50146 (.I(W4608), .ZN(W13975));
  INVX1 G50147 (.I(W7787), .ZN(W14007));
  INVX1 G50148 (.I(I278), .ZN(W36842));
  INVX1 G50149 (.I(W7858), .ZN(W13978));
  INVX1 G50150 (.I(W12814), .ZN(W13980));
  INVX1 G50151 (.I(W24802), .ZN(O8627));
  INVX1 G50152 (.I(W35362), .ZN(O8625));
  INVX1 G50153 (.I(W31509), .ZN(O8624));
  INVX1 G50154 (.I(W1409), .ZN(W13985));
  INVX1 G50155 (.I(W10485), .ZN(O8622));
  INVX1 G50156 (.I(W9611), .ZN(W13987));
  INVX1 G50157 (.I(W15088), .ZN(O8579));
  INVX1 G50158 (.I(W2421), .ZN(W14059));
  INVX1 G50159 (.I(W12085), .ZN(O8587));
  INVX1 G50160 (.I(W16212), .ZN(W36768));
  INVX1 G50161 (.I(W10417), .ZN(O8585));
  INVX1 G50162 (.I(W3046), .ZN(W14062));
  INVX1 G50163 (.I(W6763), .ZN(W14063));
  INVX1 G50164 (.I(W8402), .ZN(W14064));
  INVX1 G50165 (.I(I725), .ZN(W14066));
  INVX1 G50166 (.I(W26469), .ZN(W36757));
  INVX1 G50167 (.I(W2935), .ZN(W14057));
  INVX1 G50168 (.I(I1622), .ZN(W36755));
  INVX1 G50169 (.I(W2049), .ZN(W14070));
  INVX1 G50170 (.I(W9976), .ZN(O8578));
  INVX1 G50171 (.I(W5250), .ZN(W14078));
  INVX1 G50172 (.I(I1927), .ZN(W14079));
  INVX1 G50173 (.I(W4608), .ZN(W14080));
  INVX1 G50174 (.I(W22749), .ZN(W36747));
  INVX1 G50175 (.I(I1140), .ZN(W14082));
  INVX1 G50176 (.I(W8536), .ZN(O822));
  INVX1 G50177 (.I(W9208), .ZN(W14029));
  INVX1 G50178 (.I(W18428), .ZN(W36809));
  INVX1 G50179 (.I(W24704), .ZN(W36805));
  INVX1 G50180 (.I(W7064), .ZN(W14016));
  INVX1 G50181 (.I(W11118), .ZN(O8606));
  INVX1 G50182 (.I(W13692), .ZN(W14021));
  INVX1 G50183 (.I(W33949), .ZN(O8602));
  INVX1 G50184 (.I(W13850), .ZN(W36798));
  INVX1 G50185 (.I(W35758), .ZN(W36795));
  INVX1 G50186 (.I(I198), .ZN(W14024));
  INVX1 G50187 (.I(W5160), .ZN(W14208));
  INVX1 G50188 (.I(W10945), .ZN(W36789));
  INVX1 G50189 (.I(W4281), .ZN(O8597));
  INVX1 G50190 (.I(W13806), .ZN(O8596));
  INVX1 G50191 (.I(W5230), .ZN(W14039));
  INVX1 G50192 (.I(W6262), .ZN(W14041));
  INVX1 G50193 (.I(W12069), .ZN(W14042));
  INVX1 G50194 (.I(W19197), .ZN(O8591));
  INVX1 G50195 (.I(W12704), .ZN(W14052));
  INVX1 G50196 (.I(W9138), .ZN(W14053));
  INVX1 G50197 (.I(W5538), .ZN(W36448));
  INVX1 G50198 (.I(W24716), .ZN(O8414));
  INVX1 G50199 (.I(W11063), .ZN(W14364));
  INVX1 G50200 (.I(I620), .ZN(W14365));
  INVX1 G50201 (.I(W287), .ZN(W14370));
  INVX1 G50202 (.I(I1096), .ZN(W14373));
  INVX1 G50203 (.I(W23585), .ZN(O8407));
  INVX1 G50204 (.I(W1277), .ZN(W36457));
  INVX1 G50205 (.I(W3314), .ZN(O8405));
  INVX1 G50206 (.I(W11769), .ZN(W36452));
  INVX1 G50207 (.I(W3425), .ZN(O860));
  INVX1 G50208 (.I(W12047), .ZN(W14359));
  INVX1 G50209 (.I(W31768), .ZN(O8402));
  INVX1 G50210 (.I(W12457), .ZN(O8401));
  INVX1 G50211 (.I(W2865), .ZN(W36445));
  INVX1 G50212 (.I(W24366), .ZN(W36444));
  INVX1 G50213 (.I(W23240), .ZN(W36443));
  INVX1 G50214 (.I(W7185), .ZN(O861));
  INVX1 G50215 (.I(W33200), .ZN(W36440));
  INVX1 G50216 (.I(W7868), .ZN(O862));
  INVX1 G50217 (.I(W32796), .ZN(O8397));
  INVX1 G50218 (.I(W6217), .ZN(W14348));
  INVX1 G50219 (.I(W25055), .ZN(O8433));
  INVX1 G50220 (.I(W10152), .ZN(W14338));
  INVX1 G50221 (.I(I123), .ZN(W14339));
  INVX1 G50222 (.I(W26497), .ZN(W36493));
  INVX1 G50223 (.I(W2975), .ZN(W14340));
  INVX1 G50224 (.I(W20946), .ZN(O8429));
  INVX1 G50225 (.I(W21296), .ZN(O8428));
  INVX1 G50226 (.I(W33461), .ZN(O8427));
  INVX1 G50227 (.I(I1239), .ZN(W14344));
  INVX1 G50228 (.I(W29921), .ZN(O8396));
  INVX1 G50229 (.I(W6270), .ZN(W14349));
  INVX1 G50230 (.I(W30402), .ZN(O8423));
  INVX1 G50231 (.I(W26981), .ZN(O8422));
  INVX1 G50232 (.I(W23219), .ZN(O8420));
  INVX1 G50233 (.I(W2663), .ZN(O856));
  INVX1 G50234 (.I(W18993), .ZN(O8418));
  INVX1 G50235 (.I(W26301), .ZN(O8417));
  INVX1 G50236 (.I(W7801), .ZN(W14357));
  INVX1 G50237 (.I(W34657), .ZN(O8415));
  INVX1 G50238 (.I(W21200), .ZN(O8367));
  INVX1 G50239 (.I(W25940), .ZN(O8381));
  INVX1 G50240 (.I(W9590), .ZN(W14410));
  INVX1 G50241 (.I(W12758), .ZN(O8377));
  INVX1 G50242 (.I(W2575), .ZN(W14412));
  INVX1 G50243 (.I(W8315), .ZN(W14415));
  INVX1 G50244 (.I(W35089), .ZN(W36402));
  INVX1 G50245 (.I(W6645), .ZN(W36400));
  INVX1 G50246 (.I(W5738), .ZN(O8373));
  INVX1 G50247 (.I(W13021), .ZN(O8368));
  INVX1 G50248 (.I(I1597), .ZN(W14406));
  INVX1 G50249 (.I(W17624), .ZN(W36388));
  INVX1 G50250 (.I(W1615), .ZN(W36386));
  INVX1 G50251 (.I(W13608), .ZN(O8362));
  INVX1 G50252 (.I(W3422), .ZN(O870));
  INVX1 G50253 (.I(W31951), .ZN(W36378));
  INVX1 G50254 (.I(W803), .ZN(O871));
  INVX1 G50255 (.I(W8071), .ZN(W14442));
  INVX1 G50256 (.I(W21074), .ZN(O8357));
  INVX1 G50257 (.I(W36229), .ZN(O8356));
  INVX1 G50258 (.I(W27483), .ZN(O8388));
  INVX1 G50259 (.I(W5811), .ZN(O863));
  INVX1 G50260 (.I(W7066), .ZN(W14387));
  INVX1 G50261 (.I(W11568), .ZN(W14388));
  INVX1 G50262 (.I(W21406), .ZN(W36432));
  INVX1 G50263 (.I(W34450), .ZN(O8392));
  INVX1 G50264 (.I(W13437), .ZN(W14391));
  INVX1 G50265 (.I(W11979), .ZN(W36427));
  INVX1 G50266 (.I(W12793), .ZN(W14394));
  INVX1 G50267 (.I(W256), .ZN(W36424));
  INVX1 G50268 (.I(W25437), .ZN(O8434));
  INVX1 G50269 (.I(W17053), .ZN(O8386));
  INVX1 G50270 (.I(W7666), .ZN(W14397));
  INVX1 G50271 (.I(W547), .ZN(W14398));
  INVX1 G50272 (.I(W762), .ZN(W14400));
  INVX1 G50273 (.I(W11834), .ZN(W14401));
  INVX1 G50274 (.I(W386), .ZN(O8383));
  INVX1 G50275 (.I(W16264), .ZN(W36415));
  INVX1 G50276 (.I(W17320), .ZN(O8382));
  INVX1 G50277 (.I(W13046), .ZN(W14405));
  INVX1 G50278 (.I(W13058), .ZN(W14250));
  INVX1 G50279 (.I(I147), .ZN(W14238));
  INVX1 G50280 (.I(W11809), .ZN(W14240));
  INVX1 G50281 (.I(W3441), .ZN(W14241));
  INVX1 G50282 (.I(W12320), .ZN(W36584));
  INVX1 G50283 (.I(I1159), .ZN(W14245));
  INVX1 G50284 (.I(W26221), .ZN(O8486));
  INVX1 G50285 (.I(W33571), .ZN(W36578));
  INVX1 G50286 (.I(W7645), .ZN(W14248));
  INVX1 G50287 (.I(W20596), .ZN(O8485));
  INVX1 G50288 (.I(W4182), .ZN(W14237));
  INVX1 G50289 (.I(W12088), .ZN(W14252));
  INVX1 G50290 (.I(W6710), .ZN(W14255));
  INVX1 G50291 (.I(W14196), .ZN(O8480));
  INVX1 G50292 (.I(W9724), .ZN(W14260));
  INVX1 G50293 (.I(W445), .ZN(W14262));
  INVX1 G50294 (.I(W33721), .ZN(O8473));
  INVX1 G50295 (.I(W4288), .ZN(O8471));
  INVX1 G50296 (.I(W6925), .ZN(W14266));
  INVX1 G50297 (.I(I224), .ZN(W36557));
  INVX1 G50298 (.I(W3619), .ZN(W14223));
  INVX1 G50299 (.I(W6844), .ZN(O8505));
  INVX1 G50300 (.I(W14172), .ZN(W36618));
  INVX1 G50301 (.I(W839), .ZN(W14209));
  INVX1 G50302 (.I(W6526), .ZN(W36616));
  INVX1 G50303 (.I(W24702), .ZN(W36615));
  INVX1 G50304 (.I(W8491), .ZN(W14211));
  INVX1 G50305 (.I(W1312), .ZN(W14218));
  INVX1 G50306 (.I(W20883), .ZN(W36610));
  INVX1 G50307 (.I(W24467), .ZN(O8498));
  INVX1 G50308 (.I(W13718), .ZN(W14267));
  INVX1 G50309 (.I(W21110), .ZN(O8497));
  INVX1 G50310 (.I(W2906), .ZN(O8496));
  INVX1 G50311 (.I(W5063), .ZN(O844));
  INVX1 G50312 (.I(W13327), .ZN(W14228));
  INVX1 G50313 (.I(W9726), .ZN(W14229));
  INVX1 G50314 (.I(W27205), .ZN(O8492));
  INVX1 G50315 (.I(W5618), .ZN(W14233));
  INVX1 G50316 (.I(W2038), .ZN(W14236));
  INVX1 G50317 (.I(W16036), .ZN(O8490));
  INVX1 G50318 (.I(W9975), .ZN(O8441));
  INVX1 G50319 (.I(W6947), .ZN(W14301));
  INVX1 G50320 (.I(W21051), .ZN(O8448));
  INVX1 G50321 (.I(W3396), .ZN(O8447));
  INVX1 G50322 (.I(W11143), .ZN(O8445));
  INVX1 G50323 (.I(W13275), .ZN(W14303));
  INVX1 G50324 (.I(W24940), .ZN(W36517));
  INVX1 G50325 (.I(W10107), .ZN(W14310));
  INVX1 G50326 (.I(W13204), .ZN(O854));
  INVX1 G50327 (.I(W8589), .ZN(W14312));
  INVX1 G50328 (.I(W23976), .ZN(O8451));
  INVX1 G50329 (.I(I1378), .ZN(W14315));
  INVX1 G50330 (.I(W2768), .ZN(O8439));
  INVX1 G50331 (.I(W8025), .ZN(W14327));
  INVX1 G50332 (.I(W9800), .ZN(W14331));
  INVX1 G50333 (.I(W1494), .ZN(W14332));
  INVX1 G50334 (.I(W6938), .ZN(W36503));
  INVX1 G50335 (.I(W480), .ZN(W14333));
  INVX1 G50336 (.I(W5867), .ZN(W14337));
  INVX1 G50337 (.I(W32400), .ZN(O8435));
  INVX1 G50338 (.I(W20108), .ZN(W36541));
  INVX1 G50339 (.I(W2634), .ZN(W36555));
  INVX1 G50340 (.I(W8593), .ZN(O8468));
  INVX1 G50341 (.I(W1914), .ZN(O8467));
  INVX1 G50342 (.I(W623), .ZN(O8465));
  INVX1 G50343 (.I(W7680), .ZN(W14274));
  INVX1 G50344 (.I(W702), .ZN(W14277));
  INVX1 G50345 (.I(W11614), .ZN(W14278));
  INVX1 G50346 (.I(W11869), .ZN(W14280));
  INVX1 G50347 (.I(W12125), .ZN(O850));
  INVX1 G50348 (.I(W16839), .ZN(O8067));
  INVX1 G50349 (.I(W32707), .ZN(W36540));
  INVX1 G50350 (.I(W431), .ZN(W14285));
  INVX1 G50351 (.I(I494), .ZN(O852));
  INVX1 G50352 (.I(W13033), .ZN(W14296));
  INVX1 G50353 (.I(W11474), .ZN(W36532));
  INVX1 G50354 (.I(W33172), .ZN(O8455));
  INVX1 G50355 (.I(W1663), .ZN(W36529));
  INVX1 G50356 (.I(W6438), .ZN(W14298));
  INVX1 G50357 (.I(W28470), .ZN(O8452));
  INVX1 G50358 (.I(W612), .ZN(O1032));
  INVX1 G50359 (.I(W9698), .ZN(W15568));
  INVX1 G50360 (.I(W9450), .ZN(O7690));
  INVX1 G50361 (.I(W30039), .ZN(O7689));
  INVX1 G50362 (.I(W27611), .ZN(O7688));
  INVX1 G50363 (.I(W6807), .ZN(W15570));
  INVX1 G50364 (.I(W29376), .ZN(W35233));
  INVX1 G50365 (.I(W18108), .ZN(O7687));
  INVX1 G50366 (.I(W12828), .ZN(W15576));
  INVX1 G50367 (.I(I982), .ZN(W15577));
  INVX1 G50368 (.I(W5490), .ZN(W35229));
  INVX1 G50369 (.I(W24343), .ZN(O7694));
  INVX1 G50370 (.I(W2753), .ZN(W35227));
  INVX1 G50371 (.I(W13616), .ZN(W15583));
  INVX1 G50372 (.I(W9779), .ZN(W15587));
  INVX1 G50373 (.I(W9891), .ZN(O7683));
  INVX1 G50374 (.I(W27049), .ZN(W35220));
  INVX1 G50375 (.I(W9960), .ZN(W35219));
  INVX1 G50376 (.I(W872), .ZN(W15592));
  INVX1 G50377 (.I(W25070), .ZN(W35216));
  INVX1 G50378 (.I(W8056), .ZN(W15594));
  INVX1 G50379 (.I(W4248), .ZN(W15548));
  INVX1 G50380 (.I(W32343), .ZN(W35284));
  INVX1 G50381 (.I(W3952), .ZN(W15525));
  INVX1 G50382 (.I(W4037), .ZN(O1023));
  INVX1 G50383 (.I(W8491), .ZN(W15531));
  INVX1 G50384 (.I(W29493), .ZN(W35277));
  INVX1 G50385 (.I(W12106), .ZN(W15540));
  INVX1 G50386 (.I(W11238), .ZN(W35269));
  INVX1 G50387 (.I(W3049), .ZN(W15543));
  INVX1 G50388 (.I(W4904), .ZN(W15546));
  INVX1 G50389 (.I(W841), .ZN(W15595));
  INVX1 G50390 (.I(W16460), .ZN(O7703));
  INVX1 G50391 (.I(W1), .ZN(W15550));
  INVX1 G50392 (.I(W1275), .ZN(W15555));
  INVX1 G50393 (.I(W7759), .ZN(W15557));
  INVX1 G50394 (.I(W2256), .ZN(W15558));
  INVX1 G50395 (.I(W26160), .ZN(O7696));
  INVX1 G50396 (.I(W3444), .ZN(W35252));
  INVX1 G50397 (.I(W1234), .ZN(W15562));
  INVX1 G50398 (.I(W22963), .ZN(W35248));
  INVX1 G50399 (.I(W15130), .ZN(W15654));
  INVX1 G50400 (.I(W30336), .ZN(O7659));
  INVX1 G50401 (.I(W12822), .ZN(W15647));
  INVX1 G50402 (.I(W28513), .ZN(W35167));
  INVX1 G50403 (.I(W14665), .ZN(O1043));
  INVX1 G50404 (.I(W11138), .ZN(W15649));
  INVX1 G50405 (.I(W13296), .ZN(W15651));
  INVX1 G50406 (.I(W12432), .ZN(O7654));
  INVX1 G50407 (.I(W23585), .ZN(O7653));
  INVX1 G50408 (.I(W34909), .ZN(O7652));
  INVX1 G50409 (.I(W21161), .ZN(O7661));
  INVX1 G50410 (.I(W9365), .ZN(W15655));
  INVX1 G50411 (.I(W5891), .ZN(O1045));
  INVX1 G50412 (.I(W7119), .ZN(W15662));
  INVX1 G50413 (.I(W11842), .ZN(W35152));
  INVX1 G50414 (.I(W5865), .ZN(O7648));
  INVX1 G50415 (.I(W3027), .ZN(W35150));
  INVX1 G50416 (.I(W1270), .ZN(O1048));
  INVX1 G50417 (.I(W7204), .ZN(W15667));
  INVX1 G50418 (.I(W2503), .ZN(W15668));
  INVX1 G50419 (.I(W8219), .ZN(W35190));
  INVX1 G50420 (.I(W15324), .ZN(W35210));
  INVX1 G50421 (.I(W8976), .ZN(W15604));
  INVX1 G50422 (.I(W18699), .ZN(W35207));
  INVX1 G50423 (.I(I319), .ZN(O1037));
  INVX1 G50424 (.I(W14118), .ZN(W15616));
  INVX1 G50425 (.I(W5516), .ZN(O1039));
  INVX1 G50426 (.I(W8136), .ZN(O7673));
  INVX1 G50427 (.I(W29559), .ZN(W35195));
  INVX1 G50428 (.I(W6929), .ZN(O7672));
  INVX1 G50429 (.I(W9309), .ZN(O7714));
  INVX1 G50430 (.I(W14242), .ZN(W15631));
  INVX1 G50431 (.I(W13374), .ZN(W15636));
  INVX1 G50432 (.I(W6704), .ZN(W15637));
  INVX1 G50433 (.I(W2386), .ZN(W35181));
  INVX1 G50434 (.I(W31580), .ZN(O7663));
  INVX1 G50435 (.I(W7795), .ZN(W15640));
  INVX1 G50436 (.I(W625), .ZN(W35176));
  INVX1 G50437 (.I(W7023), .ZN(O1042));
  INVX1 G50438 (.I(W14778), .ZN(W15645));
  INVX1 G50439 (.I(W8704), .ZN(W15429));
  INVX1 G50440 (.I(W29595), .ZN(W35375));
  INVX1 G50441 (.I(W19028), .ZN(W35374));
  INVX1 G50442 (.I(W52), .ZN(W15414));
  INVX1 G50443 (.I(W10329), .ZN(O7767));
  INVX1 G50444 (.I(W12012), .ZN(W15417));
  INVX1 G50445 (.I(W5831), .ZN(O1002));
  INVX1 G50446 (.I(W14313), .ZN(W15422));
  INVX1 G50447 (.I(W5681), .ZN(W15424));
  INVX1 G50448 (.I(W12983), .ZN(W15425));
  INVX1 G50449 (.I(W19826), .ZN(W35376));
  INVX1 G50450 (.I(W888), .ZN(W15433));
  INVX1 G50451 (.I(W1590), .ZN(O7758));
  INVX1 G50452 (.I(W10794), .ZN(W35356));
  INVX1 G50453 (.I(W1486), .ZN(W35355));
  INVX1 G50454 (.I(W7885), .ZN(W15439));
  INVX1 G50455 (.I(I1447), .ZN(W35353));
  INVX1 G50456 (.I(W15135), .ZN(W35352));
  INVX1 G50457 (.I(W20073), .ZN(O7757));
  INVX1 G50458 (.I(W17985), .ZN(O7755));
  INVX1 G50459 (.I(I1133), .ZN(W35387));
  INVX1 G50460 (.I(W14212), .ZN(O7786));
  INVX1 G50461 (.I(W6896), .ZN(O7785));
  INVX1 G50462 (.I(W5147), .ZN(O7784));
  INVX1 G50463 (.I(W5180), .ZN(W15399));
  INVX1 G50464 (.I(W12547), .ZN(W15400));
  INVX1 G50465 (.I(W5504), .ZN(O7779));
  INVX1 G50466 (.I(W18618), .ZN(W35395));
  INVX1 G50467 (.I(W18152), .ZN(O7775));
  INVX1 G50468 (.I(W14135), .ZN(O7773));
  INVX1 G50469 (.I(W1440), .ZN(W15445));
  INVX1 G50470 (.I(W290), .ZN(W15411));
  INVX1 G50471 (.I(W31097), .ZN(O7772));
  INVX1 G50472 (.I(W32470), .ZN(W35384));
  INVX1 G50473 (.I(W22532), .ZN(O7771));
  INVX1 G50474 (.I(W34803), .ZN(W35382));
  INVX1 G50475 (.I(W10423), .ZN(O7770));
  INVX1 G50476 (.I(W12532), .ZN(O7769));
  INVX1 G50477 (.I(W14855), .ZN(O7768));
  INVX1 G50478 (.I(W9229), .ZN(W35377));
  INVX1 G50479 (.I(W9732), .ZN(W35306));
  INVX1 G50480 (.I(W8870), .ZN(O7734));
  INVX1 G50481 (.I(W17976), .ZN(O7732));
  INVX1 G50482 (.I(W8424), .ZN(O7731));
  INVX1 G50483 (.I(W5075), .ZN(W35313));
  INVX1 G50484 (.I(W1750), .ZN(W35311));
  INVX1 G50485 (.I(W2690), .ZN(W35310));
  INVX1 G50486 (.I(W2920), .ZN(W15490));
  INVX1 G50487 (.I(I1366), .ZN(W15491));
  INVX1 G50488 (.I(W6140), .ZN(W15493));
  INVX1 G50489 (.I(W4527), .ZN(W15483));
  INVX1 G50490 (.I(W2212), .ZN(W35303));
  INVX1 G50491 (.I(W3469), .ZN(W15500));
  INVX1 G50492 (.I(W3554), .ZN(W15502));
  INVX1 G50493 (.I(W1377), .ZN(W15505));
  INVX1 G50494 (.I(I713), .ZN(W15509));
  INVX1 G50495 (.I(W51), .ZN(O1020));
  INVX1 G50496 (.I(W425), .ZN(W15520));
  INVX1 G50497 (.I(W12323), .ZN(W15521));
  INVX1 G50498 (.I(W6807), .ZN(O7715));
  INVX1 G50499 (.I(W12143), .ZN(W15470));
  INVX1 G50500 (.I(W8738), .ZN(W15449));
  INVX1 G50501 (.I(W679), .ZN(W15450));
  INVX1 G50502 (.I(W1515), .ZN(W15451));
  INVX1 G50503 (.I(W973), .ZN(W15453));
  INVX1 G50504 (.I(W8422), .ZN(W35341));
  INVX1 G50505 (.I(W14153), .ZN(W15454));
  INVX1 G50506 (.I(W3017), .ZN(O1009));
  INVX1 G50507 (.I(W271), .ZN(O1010));
  INVX1 G50508 (.I(W10359), .ZN(O7744));
  INVX1 G50509 (.I(W12300), .ZN(W15670));
  INVX1 G50510 (.I(I1497), .ZN(O1014));
  INVX1 G50511 (.I(W32444), .ZN(W35329));
  INVX1 G50512 (.I(W3624), .ZN(W15473));
  INVX1 G50513 (.I(W11321), .ZN(O1015));
  INVX1 G50514 (.I(W16217), .ZN(W35326));
  INVX1 G50515 (.I(W3799), .ZN(W15481));
  INVX1 G50516 (.I(I424), .ZN(W15482));
  INVX1 G50517 (.I(W3286), .ZN(W35321));
  INVX1 G50518 (.I(W10310), .ZN(O7736));
  INVX1 G50519 (.I(W5698), .ZN(O1079));
  INVX1 G50520 (.I(W16018), .ZN(O7549));
  INVX1 G50521 (.I(I481), .ZN(O7548));
  INVX1 G50522 (.I(W8696), .ZN(W34977));
  INVX1 G50523 (.I(W12391), .ZN(W34976));
  INVX1 G50524 (.I(I510), .ZN(O1076));
  INVX1 G50525 (.I(W1486), .ZN(W15851));
  INVX1 G50526 (.I(W7141), .ZN(W34972));
  INVX1 G50527 (.I(W24971), .ZN(W34971));
  INVX1 G50528 (.I(W6401), .ZN(W15852));
  INVX1 G50529 (.I(W5942), .ZN(W15859));
  INVX1 G50530 (.I(W7277), .ZN(W15844));
  INVX1 G50531 (.I(W34232), .ZN(W34959));
  INVX1 G50532 (.I(W18470), .ZN(O7536));
  INVX1 G50533 (.I(W14539), .ZN(W15878));
  INVX1 G50534 (.I(W4039), .ZN(W15880));
  INVX1 G50535 (.I(W4422), .ZN(W15881));
  INVX1 G50536 (.I(W9265), .ZN(W34946));
  INVX1 G50537 (.I(W10351), .ZN(O1085));
  INVX1 G50538 (.I(W11920), .ZN(W15893));
  INVX1 G50539 (.I(W33200), .ZN(O7528));
  INVX1 G50540 (.I(W19738), .ZN(W34997));
  INVX1 G50541 (.I(W31179), .ZN(O7571));
  INVX1 G50542 (.I(W18310), .ZN(O7570));
  INVX1 G50543 (.I(W11654), .ZN(O7569));
  INVX1 G50544 (.I(W4347), .ZN(W15814));
  INVX1 G50545 (.I(W11186), .ZN(O1070));
  INVX1 G50546 (.I(W716), .ZN(W15817));
  INVX1 G50547 (.I(W9989), .ZN(W15819));
  INVX1 G50548 (.I(W10586), .ZN(W15822));
  INVX1 G50549 (.I(W2757), .ZN(W15823));
  INVX1 G50550 (.I(W1817), .ZN(W15896));
  INVX1 G50551 (.I(W30152), .ZN(W34995));
  INVX1 G50552 (.I(W20651), .ZN(W34993));
  INVX1 G50553 (.I(W6117), .ZN(W15832));
  INVX1 G50554 (.I(W7821), .ZN(O7558));
  INVX1 G50555 (.I(W9926), .ZN(O7557));
  INVX1 G50556 (.I(W15454), .ZN(O7556));
  INVX1 G50557 (.I(W6463), .ZN(W15833));
  INVX1 G50558 (.I(W34579), .ZN(W34986));
  INVX1 G50559 (.I(W5296), .ZN(O1072));
  INVX1 G50560 (.I(W32928), .ZN(W34897));
  INVX1 G50561 (.I(W8954), .ZN(W15926));
  INVX1 G50562 (.I(W22187), .ZN(O7508));
  INVX1 G50563 (.I(W5280), .ZN(W34905));
  INVX1 G50564 (.I(W8702), .ZN(W15931));
  INVX1 G50565 (.I(W23219), .ZN(O7503));
  INVX1 G50566 (.I(W33352), .ZN(O7502));
  INVX1 G50567 (.I(W9930), .ZN(W34900));
  INVX1 G50568 (.I(W190), .ZN(W15933));
  INVX1 G50569 (.I(W59), .ZN(W15935));
  INVX1 G50570 (.I(W4948), .ZN(O7509));
  INVX1 G50571 (.I(W28794), .ZN(O7500));
  INVX1 G50572 (.I(I442), .ZN(W15937));
  INVX1 G50573 (.I(W11285), .ZN(W15939));
  INVX1 G50574 (.I(W4172), .ZN(W15940));
  INVX1 G50575 (.I(W5762), .ZN(W15941));
  INVX1 G50576 (.I(W12744), .ZN(W34891));
  INVX1 G50577 (.I(W8600), .ZN(W15942));
  INVX1 G50578 (.I(W2917), .ZN(W15944));
  INVX1 G50579 (.I(I1811), .ZN(O7496));
  INVX1 G50580 (.I(W8947), .ZN(W15908));
  INVX1 G50581 (.I(W5142), .ZN(W15899));
  INVX1 G50582 (.I(W32845), .ZN(W34935));
  INVX1 G50583 (.I(W13372), .ZN(O1088));
  INVX1 G50584 (.I(W8364), .ZN(W15904));
  INVX1 G50585 (.I(I1370), .ZN(W15905));
  INVX1 G50586 (.I(W30756), .ZN(W34930));
  INVX1 G50587 (.I(W4948), .ZN(W15906));
  INVX1 G50588 (.I(W12370), .ZN(O7522));
  INVX1 G50589 (.I(W24322), .ZN(O7521));
  INVX1 G50590 (.I(W32323), .ZN(O7572));
  INVX1 G50591 (.I(W31343), .ZN(O7518));
  INVX1 G50592 (.I(W21957), .ZN(O7516));
  INVX1 G50593 (.I(W3967), .ZN(W15911));
  INVX1 G50594 (.I(I1308), .ZN(W15913));
  INVX1 G50595 (.I(W8588), .ZN(W15915));
  INVX1 G50596 (.I(W3731), .ZN(W15921));
  INVX1 G50597 (.I(W2654), .ZN(O7510));
  INVX1 G50598 (.I(W8400), .ZN(W15925));
  INVX1 G50599 (.I(W16659), .ZN(W34911));
  INVX1 G50600 (.I(W3887), .ZN(W15724));
  INVX1 G50601 (.I(W12877), .ZN(W15712));
  INVX1 G50602 (.I(W14992), .ZN(W35107));
  INVX1 G50603 (.I(W4126), .ZN(W15715));
  INVX1 G50604 (.I(I1715), .ZN(W15716));
  INVX1 G50605 (.I(W30733), .ZN(O7625));
  INVX1 G50606 (.I(W16156), .ZN(O7624));
  INVX1 G50607 (.I(W7803), .ZN(W15720));
  INVX1 G50608 (.I(W28613), .ZN(O7622));
  INVX1 G50609 (.I(W6998), .ZN(W15722));
  INVX1 G50610 (.I(W9816), .ZN(W35111));
  INVX1 G50611 (.I(W2955), .ZN(W15725));
  INVX1 G50612 (.I(W14186), .ZN(W15729));
  INVX1 G50613 (.I(W964), .ZN(W15733));
  INVX1 G50614 (.I(W12391), .ZN(W15735));
  INVX1 G50615 (.I(W7445), .ZN(W15736));
  INVX1 G50616 (.I(W5937), .ZN(W15741));
  INVX1 G50617 (.I(W1582), .ZN(O1059));
  INVX1 G50618 (.I(W14235), .ZN(W15747));
  INVX1 G50619 (.I(W33006), .ZN(O7611));
  INVX1 G50620 (.I(W3218), .ZN(W35126));
  INVX1 G50621 (.I(W11831), .ZN(W15671));
  INVX1 G50622 (.I(W13097), .ZN(W35142));
  INVX1 G50623 (.I(W15074), .ZN(W15672));
  INVX1 G50624 (.I(W5446), .ZN(O1050));
  INVX1 G50625 (.I(W3276), .ZN(W15678));
  INVX1 G50626 (.I(I514), .ZN(W15679));
  INVX1 G50627 (.I(W14518), .ZN(W15683));
  INVX1 G50628 (.I(I969), .ZN(W15688));
  INVX1 G50629 (.I(W7904), .ZN(W15690));
  INVX1 G50630 (.I(W29195), .ZN(O7610));
  INVX1 G50631 (.I(W679), .ZN(W15694));
  INVX1 G50632 (.I(I792), .ZN(O1052));
  INVX1 G50633 (.I(W15527), .ZN(W15696));
  INVX1 G50634 (.I(W26254), .ZN(O7637));
  INVX1 G50635 (.I(W11299), .ZN(O7636));
  INVX1 G50636 (.I(W13781), .ZN(W15697));
  INVX1 G50637 (.I(W1871), .ZN(W15700));
  INVX1 G50638 (.I(W9215), .ZN(W15705));
  INVX1 G50639 (.I(W23363), .ZN(O7632));
  INVX1 G50640 (.I(W25651), .ZN(O7583));
  INVX1 G50641 (.I(W678), .ZN(W35040));
  INVX1 G50642 (.I(W11797), .ZN(W15783));
  INVX1 G50643 (.I(W11345), .ZN(W15784));
  INVX1 G50644 (.I(W31953), .ZN(W35037));
  INVX1 G50645 (.I(W14316), .ZN(W35036));
  INVX1 G50646 (.I(W12511), .ZN(O1067));
  INVX1 G50647 (.I(W7513), .ZN(O1068));
  INVX1 G50648 (.I(W3947), .ZN(W15789));
  INVX1 G50649 (.I(W11051), .ZN(W15792));
  INVX1 G50650 (.I(W14904), .ZN(W15781));
  INVX1 G50651 (.I(I1942), .ZN(W15796));
  INVX1 G50652 (.I(W11191), .ZN(W35027));
  INVX1 G50653 (.I(W32595), .ZN(O7582));
  INVX1 G50654 (.I(W29776), .ZN(W35023));
  INVX1 G50655 (.I(W24558), .ZN(W35022));
  INVX1 G50656 (.I(W24326), .ZN(W35021));
  INVX1 G50657 (.I(W12222), .ZN(W15803));
  INVX1 G50658 (.I(W14238), .ZN(O1069));
  INVX1 G50659 (.I(W5681), .ZN(W15812));
  INVX1 G50660 (.I(W22359), .ZN(O7598));
  INVX1 G50661 (.I(W26022), .ZN(O7609));
  INVX1 G50662 (.I(W33968), .ZN(O7608));
  INVX1 G50663 (.I(W15462), .ZN(W35072));
  INVX1 G50664 (.I(I1812), .ZN(W15752));
  INVX1 G50665 (.I(W11146), .ZN(W15754));
  INVX1 G50666 (.I(I1277), .ZN(O7605));
  INVX1 G50667 (.I(W8796), .ZN(W15759));
  INVX1 G50668 (.I(W5016), .ZN(W15761));
  INVX1 G50669 (.I(W13444), .ZN(W15768));
  INVX1 G50670 (.I(W5099), .ZN(W15392));
  INVX1 G50671 (.I(I1775), .ZN(W15769));
  INVX1 G50672 (.I(W19935), .ZN(O7596));
  INVX1 G50673 (.I(W14033), .ZN(W15771));
  INVX1 G50674 (.I(W25767), .ZN(O7595));
  INVX1 G50675 (.I(W13336), .ZN(O1065));
  INVX1 G50676 (.I(W14810), .ZN(W15777));
  INVX1 G50677 (.I(W10560), .ZN(O7591));
  INVX1 G50678 (.I(W28646), .ZN(W35045));
  INVX1 G50679 (.I(W19069), .ZN(W35043));
  INVX1 G50680 (.I(W20249), .ZN(W35726));
  INVX1 G50681 (.I(W1677), .ZN(W15058));
  INVX1 G50682 (.I(W6029), .ZN(W15059));
  INVX1 G50683 (.I(W25192), .ZN(O7984));
  INVX1 G50684 (.I(W939), .ZN(W15063));
  INVX1 G50685 (.I(W12260), .ZN(W15064));
  INVX1 G50686 (.I(W5827), .ZN(O956));
  INVX1 G50687 (.I(W6244), .ZN(W15066));
  INVX1 G50688 (.I(I1554), .ZN(W15067));
  INVX1 G50689 (.I(W7619), .ZN(O957));
  INVX1 G50690 (.I(W3334), .ZN(W35727));
  INVX1 G50691 (.I(W15613), .ZN(O7987));
  INVX1 G50692 (.I(I578), .ZN(O7981));
  INVX1 G50693 (.I(W8229), .ZN(W15073));
  INVX1 G50694 (.I(W28013), .ZN(W35722));
  INVX1 G50695 (.I(W12297), .ZN(W15074));
  INVX1 G50696 (.I(W6690), .ZN(W15075));
  INVX1 G50697 (.I(I242), .ZN(W15077));
  INVX1 G50698 (.I(W10483), .ZN(O7975));
  INVX1 G50699 (.I(W7336), .ZN(W15081));
  INVX1 G50700 (.I(W6545), .ZN(W15084));
  INVX1 G50701 (.I(W13840), .ZN(W15035));
  INVX1 G50702 (.I(W14321), .ZN(O8002));
  INVX1 G50703 (.I(W11531), .ZN(W15025));
  INVX1 G50704 (.I(W6863), .ZN(W35762));
  INVX1 G50705 (.I(W4124), .ZN(W15026));
  INVX1 G50706 (.I(W5993), .ZN(O947));
  INVX1 G50707 (.I(W7079), .ZN(O948));
  INVX1 G50708 (.I(W14729), .ZN(W15031));
  INVX1 G50709 (.I(W3950), .ZN(W15032));
  INVX1 G50710 (.I(W5327), .ZN(O949));
  INVX1 G50711 (.I(W33448), .ZN(O7972));
  INVX1 G50712 (.I(W701), .ZN(W15038));
  INVX1 G50713 (.I(W11852), .ZN(O7996));
  INVX1 G50714 (.I(W16781), .ZN(O7995));
  INVX1 G50715 (.I(W14274), .ZN(O951));
  INVX1 G50716 (.I(W15028), .ZN(O952));
  INVX1 G50717 (.I(W14538), .ZN(W15047));
  INVX1 G50718 (.I(I1896), .ZN(O7990));
  INVX1 G50719 (.I(W19906), .ZN(O7989));
  INVX1 G50720 (.I(W396), .ZN(W15055));
  INVX1 G50721 (.I(W3870), .ZN(O7948));
  INVX1 G50722 (.I(W10944), .ZN(W35677));
  INVX1 G50723 (.I(W19895), .ZN(O7956));
  INVX1 G50724 (.I(I832), .ZN(W15132));
  INVX1 G50725 (.I(W12527), .ZN(W15135));
  INVX1 G50726 (.I(W5300), .ZN(W15136));
  INVX1 G50727 (.I(W4534), .ZN(W15140));
  INVX1 G50728 (.I(W18866), .ZN(W35666));
  INVX1 G50729 (.I(W16631), .ZN(O7949));
  INVX1 G50730 (.I(W1902), .ZN(W15147));
  INVX1 G50731 (.I(W31371), .ZN(O7957));
  INVX1 G50732 (.I(W13600), .ZN(W15148));
  INVX1 G50733 (.I(W8675), .ZN(W15150));
  INVX1 G50734 (.I(W20515), .ZN(W35660));
  INVX1 G50735 (.I(W6327), .ZN(W15151));
  INVX1 G50736 (.I(I572), .ZN(W35658));
  INVX1 G50737 (.I(W20184), .ZN(O7946));
  INVX1 G50738 (.I(W32369), .ZN(O7943));
  INVX1 G50739 (.I(W11868), .ZN(O7942));
  INVX1 G50740 (.I(W1521), .ZN(W15156));
  INVX1 G50741 (.I(W11271), .ZN(O961));
  INVX1 G50742 (.I(W25797), .ZN(W35711));
  INVX1 G50743 (.I(W23154), .ZN(W35705));
  INVX1 G50744 (.I(W13899), .ZN(W35704));
  INVX1 G50745 (.I(W11566), .ZN(W15096));
  INVX1 G50746 (.I(W908), .ZN(W15099));
  INVX1 G50747 (.I(W7389), .ZN(W15100));
  INVX1 G50748 (.I(W33701), .ZN(O7968));
  INVX1 G50749 (.I(I1121), .ZN(O7967));
  INVX1 G50750 (.I(W267), .ZN(W15108));
  INVX1 G50751 (.I(W1866), .ZN(W35765));
  INVX1 G50752 (.I(W2119), .ZN(W15111));
  INVX1 G50753 (.I(W10345), .ZN(W15112));
  INVX1 G50754 (.I(W10132), .ZN(W35693));
  INVX1 G50755 (.I(W2099), .ZN(W15116));
  INVX1 G50756 (.I(W27637), .ZN(W35688));
  INVX1 G50757 (.I(W22377), .ZN(W35687));
  INVX1 G50758 (.I(W2361), .ZN(W15119));
  INVX1 G50759 (.I(W18447), .ZN(O7961));
  INVX1 G50760 (.I(W8478), .ZN(W15131));
  INVX1 G50761 (.I(W27180), .ZN(W35851));
  INVX1 G50762 (.I(W8981), .ZN(W14930));
  INVX1 G50763 (.I(W9830), .ZN(W14931));
  INVX1 G50764 (.I(W14549), .ZN(O8046));
  INVX1 G50765 (.I(W15792), .ZN(O8045));
  INVX1 G50766 (.I(W30791), .ZN(O8044));
  INVX1 G50767 (.I(W13235), .ZN(W35855));
  INVX1 G50768 (.I(W1277), .ZN(W14934));
  INVX1 G50769 (.I(W12861), .ZN(W14935));
  INVX1 G50770 (.I(W16266), .ZN(W35852));
  INVX1 G50771 (.I(W2736), .ZN(W14924));
  INVX1 G50772 (.I(W16335), .ZN(O8043));
  INVX1 G50773 (.I(W21599), .ZN(O8042));
  INVX1 G50774 (.I(I1571), .ZN(W14943));
  INVX1 G50775 (.I(W7164), .ZN(W14944));
  INVX1 G50776 (.I(W25235), .ZN(W35838));
  INVX1 G50777 (.I(W6816), .ZN(W35837));
  INVX1 G50778 (.I(W23405), .ZN(W35835));
  INVX1 G50779 (.I(W4901), .ZN(W14951));
  INVX1 G50780 (.I(W8244), .ZN(W14952));
  INVX1 G50781 (.I(W21520), .ZN(W35877));
  INVX1 G50782 (.I(W6007), .ZN(W14900));
  INVX1 G50783 (.I(W4359), .ZN(O8065));
  INVX1 G50784 (.I(I967), .ZN(W14901));
  INVX1 G50785 (.I(W19183), .ZN(O8061));
  INVX1 G50786 (.I(W32424), .ZN(W35884));
  INVX1 G50787 (.I(W32280), .ZN(O8060));
  INVX1 G50788 (.I(W5268), .ZN(W14905));
  INVX1 G50789 (.I(W13055), .ZN(O930));
  INVX1 G50790 (.I(W14300), .ZN(W14914));
  INVX1 G50791 (.I(W9254), .ZN(O936));
  INVX1 G50792 (.I(W6920), .ZN(W35876));
  INVX1 G50793 (.I(W28441), .ZN(W35874));
  INVX1 G50794 (.I(W2554), .ZN(O8057));
  INVX1 G50795 (.I(W16142), .ZN(O8056));
  INVX1 G50796 (.I(W3768), .ZN(W14918));
  INVX1 G50797 (.I(W34529), .ZN(O8055));
  INVX1 G50798 (.I(W7118), .ZN(W14919));
  INVX1 G50799 (.I(W5559), .ZN(W14922));
  INVX1 G50800 (.I(W26515), .ZN(O8051));
  INVX1 G50801 (.I(I408), .ZN(W15009));
  INVX1 G50802 (.I(W10390), .ZN(O942));
  INVX1 G50803 (.I(I1802), .ZN(O8018));
  INVX1 G50804 (.I(W25571), .ZN(W35793));
  INVX1 G50805 (.I(W15799), .ZN(O8016));
  INVX1 G50806 (.I(I1968), .ZN(W14997));
  INVX1 G50807 (.I(W25007), .ZN(W35787));
  INVX1 G50808 (.I(W8098), .ZN(W15000));
  INVX1 G50809 (.I(W17499), .ZN(O8009));
  INVX1 G50810 (.I(W9449), .ZN(W15008));
  INVX1 G50811 (.I(W5859), .ZN(W35798));
  INVX1 G50812 (.I(W6205), .ZN(W15011));
  INVX1 G50813 (.I(W14101), .ZN(W35778));
  INVX1 G50814 (.I(W12499), .ZN(W15012));
  INVX1 G50815 (.I(W28370), .ZN(W35776));
  INVX1 G50816 (.I(W18483), .ZN(O8006));
  INVX1 G50817 (.I(W12888), .ZN(W15013));
  INVX1 G50818 (.I(W6583), .ZN(W15022));
  INVX1 G50819 (.I(W12342), .ZN(W35767));
  INVX1 G50820 (.I(W15280), .ZN(O8003));
  INVX1 G50821 (.I(W10687), .ZN(O939));
  INVX1 G50822 (.I(W8523), .ZN(W14957));
  INVX1 G50823 (.I(W11506), .ZN(O8032));
  INVX1 G50824 (.I(W3776), .ZN(W14961));
  INVX1 G50825 (.I(W6251), .ZN(W14963));
  INVX1 G50826 (.I(W90), .ZN(W14964));
  INVX1 G50827 (.I(W14093), .ZN(W14965));
  INVX1 G50828 (.I(W3587), .ZN(O8029));
  INVX1 G50829 (.I(W26776), .ZN(W35817));
  INVX1 G50830 (.I(W10945), .ZN(O938));
  INVX1 G50831 (.I(W20288), .ZN(O7940));
  INVX1 G50832 (.I(W4112), .ZN(W14976));
  INVX1 G50833 (.I(W317), .ZN(W14977));
  INVX1 G50834 (.I(W33787), .ZN(W35808));
  INVX1 G50835 (.I(W13562), .ZN(W14978));
  INVX1 G50836 (.I(W14364), .ZN(W35805));
  INVX1 G50837 (.I(I1606), .ZN(W35804));
  INVX1 G50838 (.I(W10250), .ZN(W14983));
  INVX1 G50839 (.I(W3779), .ZN(W14987));
  INVX1 G50840 (.I(W423), .ZN(O941));
  INVX1 G50841 (.I(W4455), .ZN(O7829));
  INVX1 G50842 (.I(W1338), .ZN(W35493));
  INVX1 G50843 (.I(W24610), .ZN(O7836));
  INVX1 G50844 (.I(W16327), .ZN(W35491));
  INVX1 G50845 (.I(W8259), .ZN(O7835));
  INVX1 G50846 (.I(W28672), .ZN(W35489));
  INVX1 G50847 (.I(W23504), .ZN(O7834));
  INVX1 G50848 (.I(W12952), .ZN(W15305));
  INVX1 G50849 (.I(I1086), .ZN(W15307));
  INVX1 G50850 (.I(W6479), .ZN(W15314));
  INVX1 G50851 (.I(W34268), .ZN(O7830));
  INVX1 G50852 (.I(W27879), .ZN(O7837));
  INVX1 G50853 (.I(W7248), .ZN(O7828));
  INVX1 G50854 (.I(W3368), .ZN(O7827));
  INVX1 G50855 (.I(W8874), .ZN(W35478));
  INVX1 G50856 (.I(W2155), .ZN(W35477));
  INVX1 G50857 (.I(W270), .ZN(O7825));
  INVX1 G50858 (.I(W11065), .ZN(W15321));
  INVX1 G50859 (.I(W30899), .ZN(O7823));
  INVX1 G50860 (.I(W20107), .ZN(O7822));
  INVX1 G50861 (.I(W5617), .ZN(W15323));
  INVX1 G50862 (.I(W10439), .ZN(W15287));
  INVX1 G50863 (.I(W8850), .ZN(W15275));
  INVX1 G50864 (.I(W12744), .ZN(W15276));
  INVX1 G50865 (.I(W17628), .ZN(O7857));
  INVX1 G50866 (.I(W15237), .ZN(O7854));
  INVX1 G50867 (.I(W1956), .ZN(W15282));
  INVX1 G50868 (.I(W14111), .ZN(W15284));
  INVX1 G50869 (.I(W29208), .ZN(W35512));
  INVX1 G50870 (.I(W18154), .ZN(O7850));
  INVX1 G50871 (.I(W424), .ZN(W15285));
  INVX1 G50872 (.I(W9471), .ZN(O990));
  INVX1 G50873 (.I(W10851), .ZN(W15288));
  INVX1 G50874 (.I(W6064), .ZN(O985));
  INVX1 G50875 (.I(W6031), .ZN(W15291));
  INVX1 G50876 (.I(W2525), .ZN(O986));
  INVX1 G50877 (.I(W24286), .ZN(O7844));
  INVX1 G50878 (.I(W11589), .ZN(O987));
  INVX1 G50879 (.I(W9172), .ZN(W15296));
  INVX1 G50880 (.I(W205), .ZN(W15301));
  INVX1 G50881 (.I(W8078), .ZN(W15304));
  INVX1 G50882 (.I(W10979), .ZN(W15380));
  INVX1 G50883 (.I(W2764), .ZN(W15358));
  INVX1 G50884 (.I(I1471), .ZN(W15359));
  INVX1 G50885 (.I(W530), .ZN(W35435));
  INVX1 G50886 (.I(I1381), .ZN(O7801));
  INVX1 G50887 (.I(W1114), .ZN(O7799));
  INVX1 G50888 (.I(W3841), .ZN(W15372));
  INVX1 G50889 (.I(W34662), .ZN(W35423));
  INVX1 G50890 (.I(W2623), .ZN(W15377));
  INVX1 G50891 (.I(W14394), .ZN(W15378));
  INVX1 G50892 (.I(W9581), .ZN(W15357));
  INVX1 G50893 (.I(W17539), .ZN(W35419));
  INVX1 G50894 (.I(W19331), .ZN(O7796));
  INVX1 G50895 (.I(W7513), .ZN(O997));
  INVX1 G50896 (.I(W7234), .ZN(W15382));
  INVX1 G50897 (.I(I1786), .ZN(O999));
  INVX1 G50898 (.I(W7353), .ZN(W15390));
  INVX1 G50899 (.I(W19378), .ZN(W35409));
  INVX1 G50900 (.I(W1934), .ZN(O7789));
  INVX1 G50901 (.I(W21257), .ZN(O7788));
  INVX1 G50902 (.I(W31260), .ZN(W35452));
  INVX1 G50903 (.I(I595), .ZN(W15331));
  INVX1 G50904 (.I(W3244), .ZN(W15333));
  INVX1 G50905 (.I(W29711), .ZN(O7818));
  INVX1 G50906 (.I(W5266), .ZN(O7816));
  INVX1 G50907 (.I(W26204), .ZN(W35460));
  INVX1 G50908 (.I(W15211), .ZN(W15341));
  INVX1 G50909 (.I(W11146), .ZN(W15343));
  INVX1 G50910 (.I(W32943), .ZN(W35454));
  INVX1 G50911 (.I(W11874), .ZN(O995));
  INVX1 G50912 (.I(W12138), .ZN(W35523));
  INVX1 G50913 (.I(W12306), .ZN(W15347));
  INVX1 G50914 (.I(W18390), .ZN(W35448));
  INVX1 G50915 (.I(W3466), .ZN(W15348));
  INVX1 G50916 (.I(W537), .ZN(W15349));
  INVX1 G50917 (.I(W23809), .ZN(O7808));
  INVX1 G50918 (.I(W20543), .ZN(W35442));
  INVX1 G50919 (.I(W5477), .ZN(W15352));
  INVX1 G50920 (.I(W4032), .ZN(W15356));
  INVX1 G50921 (.I(W5222), .ZN(O7806));
  INVX1 G50922 (.I(I1136), .ZN(W35602));
  INVX1 G50923 (.I(I829), .ZN(W15192));
  INVX1 G50924 (.I(W25754), .ZN(O7916));
  INVX1 G50925 (.I(W3762), .ZN(W15197));
  INVX1 G50926 (.I(W8673), .ZN(W15198));
  INVX1 G50927 (.I(W5930), .ZN(O7913));
  INVX1 G50928 (.I(W13660), .ZN(O973));
  INVX1 G50929 (.I(W4), .ZN(O7910));
  INVX1 G50930 (.I(W29216), .ZN(W35604));
  INVX1 G50931 (.I(W15472), .ZN(O7909));
  INVX1 G50932 (.I(W12208), .ZN(W35617));
  INVX1 G50933 (.I(W3392), .ZN(W35600));
  INVX1 G50934 (.I(W1974), .ZN(W15205));
  INVX1 G50935 (.I(I832), .ZN(W15208));
  INVX1 G50936 (.I(W6556), .ZN(W15212));
  INVX1 G50937 (.I(W9782), .ZN(O974));
  INVX1 G50938 (.I(W35391), .ZN(O7903));
  INVX1 G50939 (.I(W15261), .ZN(O7902));
  INVX1 G50940 (.I(I1132), .ZN(W15217));
  INVX1 G50941 (.I(W9967), .ZN(O7899));
  INVX1 G50942 (.I(W9341), .ZN(W15183));
  INVX1 G50943 (.I(I364), .ZN(O7939));
  INVX1 G50944 (.I(W12171), .ZN(W15161));
  INVX1 G50945 (.I(W22682), .ZN(O7935));
  INVX1 G50946 (.I(W29751), .ZN(O7933));
  INVX1 G50947 (.I(W2416), .ZN(O7932));
  INVX1 G50948 (.I(W119), .ZN(O7930));
  INVX1 G50949 (.I(W6112), .ZN(W15173));
  INVX1 G50950 (.I(W8561), .ZN(W15177));
  INVX1 G50951 (.I(I1289), .ZN(W15181));
  INVX1 G50952 (.I(W34533), .ZN(O7898));
  INVX1 G50953 (.I(W19198), .ZN(O7926));
  INVX1 G50954 (.I(W30224), .ZN(W35625));
  INVX1 G50955 (.I(W11863), .ZN(W15187));
  INVX1 G50956 (.I(W18398), .ZN(W35623));
  INVX1 G50957 (.I(W27397), .ZN(O7925));
  INVX1 G50958 (.I(I1554), .ZN(W15190));
  INVX1 G50959 (.I(W25621), .ZN(W35620));
  INVX1 G50960 (.I(W21208), .ZN(O7923));
  INVX1 G50961 (.I(W818), .ZN(W15191));
  INVX1 G50962 (.I(W1282), .ZN(W15257));
  INVX1 G50963 (.I(W24961), .ZN(O7877));
  INVX1 G50964 (.I(W11335), .ZN(W15251));
  INVX1 G50965 (.I(W3817), .ZN(O980));
  INVX1 G50966 (.I(W29218), .ZN(W35549));
  INVX1 G50967 (.I(W29578), .ZN(W35548));
  INVX1 G50968 (.I(W8919), .ZN(O982));
  INVX1 G50969 (.I(W14722), .ZN(O7873));
  INVX1 G50970 (.I(W10942), .ZN(O7872));
  INVX1 G50971 (.I(W29989), .ZN(O7871));
  INVX1 G50972 (.I(W6133), .ZN(W15249));
  INVX1 G50973 (.I(I499), .ZN(W15258));
  INVX1 G50974 (.I(W10324), .ZN(W15260));
  INVX1 G50975 (.I(W713), .ZN(W15262));
  INVX1 G50976 (.I(W33590), .ZN(W35535));
  INVX1 G50977 (.I(W6987), .ZN(W15265));
  INVX1 G50978 (.I(W26721), .ZN(O7863));
  INVX1 G50979 (.I(W7920), .ZN(W15267));
  INVX1 G50980 (.I(W14688), .ZN(O7860));
  INVX1 G50981 (.I(W34501), .ZN(W35525));
  INVX1 G50982 (.I(W30687), .ZN(O7887));
  INVX1 G50983 (.I(W3004), .ZN(W15222));
  INVX1 G50984 (.I(W19052), .ZN(O7896));
  INVX1 G50985 (.I(W11847), .ZN(W15225));
  INVX1 G50986 (.I(W33006), .ZN(O7892));
  INVX1 G50987 (.I(I358), .ZN(W15229));
  INVX1 G50988 (.I(W13938), .ZN(O7889));
  INVX1 G50989 (.I(W14609), .ZN(W15234));
  INVX1 G50990 (.I(W4734), .ZN(W35571));
  INVX1 G50991 (.I(W11667), .ZN(W35570));
  INVX1 G50992 (.I(W37962), .ZN(O11075));
  INVX1 G50993 (.I(W11275), .ZN(O7886));
  INVX1 G50994 (.I(W3663), .ZN(W15235));
  INVX1 G50995 (.I(W3662), .ZN(W15236));
  INVX1 G50996 (.I(W11079), .ZN(W15237));
  INVX1 G50997 (.I(W4264), .ZN(W15240));
  INVX1 G50998 (.I(W6358), .ZN(W15245));
  INVX1 G50999 (.I(W9701), .ZN(O7880));
  INVX1 G51000 (.I(W18780), .ZN(O7879));
  INVX1 G51001 (.I(I732), .ZN(W15246));
endmodule
