module hidden_1 (I0, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I16, I17, I18, I19, I20, I21, I22, I23, I24, I26, I27, I28, I29, I30, I31, I32, I34, I36, I38, I39, I40, I42, I43, I44, I45, I46, I48, I49, I50, I51, I52, I54, I55, I56, I57, I58, I60, I61, I62, I64, I65, I66, I68, I70, I71, I72, I74, I75, I76, I78, I79, I80, I81, I82, I84, I85, I86, I88, I90, I91, I92, I94, I95, I96, I98, I100, I102, I103, I104, I106, I108, I109, I110, I111, I112, I113, I114, I115, I116, I117, I118, I120, I121, I122, I123, I124, I126, I128, I130, I132, I134, I135, I136, I137, I138, I140, I142, I144, I145, I146, I147, I148, I150, I151, I152, I153, I154, I156, I157, I158, I160, I161, I162, I163, I164, I165, I166, I168, I169, I170, I171, I172, I174, I175, I176, I178, I179, I180, I181, I182, I184, I185, I186, I188, I190, I191, I192, I193, I194, I195, I196, I197, I198, I200, I202, I203, I204, I206, I207, I208, I209, I210, I212, I213, I214, I215, I216, I217, I218, I219, I220, I221, I222, I223, I224, I225, I226, I227, I228, I229, I230, I231, I232, I233, I234, I235, I236, I237, I238, I239, I240, I241, I242, I243, I244, I245, I246, I247, I248, I249, I250, I252, I253, I254, I255, I256, I257, I258, I259, I260, I261, I262, I263, I264, I266, I267, I268, I269, I270, I271, I272, I274, I276, I277, I278, I280, I282, I283, I284, I285, I286, I288, I289, I290, I291, I292, I294, I296, I297, I298, I299, I300, I301, I302, I303, I304, I305, I306, I308, I309, I310, I312, I313, I314, I315, I316, I317, I318, I319, I320, I322, I323, I324, I326, I328, I329, I330, I331, I332, I334, I335, I336, I337, I338, I339, I340, I342, I344, I346, I347, I348, I349, I350, I351, I352, I353, I354, I355, I356, I357, I358, I360, I361, I362, I364, I365, I366, I368, I370, I371, I372, I374, I375, I376, I378, I380, I382, I384, I385, I386, I387, I388, I389, I390, I391, I392, I393, I394, I396, I398, I400, I401, I402, I404, I405, I406, I407, I408, I409, I410, I412, I413, I414, I415, I416, I417, I418, I420, I421, I422, I423, I424, I426, I428, I429, I430, I431, I432, I433, I434, I435, I436, I437, I438, I439, I440, I441, I442, I443, I444, I445, I446, I447, I448, I450, I451, I452, I454, I455, I456, I457, I458, I459, I460, I462, I463, I464, I466, I467, I468, I469, I470, I471, I472, I474, I475, I476, I477, I478, I479, I480, I481, I482, I483, I484, I485, I486, I488, I489, I490, I491, I492, I493, I494, I495, I496, I498, I499, I500, I501, I502, I503, I504, I505, I506, I507, I508, I509, I510, I511, I512, I514, I516, I517, I518, I519, I520, I521, I522, I524, I525, I526, I527, I528, I530, I531, I532, I533, I534, I535, I536, I537, I538, I539, I540, I541, I542, I543, I544, I546, I547, I548, I549, I550, I551, I552, I554, I555, I556, I557, I558, I559, I560, I562, I563, I564, I565, I566, I567, I568, I570, I572, I574, I575, I576, I578, I579, I580, I581, I582, I583, I584, I586, I587, I588, I590, I592, I594, I595, I596, I597, I598, I600, I601, I602, I603, I604, I605, I606, I607, I608, I609, I610, I612, I613, I614, I615, I616, I618, I619, I620, I621, I622, I623, I624, I625, I626, I628, I629, I630, I631, I632, I633, I634, I635, I636, I637, I638, I639, I640, I641, I642, I643, I644, I646, I647, I648, I649, I650, I652, I654, I655, I656, I657, I658, I659, I660, I661, I662, I664, I665, I666, I668, I669, I670, I671, I672, I673, I674, I675, I676, I677, I678, I679, I680, I681, I682, I683, I684, I685, I686, I687, I688, I690, I691, I692, I693, I694, I695, I696, I697, I698, I700, I701, I702, I704, I705, I706, I707, I708, I710, I711, I712, I713, I714, I715, I716, I718, I719, I720, I721, I722, I723, I724, I725, I726, I727, I728, I729, I730, I731, I732, I734, I735, I736, I737, I738, I740, I741, I742, I743, I744, I745, I746, I747, I748, I750, I752, I753, I754, I755, I756, I758, I759, I760, I762, I764, I765, I766, I767, I768, I770, I771, I772, I773, I774, I776, I777, I778, I779, I780, I781, I782, I784, I785, I786, I787, I788, I790, I791, I792, I793, I794, I796, I797, I798, I799, I800, I802, I804, I806, I808, I809, I810, I811, I812, I813, I814, I815, I816, I817, I818, I819, I820, I821, I822, I824, I825, I826, I827, I828, I829, I830, I831, I832, I833, I834, I836, I838, I839, I840, I842, I843, I844, I846, I848, I849, I850, I852, I853, I854, I856, I857, I858, I859, I860, I861, I862, I863, I864, I866, I868, I870, I871, I872, I873, I874, I875, I876, I877, I878, I879, I880, I881, I882, I884, I885, I886, I887, I888, I889, I890, I892, I893, I894, I895, I896, I898, I900, I901, I902, I903, I904, I905, I906, I907, I908, I909, I910, I911, I912, I913, I914, I915, I916, I917, I918, I919, I920, I921, I922, I923, I924, I925, I926, I927, I928, I929, I930, I932, I933, I934, I936, I937, I938, I939, I940, I941, I942, I943, I944, I945, I946, I947, I948, I950, I952, I953, I954, I956, I957, I958, I960, I962, I963, I964, I965, I966, I967, I968, I969, I970, I972, I973, I974, I975, I976, I977, I978, I980, I981, I982, I983, I984, I986, I987, I988, I989, I990, I991, I992, I993, I994, I995, I996, I998, I999, O0, O1, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15, O16, O17, O18, O19, O20, O21, O22, O23, O24, O25, O26, O27, O28, O29, O30, O31, O32, O33, O34, O35, O36, O37, O38, O39, O40, O41, O42, O43, O44, O45, O46, O47, O48, O49, O50, O51, O52, O53, O54, O55, O56, O57, O58, O59, O60, O61, O62, O63, O64, O65, O66, O67, O68, O69, O70, O71, O72, O73, O74, O75, O76, O77, O78, O79, O80, O81, O82, O83, O84, O85, O86, O87, O88, O89, O90, O91, O92, O93, O94, O95, O96, O97, O98, O99, O100, O101, O102, O103, O104, O105, O106, O107, O108, O109, O110, O111, O112, O113, O114, O115, O116, O117, O118, O119, O120, O121, O122, O123, O124, O125, O126, O127, O128, O129, O130, O131, O132, O133, O134, O135, O136, O137, O138, O139, O140, O141, O142, O143, O144, O145, O146, O147, O148, O149, O150, O151, O152, O153, O154, O155, O156, O157, O158, O159, O160, O161, O162, O163, O164, O165, O166, O167, O168, O169, O170, O171, O172, O173, O174, O175, O176, O177, O178, O179, O180, O181, O182, O183, O184, O185, O186, O187, O188, O189, O190, O191, O192, O193, O194, O195, O196, O197, O198, O199, O200, O201, O202, O203, O204, O205, O206, O207, O208, O209, O210, O211, O212, O213, O214, O215, O216, O217, O218, O219, O220, O221, O222, O223, O224, O225, O226, O227, O228, O229, O230, O231, O232, O233, O234, O235, O236, O237, O238, O239, O240, O241, O242, O243, O244, O245, O246, O247, O248, O249, O250, O251, O252, O253, O254, O255, O256, O257, O258, O259, O260, O261, O262, O263, O264, O265, O266, O267, O268, O269, O270, O271, O272, O273, O274, O275, O276, O277, O278, O279, O280, O281, O282, O283, O284, O285, O286, O287, O288, O289, O290, O291, O292, O293, O294, O295, O296, O297, O298, O299, O300, O301, O302, O303, O304, O305, O306, O307, O308, O309, O310, O311, O312, O313, O314, O315, O316, O317, O318, O319, O320, O321, O322, O323, O324, O325, O326, O327, O328, O329, O330, O331, O332, O333, O334, O335, O336, O337, O338, O339, O340, O341, O342, O343, O344, O345, O346, O347, O348, O349, O350, O351, O352, O353, O354, O355, O356, O357, O358, O359, O360, O361, O362, O363, O364, O365, O366, O367, O368, O369, O370, O371, O372, O373, O374, O375, O376, O377, O378, O379, O380, O381, O382, O383, O384, O385, O386, O387, O388, O389, O390, O391, O392, O393, O394, O395, O396, O397, O398, O399, O400, O401, O402, O403, O404, O405, O406, O407, O408, O409, O410, O411, O412, O413, O414, O415, O416, O417, O418, O419, O420, O421, O422, O423, O424, O425, O426, O427, O428, O429, O430, O431, O432, O433, O434, O435, O436, O437, O438, O439, O440, O441, O442, O443, O444, O445, O446, O447, O448, O449, O450, O451, O452, O453, O454, O455, O456, O457, O458, O459, O460, O461, O462, O463, O464, O465, O466, O467, O468, O469, O470, O471, O472, O473, O474, O475, O476, O477, O478, O479, O480, O481, O482, O483, O484, O485, O486, O487, O488, O489, O490, O491, O492, O493, O494, O495, O496, O497, O498, O499, O500, O501, O502, O503, O504, O505, O506, O507, O508, O509, O510, O511, O512, O513, O514, O515, O516, O517, O518, O519, O520, O521, O522, O523, O524, O525, O526, O527, O528, O529, O530, O531, O532, O533, O534, O535, O536, O537, O538, O539, O540, O541, O542, O543, O544, O545, O546, O547, O548, O549, O550, O551, O552, O553, O554, O555, O556, O557, O558, O559, O560, O561, O562, O563, O564, O565, O566, O567, O568, O569, O570, O571, O572, O573, O574, O575, O576, O577, O578, O579, O580, O581, O582, O583, O584, O585, O586, O587, O588, O589, O590, O591, O592, O593, O594, O595, O596, O597, O598, O599, O600, O601, O602, O603, O604, O605, O606, O607, O608, O609, O610, O611, O612, O613, O614, O615, O616, O617, O618, O619, O620, O621, O622, O623, O624, O625, O626, O627, O628, O629, O630, O631, O632, O633, O634, O635, O636, O637, O638, O639, O640, O641, O642, O643, O644, O645, O646, O647, O648, O649, O650, O651, O652, O653, O654, O655, O656, O657, O658, O659, O660, O661, O662, O663, O664, O665, O666, O667, O668, O669, O670, O671, O672, O673, O674, O675, O676, O677, O678, O679, O680, O681, O682, O683, O684, O685, O686, O687, O688, O689, O690, O691, O692, O693, O694, O695, O696, O697, O698, O699, O700, O701, O702, O703, O704, O705, O706, O707, O708, O709, O710, O711, O712, O713, O714, O715, O716, O717, O718, O719, O720, O721, O722, O723, O724, O725, O726, O727, O728, O729, O730, O731, O732, O733, O734, O735, O736, O737, O738, O739, O740, O741, O742, O743, O744, O745, O746, O747, O748, O749, O750, O751, O752, O753, O754, O755, O756, O757, O758, O759, O760, O761, O762, O763, O764, O765, O766, O767, O768, O769, O770, O771, O772, O773, O774, O775, O776, O777, O778, O779, O780, O781, O782, O783, O784, O785, O786, O787, O788, O789, O790, O791, O792, O793, O794, O795, O796, O797, O798, O799, O800, O801, O802, O803, O804, O805, O806, O807, O808, O809, O810, O811, O812, O813, O814, O815, O816, O817, O818, O819, O820, O821, O822, O823, O824, O825, O826, O827, O828, O829, O830, O831, O832, O833, O834, O835, O836, O837, O838, O839, O840, O841, O842, O843, O844, O845, O846, O847, O848, O849, O850, O851, O852, O853, O854, O855, O856, O857, O858, O859, O860, O861, O862, O863, O864, O865, O866, O867, O868, O869, O870, O871, O872, O873, O874, O875, O876, O877, O878, O879, O880, O881, O882, O883, O884, O885, O886, O887, O888, O889, O890, O891, O892, O893, O894, O895, O896, O897, O898, O899, O900, O901, O902, O903, O904, O905, O906, O907, O908, O909, O910, O911, O912, O913, O914, O915, O916, O917, O918, O919, O920, O921, O922, O923, O924, O925, O926, O927, O928, O929, O930, O931, O932, O933, O934, O935, O936, O937, O938, O939, O940, O941, O942, O943, O944, O945, O946, O947, O948, O949, O950, O951, O952, O953, O954, O955, O956, O957, O958, O959, O960, O961, O962, O963, O964, O965, O966, O967, O968, O969, O970, O971, O972, O973, O974, O975, O976, O977, O978, O979, O980, O981, O982, O983, O984, O985, O986, O987, O988, O989, O990, O991, O992, O993, O994, O995, O996, O997, O998, O999, O1000, O1001, O1002, O1003, O1004, O1005, O1006, O1007, O1008, O1009, O1010, O1011, O1012, O1013, O1014, O1015, O1016, O1017, O1018, O1019, O1020, O1021, O1022, O1023, O1024, O1025, O1026, O1027, O1028, O1029, O1030, O1031, O1032, O1033, O1034, O1035, O1036, O1037, O1038, O1039, O1040, O1041, O1042, O1043, O1044, O1045, O1046, O1047, O1048, O1049, O1050, O1051, O1052, O1053, O1054, O1055, O1056, O1057, O1058, O1059, O1060, O1061, O1062, O1063, O1064, O1065, O1066, O1067, O1068, O1069, O1070, O1071, O1072, O1073, O1074, O1075, O1076, O1077, O1078, O1079, O1080, O1081, O1082, O1083, O1084, O1085, O1086, O1087, O1088, O1089, O1090, O1091, O1092, O1093, O1094, O1095, O1096, O1097, O1098, O1099, O1100, O1101, O1102, O1103, O1104, O1105, O1106, O1107, O1108, O1109, O1110, O1111, O1112, O1113, O1114, O1115, O1116, O1117, O1118, O1119, O1120, O1121, O1122, O1123, O1124, O1125, O1126, O1127, O1128, O1129, O1130, O1131, O1132, O1133, O1134, O1135, O1136, O1137, O1138, O1139, O1140, O1141, O1142, O1143, O1144, O1145, O1146, O1147, O1148, O1149, O1150, O1151, O1152, O1153, O1154, O1155, O1156, O1157, O1158, O1159, O1160, O1161, O1162, O1163, O1164, O1165, O1166, O1167, O1168, O1169, O1170, O1171, O1172, O1173, O1174, O1175, O1176, O1177, O1178, O1179, O1180, O1181, O1182, O1183, O1184, O1185, O1186, O1187, O1188, O1189, O1190, O1191, O1192, O1193, O1194, O1195, O1196, O1197, O1198, O1199, O1200, O1201, O1202, O1203, O1204, O1205, O1206, O1207, O1208, O1209, O1210, O1211, O1212, O1213, O1214, O1215, O1216, O1217, O1218, O1219, O1220, O1221, O1222, O1223, O1224, O1225, O1226, O1227, O1228, O1229, O1230, O1231, O1232, O1233, O1234, O1235, O1236, O1237, O1238, O1239, O1240, O1241, O1242, O1243, O1244, O1245, O1246, O1247, O1248, O1249, O1250, O1251, O1252, O1253, O1254, O1255, O1256, O1257, O1258, O1259, O1260, O1261, O1262, O1263, O1264, O1265, O1266, O1267, O1268, O1269, O1270, O1271, O1272, O1273, O1274, O1275, O1276, O1277, O1278, O1279, O1280, O1281, O1282, O1283, O1284, O1285, O1286, O1287, O1288, O1289, O1290, O1291, O1292, O1293, O1294, O1295, O1296, O1297, O1298, O1299, O1300, O1301, O1302, O1303, O1304, O1305, O1306, O1307, O1308, O1309, O1310, O1311, O1312, O1313, O1314, O1315, O1316, O1317, O1318, O1319, O1320, O1321, O1322, O1323, O1324, O1325, O1326, O1327, O1328, O1329, O1330, O1331, O1332, O1333, O1334, O1335, O1336, O1337, O1338, O1339, O1340, O1341, O1342, O1343, O1344, O1345, O1346, O1347, O1348, O1349, O1350, O1351, O1352, O1353, O1354, O1355, O1356, O1357, O1358, O1359, O1360, O1361, O1362, O1363, O1364, O1365, O1366, O1367, O1368, O1369, O1370, O1371, O1372, O1373, O1374, O1375, O1376, O1377, O1378, O1379, O1380, O1381, O1382, O1383, O1384, O1385, O1386, O1387, O1388, O1389, O1390, O1391, O1392, O1393, O1394, O1395, O1396, O1397, O1398, O1399, O1400, O1401, O1402, O1403, O1404, O1405, O1406, O1407, O1408, O1409, O1410, O1411, O1412, O1413, O1414, O1415, O1416, O1417, O1418, O1419, O1420, O1421, O1422, O1423, O1424, O1425, O1426, O1427, O1428, O1429, O1430, O1431, O1432, O1433, O1434, O1435, O1436, O1437, O1438, O1439, O1440, O1441, O1442, O1443, O1444, O1445, O1446, O1447, O1448, O1449, O1450, O1451, O1452, O1453, O1454, O1455, O1456, O1457, O1458, O1459, O1460, O1461, O1462, O1463, O1464, O1465, O1466, O1467, O1468, O1469, O1470, O1471, O1472, O1473, O1474, O1475, O1476, O1477, O1478, O1479, O1480, O1481, O1482, O1483, O1484, O1485, O1486, O1487, O1488, O1489, O1490, O1491, O1492, O1493, O1494, O1495, O1496, O1497, O1498, O1499, O1500, O1501, O1502, O1503, O1504, O1505, O1506, O1507, O1508, O1509, O1510, O1511, O1512, O1513, O1514, O1515, O1516, O1517, O1518, O1519, O1520, O1521, O1522, O1523, O1524, O1525, O1526, O1527, O1528, O1529, O1530, O1531, O1532, O1533, O1534, O1535, O1536, O1537, O1538, O1539, O1540, O1541, O1542, O1543, O1544, O1545, O1546, O1547, O1548, O1549, O1550, O1551, O1552, O1553, O1554, O1555, O1556, O1557, O1558, O1559, O1560, O1561, O1562, O1563, O1564, O1565, O1566, O1567, O1568, O1569, O1570, O1571, O1572, O1573, O1574, O1575, O1576, O1577, O1578, O1579, O1580, O1581, O1582, O1583, O1584, O1585, O1586, O1587, O1588, O1589, O1590, O1591, O1592, O1593, O1594, O1595, O1596, O1597, O1598, O1599, O1600, O1601, O1602, O1603, O1604, O1605, O1606, O1607, O1608, O1609, O1610, O1611, O1612, O1613, O1614, O1615, O1616, O1617, O1618, O1619, O1620, O1621, O1622, O1623, O1624, O1625, O1626, O1627, O1628, O1629, O1630, O1631, O1632, O1633, O1634, O1635, O1636, O1637, O1638, O1639, O1640, O1641, O1642, O1643, O1644, O1645, O1646, O1647, O1648, O1649, O1650, O1651, O1652, O1653, O1654, O1655, O1656, O1657, O1658, O1659, O1660, O1661, O1662, O1663, O1664, O1665, O1666, O1667, O1668, O1669, O1670, O1671, O1672, O1673, O1674, O1675, O1676, O1677, O1678, O1679, O1680, O1681, O1682, O1683, O1684, O1685, O1686, O1687, O1688, O1689, O1690, O1691, O1692, O1693, O1694, O1695, O1696, O1697, O1698, O1699, O1700, O1701, O1702, O1703, O1704, O1705, O1706, O1707, O1708, O1709, O1710, O1711, O1712, O1713, O1714, O1715, O1716, O1717, O1718, O1719, O1720, O1721, O1722, O1723, O1724, O1725, O1726, O1727, O1728, O1729, O1730, O1731, O1732, O1733, O1734, O1735, O1736, O1737, O1738, O1739, O1740, O1741, O1742, O1743, O1744, O1745, O1746, O1747, O1748, O1749, O1750, O1751, O1752, O1753, O1754, O1755, O1756, O1757, O1758, O1759, O1760, O1761, O1762, O1763, O1764, O1765, O1766, O1767, O1768, O1769, O1770, O1771, O1772, O1773, O1774, O1775, O1776, O1777, O1778, O1779, O1780, O1781, O1782, O1783, O1784, O1785, O1786, O1787, O1788, O1789, O1790, O1791, O1792, O1793, O1794, O1795, O1796, O1797, O1798, O1799, O1800, O1801, O1802, O1803, O1804, O1805, O1806, O1807, O1808, O1809, O1810, O1811, O1812, O1813, O1814, O1815, O1816, O1817, O1818, O1819, O1820, O1821, O1822, O1823, O1824, O1825, O1826, O1827, O1828, O1829, O1830, O1831, O1832, O1833, O1834, O1835, O1836, O1837, O1838, O1839, O1840, O1841, O1842, O1843, O1844, O1845, O1846, O1847, O1848, O1849, O1850, O1851, O1852, O1853, O1854, O1855, O1856, O1857, O1858, O1859, O1860, O1861, O1862, O1863, O1864, O1865, O1866, O1867, O1868, O1869, O1870, O1871, O1872, O1873, O1874, O1875, O1876, O1877, O1878, O1879, O1880, O1881, O1882, O1883, O1884, O1885, O1886, O1887, O1888, O1889, O1890, O1891, O1892, O1893, O1894, O1895, O1896, O1897, O1898, O1899, O1900, O1901, O1902, O1903, O1904, O1905, O1906, O1907, O1908, O1909, O1910, O1911, O1912, O1913, O1914, O1915, O1916, O1917, O1918, O1919, O1920, O1921, O1922, O1923, O1924, O1925, O1926, O1927, O1928, O1929, O1930, O1931, O1932, O1933, O1934, O1935, O1936, O1937, O1938, O1939, O1940, O1941, O1942, O1943, O1944, O1945, O1946, O1947, O1948, O1949, O1950, O1951, O1952, O1953, O1954, O1955, O1956, O1957, O1958, O1959, O1960, O1961, O1962, O1963, O1964, O1965, O1966, O1967, O1968, O1969, O1970, O1971, O1972, O1973, O1974, O1975, O1976, O1977, O1978, O1979, O1980, O1981, O1982, O1983, O1984, O1985, O1986, O1987, O1988, O1989, O1990, O1991, O1992, O1993, O1994, O1995, O1996, O1997, O1998, O1999, O2000, O2001, O2002, O2003, O2004, O2005, O2006, O2007, O2008, O2009, O2010, O2011, O2012, O2013, O2014, O2015, O2016, O2017, O2018, O2019, O2020, O2021, O2022, O2023, O2024, O2025, O2026, O2027, O2028, O2029, O2030, O2031, O2032, O2033, O2034, O2035, O2036, O2037, O2038, O2039, O2040, O2041, O2042, O2043, O2044, O2045, O2046, O2047, O2048, O2049, O2050, O2051, O2052, O2053, O2054, O2055, O2056, O2057, O2058, O2059, O2060, O2061, O2062, O2063, O2064, O2065, O2066, O2067, O2068, O2069, O2070, O2071, O2072, O2073, O2074, O2075, O2076, O2077, O2078, O2079, O2080, O2081, O2082, O2083, O2084, O2085, O2086, O2087, O2088, O2089, O2090, O2091, O2092, O2093, O2094, O2095, O2096, O2097, O2098, O2099, O2100, O2101, O2102, O2103, O2104, O2105, O2106, O2107, O2108, O2109, O2110, O2111, O2112, O2113, O2114, O2115, O2116, O2117, O2118, O2119, O2120, O2121, O2122, O2123, O2124, O2125, O2126, O2127, O2128, O2129, O2130, O2131, O2132, O2133, O2134, O2135, O2136, O2137, O2138, O2139, O2140, O2141, O2142, O2143, O2144, O2145, O2146, O2147, O2148, O2149, O2150, O2151, O2152, O2153, O2154, O2155, O2156, O2157, O2158, O2159, O2160, O2161, O2162, O2163, O2164, O2165, O2166, O2167, O2168, O2169, O2170, O2171, O2172, O2173, O2174, O2175, O2176, O2177, O2178, O2179, O2180, O2181, O2182, O2183, O2184, O2185, O2186, O2187, O2188, O2189, O2190, O2191, O2192, O2193, O2194, O2195, O2196, O2197, O2198, O2199, O2200, O2201, O2202, O2203, O2204, O2205, O2206, O2207, O2208, O2209, O2210, O2211, O2212, O2213, O2214, O2215, O2216, O2217, O2218, O2219, O2220, O2221, O2222, O2223, O2224, O2225, O2226, O2227, O2228, O2229, O2230, O2231, O2232, O2233, O2234, O2235, O2236, O2237, O2238, O2239, O2240, O2241, O2242, O2243, O2244, O2245, O2246, O2247, O2248, O2249, O2250, O2251, O2252, O2253, O2254, O2255, O2256, O2257, O2258, O2259, O2260, O2261, O2262, O2263, O2264, O2265, O2266, O2267, O2268, O2269, O2270, O2271, O2272, O2273, O2274, O2275, O2276, O2277, O2278, O2279, O2280, O2281, O2282, O2283, O2284, O2285, O2286, O2287, O2288, O2289, O2290, O2291, O2292, O2293, O2294, O2295, O2296, O2297, O2298, O2299, O2300, O2301, O2302, O2303, O2304, O2305, O2306, O2307, O2308, O2309, O2310, O2311, O2312, O2313, O2314, O2315, O2316, O2317, O2318, O2319, O2320, O2321, O2322, O2323, O2324, O2325, O2326, O2327, O2328, O2329, O2330, O2331, O2332, O2333, O2334, O2335, O2336, O2337, O2338, O2339, O2340, O2341, O2342, O2343, O2344, O2345, O2346, O2347, O2348, O2349, O2350, O2351, O2352, O2353, O2354, O2355, O2356, O2357, O2358, O2359, O2360, O2361, O2362, O2363, O2364, O2365, O2366, O2367, O2368, O2369, O2370, O2371, O2372, O2373, O2374, O2375, O2376, O2377, O2378, O2379, O2380, O2381, O2382, O2383, O2384, O2385, O2386, O2387, O2388, O2389, O2390, O2391, O2392, O2393, O2394, O2395, O2396, O2397, O2398, O2399, O2400, O2401, O2402, O2403, O2404, O2405, O2406, O2407, O2408, O2409, O2410, O2411, O2412, O2413, O2414, O2415, O2416, O2417, O2418, O2419, O2420, O2421, O2422, O2423, O2424, O2425, O2426, O2427, O2428, O2429, O2430, O2431, O2432, O2433, O2434, O2435, O2436, O2437, O2438, O2439, O2440, O2441, O2442, O2443, O2444, O2445, O2446, O2447, O2448);
  input I0, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I16, I17, I18, I19, I20, I21, I22, I23, I24, I26, I27, I28, I29, I30, I31, I32, I34, I36, I38, I39, I40, I42, I43, I44, I45, I46, I48, I49, I50, I51, I52, I54, I55, I56, I57, I58, I60, I61, I62, I64, I65, I66, I68, I70, I71, I72, I74, I75, I76, I78, I79, I80, I81, I82, I84, I85, I86, I88, I90, I91, I92, I94, I95, I96, I98, I100, I102, I103, I104, I106, I108, I109, I110, I111, I112, I113, I114, I115, I116, I117, I118, I120, I121, I122, I123, I124, I126, I128, I130, I132, I134, I135, I136, I137, I138, I140, I142, I144, I145, I146, I147, I148, I150, I151, I152, I153, I154, I156, I157, I158, I160, I161, I162, I163, I164, I165, I166, I168, I169, I170, I171, I172, I174, I175, I176, I178, I179, I180, I181, I182, I184, I185, I186, I188, I190, I191, I192, I193, I194, I195, I196, I197, I198, I200, I202, I203, I204, I206, I207, I208, I209, I210, I212, I213, I214, I215, I216, I217, I218, I219, I220, I221, I222, I223, I224, I225, I226, I227, I228, I229, I230, I231, I232, I233, I234, I235, I236, I237, I238, I239, I240, I241, I242, I243, I244, I245, I246, I247, I248, I249, I250, I252, I253, I254, I255, I256, I257, I258, I259, I260, I261, I262, I263, I264, I266, I267, I268, I269, I270, I271, I272, I274, I276, I277, I278, I280, I282, I283, I284, I285, I286, I288, I289, I290, I291, I292, I294, I296, I297, I298, I299, I300, I301, I302, I303, I304, I305, I306, I308, I309, I310, I312, I313, I314, I315, I316, I317, I318, I319, I320, I322, I323, I324, I326, I328, I329, I330, I331, I332, I334, I335, I336, I337, I338, I339, I340, I342, I344, I346, I347, I348, I349, I350, I351, I352, I353, I354, I355, I356, I357, I358, I360, I361, I362, I364, I365, I366, I368, I370, I371, I372, I374, I375, I376, I378, I380, I382, I384, I385, I386, I387, I388, I389, I390, I391, I392, I393, I394, I396, I398, I400, I401, I402, I404, I405, I406, I407, I408, I409, I410, I412, I413, I414, I415, I416, I417, I418, I420, I421, I422, I423, I424, I426, I428, I429, I430, I431, I432, I433, I434, I435, I436, I437, I438, I439, I440, I441, I442, I443, I444, I445, I446, I447, I448, I450, I451, I452, I454, I455, I456, I457, I458, I459, I460, I462, I463, I464, I466, I467, I468, I469, I470, I471, I472, I474, I475, I476, I477, I478, I479, I480, I481, I482, I483, I484, I485, I486, I488, I489, I490, I491, I492, I493, I494, I495, I496, I498, I499, I500, I501, I502, I503, I504, I505, I506, I507, I508, I509, I510, I511, I512, I514, I516, I517, I518, I519, I520, I521, I522, I524, I525, I526, I527, I528, I530, I531, I532, I533, I534, I535, I536, I537, I538, I539, I540, I541, I542, I543, I544, I546, I547, I548, I549, I550, I551, I552, I554, I555, I556, I557, I558, I559, I560, I562, I563, I564, I565, I566, I567, I568, I570, I572, I574, I575, I576, I578, I579, I580, I581, I582, I583, I584, I586, I587, I588, I590, I592, I594, I595, I596, I597, I598, I600, I601, I602, I603, I604, I605, I606, I607, I608, I609, I610, I612, I613, I614, I615, I616, I618, I619, I620, I621, I622, I623, I624, I625, I626, I628, I629, I630, I631, I632, I633, I634, I635, I636, I637, I638, I639, I640, I641, I642, I643, I644, I646, I647, I648, I649, I650, I652, I654, I655, I656, I657, I658, I659, I660, I661, I662, I664, I665, I666, I668, I669, I670, I671, I672, I673, I674, I675, I676, I677, I678, I679, I680, I681, I682, I683, I684, I685, I686, I687, I688, I690, I691, I692, I693, I694, I695, I696, I697, I698, I700, I701, I702, I704, I705, I706, I707, I708, I710, I711, I712, I713, I714, I715, I716, I718, I719, I720, I721, I722, I723, I724, I725, I726, I727, I728, I729, I730, I731, I732, I734, I735, I736, I737, I738, I740, I741, I742, I743, I744, I745, I746, I747, I748, I750, I752, I753, I754, I755, I756, I758, I759, I760, I762, I764, I765, I766, I767, I768, I770, I771, I772, I773, I774, I776, I777, I778, I779, I780, I781, I782, I784, I785, I786, I787, I788, I790, I791, I792, I793, I794, I796, I797, I798, I799, I800, I802, I804, I806, I808, I809, I810, I811, I812, I813, I814, I815, I816, I817, I818, I819, I820, I821, I822, I824, I825, I826, I827, I828, I829, I830, I831, I832, I833, I834, I836, I838, I839, I840, I842, I843, I844, I846, I848, I849, I850, I852, I853, I854, I856, I857, I858, I859, I860, I861, I862, I863, I864, I866, I868, I870, I871, I872, I873, I874, I875, I876, I877, I878, I879, I880, I881, I882, I884, I885, I886, I887, I888, I889, I890, I892, I893, I894, I895, I896, I898, I900, I901, I902, I903, I904, I905, I906, I907, I908, I909, I910, I911, I912, I913, I914, I915, I916, I917, I918, I919, I920, I921, I922, I923, I924, I925, I926, I927, I928, I929, I930, I932, I933, I934, I936, I937, I938, I939, I940, I941, I942, I943, I944, I945, I946, I947, I948, I950, I952, I953, I954, I956, I957, I958, I960, I962, I963, I964, I965, I966, I967, I968, I969, I970, I972, I973, I974, I975, I976, I977, I978, I980, I981, I982, I983, I984, I986, I987, I988, I989, I990, I991, I992, I993, I994, I995, I996, I998, I999;
  output O0, O1, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15, O16, O17, O18, O19, O20, O21, O22, O23, O24, O25, O26, O27, O28, O29, O30, O31, O32, O33, O34, O35, O36, O37, O38, O39, O40, O41, O42, O43, O44, O45, O46, O47, O48, O49, O50, O51, O52, O53, O54, O55, O56, O57, O58, O59, O60, O61, O62, O63, O64, O65, O66, O67, O68, O69, O70, O71, O72, O73, O74, O75, O76, O77, O78, O79, O80, O81, O82, O83, O84, O85, O86, O87, O88, O89, O90, O91, O92, O93, O94, O95, O96, O97, O98, O99, O100, O101, O102, O103, O104, O105, O106, O107, O108, O109, O110, O111, O112, O113, O114, O115, O116, O117, O118, O119, O120, O121, O122, O123, O124, O125, O126, O127, O128, O129, O130, O131, O132, O133, O134, O135, O136, O137, O138, O139, O140, O141, O142, O143, O144, O145, O146, O147, O148, O149, O150, O151, O152, O153, O154, O155, O156, O157, O158, O159, O160, O161, O162, O163, O164, O165, O166, O167, O168, O169, O170, O171, O172, O173, O174, O175, O176, O177, O178, O179, O180, O181, O182, O183, O184, O185, O186, O187, O188, O189, O190, O191, O192, O193, O194, O195, O196, O197, O198, O199, O200, O201, O202, O203, O204, O205, O206, O207, O208, O209, O210, O211, O212, O213, O214, O215, O216, O217, O218, O219, O220, O221, O222, O223, O224, O225, O226, O227, O228, O229, O230, O231, O232, O233, O234, O235, O236, O237, O238, O239, O240, O241, O242, O243, O244, O245, O246, O247, O248, O249, O250, O251, O252, O253, O254, O255, O256, O257, O258, O259, O260, O261, O262, O263, O264, O265, O266, O267, O268, O269, O270, O271, O272, O273, O274, O275, O276, O277, O278, O279, O280, O281, O282, O283, O284, O285, O286, O287, O288, O289, O290, O291, O292, O293, O294, O295, O296, O297, O298, O299, O300, O301, O302, O303, O304, O305, O306, O307, O308, O309, O310, O311, O312, O313, O314, O315, O316, O317, O318, O319, O320, O321, O322, O323, O324, O325, O326, O327, O328, O329, O330, O331, O332, O333, O334, O335, O336, O337, O338, O339, O340, O341, O342, O343, O344, O345, O346, O347, O348, O349, O350, O351, O352, O353, O354, O355, O356, O357, O358, O359, O360, O361, O362, O363, O364, O365, O366, O367, O368, O369, O370, O371, O372, O373, O374, O375, O376, O377, O378, O379, O380, O381, O382, O383, O384, O385, O386, O387, O388, O389, O390, O391, O392, O393, O394, O395, O396, O397, O398, O399, O400, O401, O402, O403, O404, O405, O406, O407, O408, O409, O410, O411, O412, O413, O414, O415, O416, O417, O418, O419, O420, O421, O422, O423, O424, O425, O426, O427, O428, O429, O430, O431, O432, O433, O434, O435, O436, O437, O438, O439, O440, O441, O442, O443, O444, O445, O446, O447, O448, O449, O450, O451, O452, O453, O454, O455, O456, O457, O458, O459, O460, O461, O462, O463, O464, O465, O466, O467, O468, O469, O470, O471, O472, O473, O474, O475, O476, O477, O478, O479, O480, O481, O482, O483, O484, O485, O486, O487, O488, O489, O490, O491, O492, O493, O494, O495, O496, O497, O498, O499, O500, O501, O502, O503, O504, O505, O506, O507, O508, O509, O510, O511, O512, O513, O514, O515, O516, O517, O518, O519, O520, O521, O522, O523, O524, O525, O526, O527, O528, O529, O530, O531, O532, O533, O534, O535, O536, O537, O538, O539, O540, O541, O542, O543, O544, O545, O546, O547, O548, O549, O550, O551, O552, O553, O554, O555, O556, O557, O558, O559, O560, O561, O562, O563, O564, O565, O566, O567, O568, O569, O570, O571, O572, O573, O574, O575, O576, O577, O578, O579, O580, O581, O582, O583, O584, O585, O586, O587, O588, O589, O590, O591, O592, O593, O594, O595, O596, O597, O598, O599, O600, O601, O602, O603, O604, O605, O606, O607, O608, O609, O610, O611, O612, O613, O614, O615, O616, O617, O618, O619, O620, O621, O622, O623, O624, O625, O626, O627, O628, O629, O630, O631, O632, O633, O634, O635, O636, O637, O638, O639, O640, O641, O642, O643, O644, O645, O646, O647, O648, O649, O650, O651, O652, O653, O654, O655, O656, O657, O658, O659, O660, O661, O662, O663, O664, O665, O666, O667, O668, O669, O670, O671, O672, O673, O674, O675, O676, O677, O678, O679, O680, O681, O682, O683, O684, O685, O686, O687, O688, O689, O690, O691, O692, O693, O694, O695, O696, O697, O698, O699, O700, O701, O702, O703, O704, O705, O706, O707, O708, O709, O710, O711, O712, O713, O714, O715, O716, O717, O718, O719, O720, O721, O722, O723, O724, O725, O726, O727, O728, O729, O730, O731, O732, O733, O734, O735, O736, O737, O738, O739, O740, O741, O742, O743, O744, O745, O746, O747, O748, O749, O750, O751, O752, O753, O754, O755, O756, O757, O758, O759, O760, O761, O762, O763, O764, O765, O766, O767, O768, O769, O770, O771, O772, O773, O774, O775, O776, O777, O778, O779, O780, O781, O782, O783, O784, O785, O786, O787, O788, O789, O790, O791, O792, O793, O794, O795, O796, O797, O798, O799, O800, O801, O802, O803, O804, O805, O806, O807, O808, O809, O810, O811, O812, O813, O814, O815, O816, O817, O818, O819, O820, O821, O822, O823, O824, O825, O826, O827, O828, O829, O830, O831, O832, O833, O834, O835, O836, O837, O838, O839, O840, O841, O842, O843, O844, O845, O846, O847, O848, O849, O850, O851, O852, O853, O854, O855, O856, O857, O858, O859, O860, O861, O862, O863, O864, O865, O866, O867, O868, O869, O870, O871, O872, O873, O874, O875, O876, O877, O878, O879, O880, O881, O882, O883, O884, O885, O886, O887, O888, O889, O890, O891, O892, O893, O894, O895, O896, O897, O898, O899, O900, O901, O902, O903, O904, O905, O906, O907, O908, O909, O910, O911, O912, O913, O914, O915, O916, O917, O918, O919, O920, O921, O922, O923, O924, O925, O926, O927, O928, O929, O930, O931, O932, O933, O934, O935, O936, O937, O938, O939, O940, O941, O942, O943, O944, O945, O946, O947, O948, O949, O950, O951, O952, O953, O954, O955, O956, O957, O958, O959, O960, O961, O962, O963, O964, O965, O966, O967, O968, O969, O970, O971, O972, O973, O974, O975, O976, O977, O978, O979, O980, O981, O982, O983, O984, O985, O986, O987, O988, O989, O990, O991, O992, O993, O994, O995, O996, O997, O998, O999, O1000, O1001, O1002, O1003, O1004, O1005, O1006, O1007, O1008, O1009, O1010, O1011, O1012, O1013, O1014, O1015, O1016, O1017, O1018, O1019, O1020, O1021, O1022, O1023, O1024, O1025, O1026, O1027, O1028, O1029, O1030, O1031, O1032, O1033, O1034, O1035, O1036, O1037, O1038, O1039, O1040, O1041, O1042, O1043, O1044, O1045, O1046, O1047, O1048, O1049, O1050, O1051, O1052, O1053, O1054, O1055, O1056, O1057, O1058, O1059, O1060, O1061, O1062, O1063, O1064, O1065, O1066, O1067, O1068, O1069, O1070, O1071, O1072, O1073, O1074, O1075, O1076, O1077, O1078, O1079, O1080, O1081, O1082, O1083, O1084, O1085, O1086, O1087, O1088, O1089, O1090, O1091, O1092, O1093, O1094, O1095, O1096, O1097, O1098, O1099, O1100, O1101, O1102, O1103, O1104, O1105, O1106, O1107, O1108, O1109, O1110, O1111, O1112, O1113, O1114, O1115, O1116, O1117, O1118, O1119, O1120, O1121, O1122, O1123, O1124, O1125, O1126, O1127, O1128, O1129, O1130, O1131, O1132, O1133, O1134, O1135, O1136, O1137, O1138, O1139, O1140, O1141, O1142, O1143, O1144, O1145, O1146, O1147, O1148, O1149, O1150, O1151, O1152, O1153, O1154, O1155, O1156, O1157, O1158, O1159, O1160, O1161, O1162, O1163, O1164, O1165, O1166, O1167, O1168, O1169, O1170, O1171, O1172, O1173, O1174, O1175, O1176, O1177, O1178, O1179, O1180, O1181, O1182, O1183, O1184, O1185, O1186, O1187, O1188, O1189, O1190, O1191, O1192, O1193, O1194, O1195, O1196, O1197, O1198, O1199, O1200, O1201, O1202, O1203, O1204, O1205, O1206, O1207, O1208, O1209, O1210, O1211, O1212, O1213, O1214, O1215, O1216, O1217, O1218, O1219, O1220, O1221, O1222, O1223, O1224, O1225, O1226, O1227, O1228, O1229, O1230, O1231, O1232, O1233, O1234, O1235, O1236, O1237, O1238, O1239, O1240, O1241, O1242, O1243, O1244, O1245, O1246, O1247, O1248, O1249, O1250, O1251, O1252, O1253, O1254, O1255, O1256, O1257, O1258, O1259, O1260, O1261, O1262, O1263, O1264, O1265, O1266, O1267, O1268, O1269, O1270, O1271, O1272, O1273, O1274, O1275, O1276, O1277, O1278, O1279, O1280, O1281, O1282, O1283, O1284, O1285, O1286, O1287, O1288, O1289, O1290, O1291, O1292, O1293, O1294, O1295, O1296, O1297, O1298, O1299, O1300, O1301, O1302, O1303, O1304, O1305, O1306, O1307, O1308, O1309, O1310, O1311, O1312, O1313, O1314, O1315, O1316, O1317, O1318, O1319, O1320, O1321, O1322, O1323, O1324, O1325, O1326, O1327, O1328, O1329, O1330, O1331, O1332, O1333, O1334, O1335, O1336, O1337, O1338, O1339, O1340, O1341, O1342, O1343, O1344, O1345, O1346, O1347, O1348, O1349, O1350, O1351, O1352, O1353, O1354, O1355, O1356, O1357, O1358, O1359, O1360, O1361, O1362, O1363, O1364, O1365, O1366, O1367, O1368, O1369, O1370, O1371, O1372, O1373, O1374, O1375, O1376, O1377, O1378, O1379, O1380, O1381, O1382, O1383, O1384, O1385, O1386, O1387, O1388, O1389, O1390, O1391, O1392, O1393, O1394, O1395, O1396, O1397, O1398, O1399, O1400, O1401, O1402, O1403, O1404, O1405, O1406, O1407, O1408, O1409, O1410, O1411, O1412, O1413, O1414, O1415, O1416, O1417, O1418, O1419, O1420, O1421, O1422, O1423, O1424, O1425, O1426, O1427, O1428, O1429, O1430, O1431, O1432, O1433, O1434, O1435, O1436, O1437, O1438, O1439, O1440, O1441, O1442, O1443, O1444, O1445, O1446, O1447, O1448, O1449, O1450, O1451, O1452, O1453, O1454, O1455, O1456, O1457, O1458, O1459, O1460, O1461, O1462, O1463, O1464, O1465, O1466, O1467, O1468, O1469, O1470, O1471, O1472, O1473, O1474, O1475, O1476, O1477, O1478, O1479, O1480, O1481, O1482, O1483, O1484, O1485, O1486, O1487, O1488, O1489, O1490, O1491, O1492, O1493, O1494, O1495, O1496, O1497, O1498, O1499, O1500, O1501, O1502, O1503, O1504, O1505, O1506, O1507, O1508, O1509, O1510, O1511, O1512, O1513, O1514, O1515, O1516, O1517, O1518, O1519, O1520, O1521, O1522, O1523, O1524, O1525, O1526, O1527, O1528, O1529, O1530, O1531, O1532, O1533, O1534, O1535, O1536, O1537, O1538, O1539, O1540, O1541, O1542, O1543, O1544, O1545, O1546, O1547, O1548, O1549, O1550, O1551, O1552, O1553, O1554, O1555, O1556, O1557, O1558, O1559, O1560, O1561, O1562, O1563, O1564, O1565, O1566, O1567, O1568, O1569, O1570, O1571, O1572, O1573, O1574, O1575, O1576, O1577, O1578, O1579, O1580, O1581, O1582, O1583, O1584, O1585, O1586, O1587, O1588, O1589, O1590, O1591, O1592, O1593, O1594, O1595, O1596, O1597, O1598, O1599, O1600, O1601, O1602, O1603, O1604, O1605, O1606, O1607, O1608, O1609, O1610, O1611, O1612, O1613, O1614, O1615, O1616, O1617, O1618, O1619, O1620, O1621, O1622, O1623, O1624, O1625, O1626, O1627, O1628, O1629, O1630, O1631, O1632, O1633, O1634, O1635, O1636, O1637, O1638, O1639, O1640, O1641, O1642, O1643, O1644, O1645, O1646, O1647, O1648, O1649, O1650, O1651, O1652, O1653, O1654, O1655, O1656, O1657, O1658, O1659, O1660, O1661, O1662, O1663, O1664, O1665, O1666, O1667, O1668, O1669, O1670, O1671, O1672, O1673, O1674, O1675, O1676, O1677, O1678, O1679, O1680, O1681, O1682, O1683, O1684, O1685, O1686, O1687, O1688, O1689, O1690, O1691, O1692, O1693, O1694, O1695, O1696, O1697, O1698, O1699, O1700, O1701, O1702, O1703, O1704, O1705, O1706, O1707, O1708, O1709, O1710, O1711, O1712, O1713, O1714, O1715, O1716, O1717, O1718, O1719, O1720, O1721, O1722, O1723, O1724, O1725, O1726, O1727, O1728, O1729, O1730, O1731, O1732, O1733, O1734, O1735, O1736, O1737, O1738, O1739, O1740, O1741, O1742, O1743, O1744, O1745, O1746, O1747, O1748, O1749, O1750, O1751, O1752, O1753, O1754, O1755, O1756, O1757, O1758, O1759, O1760, O1761, O1762, O1763, O1764, O1765, O1766, O1767, O1768, O1769, O1770, O1771, O1772, O1773, O1774, O1775, O1776, O1777, O1778, O1779, O1780, O1781, O1782, O1783, O1784, O1785, O1786, O1787, O1788, O1789, O1790, O1791, O1792, O1793, O1794, O1795, O1796, O1797, O1798, O1799, O1800, O1801, O1802, O1803, O1804, O1805, O1806, O1807, O1808, O1809, O1810, O1811, O1812, O1813, O1814, O1815, O1816, O1817, O1818, O1819, O1820, O1821, O1822, O1823, O1824, O1825, O1826, O1827, O1828, O1829, O1830, O1831, O1832, O1833, O1834, O1835, O1836, O1837, O1838, O1839, O1840, O1841, O1842, O1843, O1844, O1845, O1846, O1847, O1848, O1849, O1850, O1851, O1852, O1853, O1854, O1855, O1856, O1857, O1858, O1859, O1860, O1861, O1862, O1863, O1864, O1865, O1866, O1867, O1868, O1869, O1870, O1871, O1872, O1873, O1874, O1875, O1876, O1877, O1878, O1879, O1880, O1881, O1882, O1883, O1884, O1885, O1886, O1887, O1888, O1889, O1890, O1891, O1892, O1893, O1894, O1895, O1896, O1897, O1898, O1899, O1900, O1901, O1902, O1903, O1904, O1905, O1906, O1907, O1908, O1909, O1910, O1911, O1912, O1913, O1914, O1915, O1916, O1917, O1918, O1919, O1920, O1921, O1922, O1923, O1924, O1925, O1926, O1927, O1928, O1929, O1930, O1931, O1932, O1933, O1934, O1935, O1936, O1937, O1938, O1939, O1940, O1941, O1942, O1943, O1944, O1945, O1946, O1947, O1948, O1949, O1950, O1951, O1952, O1953, O1954, O1955, O1956, O1957, O1958, O1959, O1960, O1961, O1962, O1963, O1964, O1965, O1966, O1967, O1968, O1969, O1970, O1971, O1972, O1973, O1974, O1975, O1976, O1977, O1978, O1979, O1980, O1981, O1982, O1983, O1984, O1985, O1986, O1987, O1988, O1989, O1990, O1991, O1992, O1993, O1994, O1995, O1996, O1997, O1998, O1999, O2000, O2001, O2002, O2003, O2004, O2005, O2006, O2007, O2008, O2009, O2010, O2011, O2012, O2013, O2014, O2015, O2016, O2017, O2018, O2019, O2020, O2021, O2022, O2023, O2024, O2025, O2026, O2027, O2028, O2029, O2030, O2031, O2032, O2033, O2034, O2035, O2036, O2037, O2038, O2039, O2040, O2041, O2042, O2043, O2044, O2045, O2046, O2047, O2048, O2049, O2050, O2051, O2052, O2053, O2054, O2055, O2056, O2057, O2058, O2059, O2060, O2061, O2062, O2063, O2064, O2065, O2066, O2067, O2068, O2069, O2070, O2071, O2072, O2073, O2074, O2075, O2076, O2077, O2078, O2079, O2080, O2081, O2082, O2083, O2084, O2085, O2086, O2087, O2088, O2089, O2090, O2091, O2092, O2093, O2094, O2095, O2096, O2097, O2098, O2099, O2100, O2101, O2102, O2103, O2104, O2105, O2106, O2107, O2108, O2109, O2110, O2111, O2112, O2113, O2114, O2115, O2116, O2117, O2118, O2119, O2120, O2121, O2122, O2123, O2124, O2125, O2126, O2127, O2128, O2129, O2130, O2131, O2132, O2133, O2134, O2135, O2136, O2137, O2138, O2139, O2140, O2141, O2142, O2143, O2144, O2145, O2146, O2147, O2148, O2149, O2150, O2151, O2152, O2153, O2154, O2155, O2156, O2157, O2158, O2159, O2160, O2161, O2162, O2163, O2164, O2165, O2166, O2167, O2168, O2169, O2170, O2171, O2172, O2173, O2174, O2175, O2176, O2177, O2178, O2179, O2180, O2181, O2182, O2183, O2184, O2185, O2186, O2187, O2188, O2189, O2190, O2191, O2192, O2193, O2194, O2195, O2196, O2197, O2198, O2199, O2200, O2201, O2202, O2203, O2204, O2205, O2206, O2207, O2208, O2209, O2210, O2211, O2212, O2213, O2214, O2215, O2216, O2217, O2218, O2219, O2220, O2221, O2222, O2223, O2224, O2225, O2226, O2227, O2228, O2229, O2230, O2231, O2232, O2233, O2234, O2235, O2236, O2237, O2238, O2239, O2240, O2241, O2242, O2243, O2244, O2245, O2246, O2247, O2248, O2249, O2250, O2251, O2252, O2253, O2254, O2255, O2256, O2257, O2258, O2259, O2260, O2261, O2262, O2263, O2264, O2265, O2266, O2267, O2268, O2269, O2270, O2271, O2272, O2273, O2274, O2275, O2276, O2277, O2278, O2279, O2280, O2281, O2282, O2283, O2284, O2285, O2286, O2287, O2288, O2289, O2290, O2291, O2292, O2293, O2294, O2295, O2296, O2297, O2298, O2299, O2300, O2301, O2302, O2303, O2304, O2305, O2306, O2307, O2308, O2309, O2310, O2311, O2312, O2313, O2314, O2315, O2316, O2317, O2318, O2319, O2320, O2321, O2322, O2323, O2324, O2325, O2326, O2327, O2328, O2329, O2330, O2331, O2332, O2333, O2334, O2335, O2336, O2337, O2338, O2339, O2340, O2341, O2342, O2343, O2344, O2345, O2346, O2347, O2348, O2349, O2350, O2351, O2352, O2353, O2354, O2355, O2356, O2357, O2358, O2359, O2360, O2361, O2362, O2363, O2364, O2365, O2366, O2367, O2368, O2369, O2370, O2371, O2372, O2373, O2374, O2375, O2376, O2377, O2378, O2379, O2380, O2381, O2382, O2383, O2384, O2385, O2386, O2387, O2388, O2389, O2390, O2391, O2392, O2393, O2394, O2395, O2396, O2397, O2398, O2399, O2400, O2401, O2402, O2403, O2404, O2405, O2406, O2407, O2408, O2409, O2410, O2411, O2412, O2413, O2414, O2415, O2416, O2417, O2418, O2419, O2420, O2421, O2422, O2423, O2424, O2425, O2426, O2427, O2428, O2429, O2430, O2431, O2432, O2433, O2434, O2435, O2436, O2437, O2438, O2439, O2440, O2441, O2442, O2443, O2444, O2445, O2446, O2447, O2448;
  wire W3276, W3244, W3245, W3246, W3247, W3255, W3256, W3263, W3278, W3279, W3284, W3285, W3291, W3294, W3296, W3299, W3300, W3301, W3210, W3181, W3185, W3186, W3187, W3190, W3200, W3205, W3206, W3209, W3215, W3216, W3217, W3222, W3223, W3224, W3229, W3232, W3233, W3237, W3238, W3239, W3381, W3383, W3389, W3391, W3398, W3399, W3401, W3404, W3409, W3412, W3417, W3379, W3423, W3426, W3438, W3450, W3452, W3454, W3308, W3310, W3316, W3325, W3335, W3336, W3337, W3338, W3339, W3344, W3351, W3362, W3374, W3376, W3378, W2996, W2949, W2952, W2955, W2961, W2963, W2969, W2970, W2974, W2977, W2982, W2986, W2989, W3002, W3003, W3007, W3013, W3015, W3017, W3018, W3019, W3020, W3022, W2911, W2875, W2877, W2878, W2886, W2891, W2898, W2899, W2900, W2905, W3026, W2927, W2928, W2934, W2937, W2940, W2942, W2944, W2945, W2946, W3100, W3104, W3105, W3107, W3111, W3113, W3117, W3118, W3119, W3122, W3093, W3134, W3135, W3141, W3142, W3154, W3171, W3062, W3027, W3029, W3030, W3036, W3041, W3047, W3056, W3063, W3064, W3067, W3070, W3071, W3078, W3081, W3084, W3088, W3090, W3880, W3891, W3901, W3902, W3910, W3914, W3917, W3918, W3877, W3929, W3932, W3933, W3945, W3946, W3947, W3813, W3816, W3820, W3826, W3827, W3830, W3831, W3832, W3838, W3844, W3862, W3863, W3865, W3870, W4064, W4036, W4047, W4054, W4063, W4025, W4078, W4081, W4084, W3960, W3963, W3966, W3968, W3974, W3979, W3980, W3812, W3991, W4007, W4008, W4012, W3549, W3554, W3556, W3560, W3575, W3577, W3580, W3582, W3583, W3544, W3594, W3599, W3606, W3609, W3623, W3624, W3503, W3461, W3464, W3472, W3473, W3480, W3489, W3490, W3496, W3505, W3509, W3511, W3519, W3523, W3525, W3528, W3533, W3538, W3542, W3543, W3722, W3734, W3735, W3736, W3744, W3749, W3750, W3709, W3761, W3764, W3769, W3780, W3793, W3811, W3636, W3639, W3642, W3659, W3661, W3664, W3672, W2874, W3683, W3687, W3690, W3691, W3695, W3697, W3698, W3705, W3708, W2047, W1999, W2000, W2002, W2006, W2014, W2029, W2040, W2044, W2046, W2048, W2051, W2054, W2055, W2057, W2058, W2062, W2063, W2068, W2070, W1963, W1928, W1931, W1932, W1938, W1942, W1944, W1945, W1947, W1949, W1950, W1955, W1956, W2076, W1966, W1968, W1969, W1970, W1974, W1980, W1988, W1990, W1991, W1993, W2172, W2147, W2150, W2155, W2158, W2159, W2160, W2161, W2162, W2164, W2168, W2169, W2178, W2180, W2185, W2188, W2190, W2192, W2193, W2195, W2078, W2080, W2082, W2085, W2088, W2089, W2093, W2099, W2106, W1922, W2111, W2116, W2122, W2128, W2130, W2131, W2133, W2138, W2140, W2141, W1735, W1707, W1709, W1711, W1720, W1721, W1722, W1731, W1705, W1737, W1740, W1741, W1743, W1744, W1745, W1746, W1748, W1749, W1752, W1755, W1756, W1673, W1640, W1642, W1643, W1645, W1648, W1651, W1652, W1659, W1661, W1665, W1668, W1672, W1761, W1680, W1689, W1691, W1692, W1693, W1695, W1697, W1699, W1701, W1702, W1884, W1845, W1846, W1851, W1853, W1854, W1860, W1865, W1866, W1873, W1876, W1881, W1844, W1886, W1887, W1890, W1895, W1897, W1907, W1909, W1916, W1919, W1811, W1762, W1763, W1764, W1779, W1785, W1789, W1797, W1801, W1804, W2214, W1813, W1819, W1821, W1824, W1825, W1832, W1834, W1835, W1841, W1842, W2632, W2640, W2641, W2646, W2652, W2659, W2660, W2630, W2674, W2675, W2680, W2682, W2687, W2694, W2703, W2708, W2710, W2714, W2584, W2556, W2562, W2567, W2571, W2572, W2573, W2574, W2575, W2579, W2582, W2716, W2588, W2591, W2595, W2599, W2601, W2622, W2624, W2625, W2829, W2804, W2805, W2807, W2812, W2815, W2816, W2817, W2801, W2834, W2845, W2847, W2856, W2859, W2863, W2864, W2871, W2872, W2751, W2720, W2721, W2729, W2730, W2731, W2736, W2737, W2739, W2749, W2536, W2758, W2759, W2769, W2774, W2777, W2781, W2789, W2793, W2795, W2290, W2291, W2293, W2296, W2308, W2310, W2314, W2324, W2325, W2289, W2337, W2338, W2347, W2350, W2351, W2354, W2357, W2358, W2371, W2374, W2378, W2259, W2216, W2222, W2223, W2225, W2233, W2234, W2239, W2241, W2243, W2385, W2260, W2265, W2266, W2268, W2270, W2273, W2275, W2276, W2278, W2279, W2281, W2498, W2463, W2467, W2468, W2470, W2474, W2479, W2483, W2486, W2490, W2494, W2496, W2455, W2506, W2508, W2512, W2513, W2519, W2520, W2521, W2534, W2424, W2388, W2393, W2394, W2395, W2396, W2399, W2400, W2402, W2403, W2405, W2408, W2415, W2425, W2430, W2439, W2441, W2442, W2446, W2447, W2448, W2452, W5710, W5737, W5637, W5638, W5658, W5659, W5763, W5674, W5679, W5680, W5852, W5848, W5807, W5788, W5824, W5836, W5454, W5436, W5437, W5442, W5452, W5468, W5470, W5483, W5348, W5351, W5354, W5363, W5371, W5400, W5408, W5409, W5564, W5567, W5588, W5616, W5494, W5511, W5529, W5547, W6329, W6334, W6267, W6262, W6022, W6015, W6055, W6075, W5936, W5938, W5964, W5985, W6009, W6232, W6082, W6133, W4559, W4535, W4542, W4558, W4569, W4578, W4585, W4588, W4589, W4602, W4604, W4480, W4452, W4454, W4467, W4607, W4491, W4506, W4514, W4515, W4517, W4520, W4521, W4522, W4527, W4684, W4686, W4695, W4707, W4675, W4723, W4725, W4736, W4748, W4749, W4608, W4613, W4615, W4622, W4627, W4630, W4640, W4647, W4653, W4657, W4659, W4669, W4170, W4174, W4176, W4177, W4194, W4203, W4215, W4216, W4168, W4236, W4245, W4250, W4253, W4262, W4264, W4131, W4094, W4099, W4100, W4102, W4103, W4106, W4120, W4128, W4267, W4132, W4142, W4146, W4147, W4157, W4390, W4357, W4359, W4364, W4371, W4380, W4381, W4382, W4383, W4386, W4389, W4392, W4398, W4405, W4413, W4423, W4270, W4280, W4281, W4290, W4293, W4296, W4301, W4302, W4304, W4755, W4313, W4336, W4337, W4343, W4346, W5136, W5141, W5143, W5144, W5165, W5176, W5181, W5183, W5186, W5090, W5062, W5067, W5072, W5075, W5076, W5085, W5101, W5118, W5274, W5282, W5283, W5286, W5296, W5301, W5302, W5206, W5208, W5218, W5250, W5254, W4824, W4827, W4830, W4833, W4848, W4851, W4869, W4879, W4881, W4889, W4762, W4766, W4767, W4769, W4780, W4783, W4789, W4800, W4801, W4808, W4810, W4985, W4999, W5005, W5007, W5011, W5030, W5031, W4916, W4918, W4934, W4935, W4938, W4939, W3251, W4962, W4964, W4969, W4977, W790, W797, W1427, W1147, W1426, W329, W1149, W334, W335, W336, W337, W338, W324, W339, W340, W341, W1418, W1154, W1416, W788, W787, W1414, W347, W1433, W307, W309, W1436, W310, W312, W1434, W314, W801, W315, W316, W799, W1411, W798, W1143, W318, W319, W1430, W320, W1145, W323, W1392, W372, W772, W1397, W1396, W376, W771, W1168, W770, W382, W383, W768, W774, W388, W389, W390, W1389, W1173, W392, W393, W1178, W395, W396, W757, W1401, W1410, W350, W1409, W784, W353, W781, W355, W356, W1404, W1159, W1160, W306, W361, W1163, W362, W363, W364, W365, W778, W777, W1166, W368, W853, W1109, W231, W1110, W860, W1488, W1112, W233, W857, W234, W856, W1108, W850, W1482, W1481, W240, W242, W845, W1119, W1474, W246, W222, W886, W1505, W210, W1096, W1504, W1098, W215, W1503, W217, W220, W221, W247, W223, W867, W1498, W1497, W1496, W227, W1107, W866, W229, W279, W821, W281, W283, W1129, W1130, W1449, W289, W1448, W1447, W291, W278, W811, W1445, W1135, W1442, W1137, W1441, W808, W806, W303, W804, W262, W1122, W1123, W838, W255, W837, W835, W258, W1128, W259, W260, W404, W263, W265, W269, W1460, W270, W273, W1458, W274, W275, W277, W665, W542, W1239, W1311, W546, W668, W547, W548, W667, W666, W541, W1305, W664, W663, W550, W1302, W657, W655, W1301, W1300, W1299, W653, W527, W515, W1229, W1230, W520, W1319, W521, W523, W524, W525, W678, W652, W676, W1234, W675, W673, W535, W1237, W672, W538, W539, W670, W1280, W642, W641, W582, W639, W633, W1259, W1283, W632, W1281, W1261, W574, W590, W591, W623, W622, W596, W1265, W606, W613, W1267, W1270, W617, W1253, W651, W1247, W561, W562, W650, W1249, W1250, W649, W647, W565, W646, W1324, W644, W567, W1291, W643, W569, W570, W571, W1289, W1288, W573, W1363, W431, W1369, W1368, W437, W739, W440, W442, W735, W1364, W430, W734, W733, W732, W444, W447, W730, W1356, W723, W454, W750, W407, W408, W409, W1185, W1186, W412, W1381, W415, W1379, W1189, W457, W749, W416, W748, W1374, W419, W1192, W426, W428, W429, W505, W1332, W494, W495, W499, W698, W500, W697, W695, W1329, W504, W1333, W692, W508, W689, W1225, W688, W511, W512, W513, W1226, W1227, W1345, W1206, W458, W1207, W1209, W461, W462, W718, W464, W468, W471, W1438, W1213, W1214, W478, W715, W484, W1339, W487, W1336, W1335, W491, W1565, W208, W955, W954, W1046, W1570, W115, W1047, W117, W1566, W112, W1048, W120, W1049, W948, W122, W1562, W1561, W123, W124, W961, W89, W90, W92, W95, W96, W965, W963, W1039, W1040, W126, W1041, W960, W1042, W959, W108, W1573, W109, W1537, W937, W935, W1543, W933, W1063, W932, W158, W925, W1549, W1536, W922, W921, W165, W1535, W167, W168, W169, W945, W1052, W128, W1558, W1055, W130, W1556, W947, W131, W1555, W87, W1057, W1058, W943, W133, W1551, W135, W1059, W141, W32, W1000, W998, W24, W25, W991, W28, W1621, W1620, W1617, W1017, W1615, W988, W35, W1021, W37, W1611, W1610, W985, W39, W13, W1638, W3, W1634, W4, W5, W1005, W10, W1630, W40, W1629, W1628, W15, W1014, W1627, W1015, W21, W1625, W968, W976, W1589, W1588, W73, W969, W1586, W1585, W75, W1583, W1592, W76, W967, W80, W81, W1035, W84, W1582, W979, W1023, W1024, W1607, W45, W55, W56, W57, W1572, W1027, W1028, W1600, W1599, W60, W61, W1596, W977, W1075, W1078, W894, W200, W892, W1091, W203, W1508, W1076, W1511, W888, W1531, W918, W206, W207, W1092, W1094, W1525, W1089, W1513, W182, W1514, W896, W192, W906, W1086, W1516, W187, W1084, W1085, W902, W1518, W920, W919, W887, W173, W1072, W693, W3616, W898, W694, W3983, W3614, W4528, W978, W4534, W4502, W4485, W972, W702, W3629, W973, W3625, W4495, W4498, W4504, W4508, W975, W3618, W683, W983, W982, W679, W4554, W3601, W4553, W3603, W682, W4740, W4547, W3608, W687, W3884, W3879, W618, W859, W3875, W685, W686, W3641, W4747, W4430, W719, W3644, W4437, W4009, W1639, W4438, W4439, W717, W849, W899, W4016, W4416, W724, W3652, W4421, W722, W903, W966, W848, W4010, W3648, W4429, W4468, W4743, W4463, W855, W970, W3634, W711, W707, W3866, W3867, W4564, W4458, W854, W3638, W712, W713, W714, W3992, W4450, W1008, W4446, W4003, W3510, W1001, W874, W3541, W877, W4661, W3905, W627, W4662, W4663, W3540, W891, W4651, W3900, W4724, W648, W3547, W997, W3552, W995, W873, W4642, W4700, W3527, W3927, W4694, W1006, W4690, W4702, W3518, W3517, W629, W635, W3529, W640, W3909, W4671, W880, W4715, W3535, W4667, W621, W671, W3896, W4590, W3590, W4600, W3588, W3587, W3957, W989, W4581, W984, W3512, W674, W3970, W4574, W619, W4572, W628, W656, W994, W3563, W4635, W654, W4633, W3568, W3570, W4632, W4631, W625, W3571, W3899, W4629, W881, W3977, W872, W658, W659, W4621, W3576, W990, W3578, W3954, W4184, W915, W4191, W3829, W824, W4183, W3737, W942, W4080, W4169, W939, W940, W793, W4172, W3825, W3747, W944, W792, W791, W822, W4178, W4182, W3745, W3742, W831, W4235, W779, W912, W4239, W3716, W4243, W776, W3711, W783, W826, W3729, W827, W946, W794, W828, W780, W829, W3721, W924, W3810, W4130, W818, W1009, W3809, W3806, W819, W923, W4134, W4136, W803, W802, W4141, W4101, W3815, W813, W812, W3814, W4109, W4112, W4115, W4118, W810, W4121, W934, W4150, W3819, W3763, W4088, W4159, W3759, W4161, W795, W930, W3797, W3796, W4144, W3794, W3792, W928, W3778, W3773, W4148, W3768, W4149, W3818, W745, W4348, W744, W4029, W4354, W4028, W3673, W743, W741, W4361, W962, W4362, W844, W4035, W4329, W4335, W957, W3688, W3849, W841, W4363, W3682, W4342, W746, W731, W3653, W729, W4394, W4399, W816, W726, W4378, W4368, W738, W3665, W4373, W737, W964, W736, W3657, W3656, W4021, W4283, W4268, W4274, W3706, W4276, W765, W4282, W3840, W4053, W4284, W4052, W950, W3704, W764, W832, W4247, W775, W3710, W4065, W911, W3837, W4254, W4260, W4061, W949, W3707, W769, W4317, W752, W4046, W953, W4041, W840, W4320, W3847, W4321, W4322, W4323, W956, W4298, W3701, W761, W4295, W3699, W3841, W4300, W907, W756, W4305, W755, W754, W952, W211, W5910, W204, W202, W5855, W228, W5863, W225, W219, W218, W5891, W216, W214, W180, W178, W177, W6006, W176, W175, W174, W196, W195, W194, W193, W5968, W5987, W185, W5725, W5686, W282, W5698, W271, W268, W287, W267, W266, W5748, W298, W304, W301, W300, W297, W5662, W5665, W5666, W293, W290, W237, W5815, W241, W5820, W239, W238, W244, W235, W5841, W5766, W5767, W254, W253, W252, W251, W250, W249, W245, W58, W67, W68, W54, W51, W42, W82, W97, W6283, W78, W72, W11, W22, W19, W14, W9, W8, W6, W2, W1, W30, W98, W27, W138, W145, W144, W142, W148, W6129, W134, W164, W6058, W161, W159, W157, W156, W154, W152, W151, W150, W149, W113, W111, W110, W107, W6226, W114, W106, W104, W103, W101, W6154, W129, W127, W5629, W121, W119, W118, W6197, W116, W5047, W522, W5025, W519, W5028, W517, W5037, W5056, W509, W507, W4996, W544, W543, W4972, W4978, W4984, W536, W533, W5074, W4997, W532, W5000, W531, W5004, W530, W529, W526, W5121, W5124, W486, W483, W482, W5140, W481, W476, W473, W472, W5164, W470, W469, W466, W5185, W503, W502, W5087, W5088, W5093, W497, W496, W545, W493, W5111, W5113, W490, W488, W4828, W4811, W589, W4816, W588, W587, W4826, W584, W4839, W4849, W579, W4855, W576, W4864, W4754, W611, W608, W603, W598, W595, W4797, W4798, W594, W592, W4937, W4922, W556, W4924, W4927, W4928, W555, W554, W553, W551, W4940, W4949, W4965, W4871, W4872, W4878, W568, W4891, W4893, W463, W564, W4906, W560, W559, W557, W5471, W5484, W360, W5487, W359, W5492, W5493, W357, W5506, W352, W386, W385, W5424, W5425, W5438, W379, W377, W5448, W373, W371, W370, W5595, W328, W5576, W5577, W327, W5587, W321, W5591, W330, W5613, W311, W348, W346, W345, W5525, W5527, W343, W342, W5546, W5558, W332, W5233, W5239, W443, W5253, W5232, W439, W438, W5267, W436, W5273, W5213, W5191, W460, W5199, W453, W452, W5210, W5211, W451, W450, W5221, W5222, W5225, W5228, W410, W5338, W406, W405, W5362, W413, W399, W398, W5381, W5396, W5288, W424, W5298, W5300, W421, W5307, W616, W5325, W414, W5331, W2611, W1317, W1315, W3508, W2597, W2602, W2603, W2606, W2607, W2586, W2612, W2613, W2614, W2616, W2619, W2623, W1310, W2631, W2634, W2563, W2545, W2549, W2552, W2557, W2559, W2561, W1327, W2637, W2565, W1326, W1323, W1322, W1321, W2576, W2580, W2683, W1287, W2688, W2690, W2695, W2699, W2700, W2701, W2706, W2709, W1282, W2717, W2719, W1278, W2722, W2726, W1277, W1294, W2638, W2639, W2643, W2648, W2651, W1297, W1295, W2544, W2664, W2666, W2668, W2669, W2671, W1293, W2676, W2677, W2453, W2426, W2443, W1362, W1360, W2449, W2451, W1358, W2423, W2454, W1357, W2457, W2458, W2459, W2460, W2461, W2462, W1355, W2397, W2386, W2387, W2389, W2391, W2392, W1380, W1378, W1377, W1354, W2398, W1376, W2401, W1373, W2412, W1370, W2421, W2422, W2526, W2505, W1341, W2507, W1340, W2509, W2511, W2516, W2522, W2523, W2504, W2528, W2531, W2537, W2539, W2540, W2542, W2488, W1353, W2471, W2472, W2473, W2477, W1351, W2482, W1349, W2487, W1276, W2489, W1348, W1347, W1346, W2497, W1344, W1343, W2503, W2997, W2971, W1196, W2976, W2980, W2983, W2984, W2993, W2994, W2999, W3001, W3005, W1187, W3009, W3011, W2951, W2926, W2931, W2932, W2941, W1208, W1205, W1203, W3016, W1201, W2958, W2959, W1200, W1199, W2964, W2965, W2968, W1198, W1161, W3069, W3074, W3076, W1158, W3080, W1157, W1164, W1156, W3087, W1155, W3092, W1152, W1150, W1183, W1179, W3023, W3025, W3028, W1175, W3031, W1174, W3039, W2923, W3042, W3045, W1169, W3049, W3050, W1167, W3055, W3060, W1165, W2806, W1258, W2791, W2792, W2794, W2796, W2797, W2800, W2802, W2803, W1254, W1252, W2808, W1248, W2814, W1245, W2819, W1244, W2823, W1266, W2733, W2735, W1272, W2740, W2747, W1268, W2752, W2753, W2825, W1264, W2764, W1263, W1262, W2770, W1260, W2786, W2884, W2887, W2892, W2893, W2894, W1231, W1221, W1220, W2901, W2902, W1216, W2913, W2921, W2831, W2833, W1241, W2841, W2842, W2844, W2383, W2860, W1232, W2865, W2866, W2867, W2869, W1540, W1879, W1880, W1550, W1885, W1548, W1891, W1541, W1904, W1905, W1875, W1911, W1913, W1914, W1917, W1918, W1924, W1926, W1557, W1833, W1836, W1837, W1839, W1840, W1564, W1560, W1847, W1559, W1929, W1855, W1857, W1858, W1861, W1863, W1553, W1870, W1872, W1552, W1982, W1520, W1971, W1973, W1977, W1978, W1981, W1962, W1985, W1986, W1994, W1995, W1997, W1998, W2001, W2005, W1506, W1528, W1930, W1934, W1935, W1936, W1937, W1940, W1946, W1830, W1948, W1527, W1526, W1952, W1524, W1957, W1960, W1700, W1681, W1683, W1686, W1688, W1690, W1694, W1696, W1616, W1624, W1704, W1713, W1718, W1605, W1723, W1730, W1732, W1733, W1663, W1637, W1644, W1649, W1631, W1654, W1657, W1660, W1736, W1664, W1666, W1671, W1626, W1675, W1676, W1677, W1678, W1679, W1574, W1794, W1799, W1800, W1577, W1802, W1805, W1807, W1575, W1810, W1790, W1812, W1815, W1816, W1817, W1822, W1823, W1569, W1568, W1584, W1738, W1747, W1750, W1751, W1754, W1758, W1759, W2008, W1768, W1772, W1773, W1774, W1775, W1776, W1777, W1579, W2272, W2253, W1421, W1419, W2263, W1417, W2267, W1415, W2249, W1413, W1412, W2280, W2284, W2286, W1408, W1407, W2294, W2219, W1440, W2197, W1435, W2210, W2211, W2212, W2295, W1431, W2226, W2230, W2240, W1425, W1423, W2246, W2247, W2352, W1395, W2336, W1393, W2339, W2341, W2343, W2349, W1390, W2332, W2356, W1387, W2361, W2364, W2369, W2370, W2376, W2382, W2311, W2297, W2298, W1402, W2300, W2302, W2305, W2306, W2309, W1399, W2187, W2312, W2313, W2316, W2318, W2320, W2321, W2322, W2323, W2079, W1493, W2059, W1490, W2065, W2066, W2069, W2072, W1484, W1483, W2053, W2081, W2083, W1478, W2090, W1476, W1475, W2098, W2026, W2011, W2013, W2017, W2018, W2019, W2023, W2025, W1473, W2030, W2033, W2034, W1502, W2042, W1500, W2050, W2149, W1456, W2153, W2154, W1455, W1454, W1453, W1451, W2163, W1457, W2167, W2170, W2171, W1446, W2174, W2175, W2177, W2179, W2181, W2124, W2100, W1472, W1471, W1470, W2113, W2119, W2129, W1466, W1465, W2132, W2134, W1463, W1461, W2142, W2146, W3333, W3140, W3429, W1133, W1054, W3271, W3230, W3371, W3196, W3370, W1033, W1018, W3334, W3148, W3189, W1090, W1121, W1067, W1032, W1051, W3202, W3321, W1016, W3385, W3384, W1138, W3420, W3281, W3280, W1036, W3328, W3329, W3277, W3199, W3377, W3484, W3447, W3359, W3444, W3358, W3462, W1095, W3164, W3242, W1022, W3355, W3243, W3167, W3353, W3250, W3248, W3455, W3352, W3349, W1025, W3350, W1031, W3152, W3155, W3156, W3182, W3262, W1066, W1064, W3160, W3331, W3259, W3179, W1062, W3258, W1093, W1127, W1061, W3163, W1102, W3442, W3468, W3312, W3121, W1045, W3287, W1073, W1141, W3212, W1117, W3106, W3109, W3302, W3123, W3414, W3390, W1114, W1113, W3495, W3408, W3293, W3112, W3411, W1146, W3410, W3320, W3115, W3292, W1115, W3396, W3307, W3116, W1082, W1074, W3120, W3288, W3110, W3298, W1077, W3400, W3319, W1043, W3318, W3218, W1071, W3315, W3314, W1139, W1462, W288, W224, W3731, W213, W3689, W5682, W2139, W1056, W3733, W2041, W2157, W5874, W2024, W5866, W292, W3366, W3748, W264, W1464, W212, W2045, W3730, W3395, W2135, W1459, W1044, W2151, W2036, W2035, W280, W2028, W958, W3738, W1452, W285, W2032, W2031, W284, W2027, W3361, W272, W1501, W2144, W1450, W2039, W5700, W3364, W2148, W286, W2037, W276, W941, W3360, W243, W5843, W5806, W1489, W2060, W3388, W3712, W2095, W3713, W1053, W3715, W230, W1492, W248, W3703, W1486, W3386, W1487, W2073, W2074, W236, W2102, W2077, W232, W2067, W1479, W2086, W2087, W1050, W1477, W2049, W256, W5860, W257, W2120, W2121, W1468, W2123, W2118, W2125, W2126, W2127, W3726, W226, W261, W3727, W5776, W2104, W2056, W3393, W3719, W2108, W1494, W2109, W2110, W3720, W2112, W5858, W3368, W1469, W2117, W5482, W5474, W1400, W2307, W1070, W2304, W2303, W3801, W1069, W3798, W1403, W375, W2326, W374, W5453, W3317, W5457, W2319, W369, W1398, W366, W3808, W5519, W351, W2282, W927, W5515, W349, W2277, W3789, W5510, W2274, W344, W3786, W1068, W2269, W2287, W3327, W1405, W358, W1406, W5496, W926, W3330, W2285, W3791, W3305, W2355, W1388, W2353, W3828, W5399, W391, W3304, W5404, W916, W3839, W397, W2363, W2362, W913, W2360, W1391, W2359, W5386, W394, W1386, W380, W3309, W2334, W5435, W2333, W1394, W378, W2330, W2329, W2328, W387, W2346, W3306, W5414, W2340, W917, W2198, W5622, W5623, W3345, W5627, W2201, W2200, W3343, W308, W2365, W3346, W2196, W305, W2215, W2213, W3765, W1437, W2209, W5615, W313, W2206, W5619, W295, W299, W5657, W1444, W3347, W3348, W938, W296, W2173, W294, W2194, W1439, W2191, W3757, W2189, W936, W2217, W2183, W5653, W3776, W2256, W2255, W2252, W2251, W2257, W2248, W3775, W5561, W3774, W3784, W3783, W5531, W2264, W929, W2262, W2261, W333, W5543, W2228, W5582, W326, W325, W3770, W2229, W322, W5581, W2227, W931, W1429, W2221, W2220, W2218, W2232, W1428, W2235, W2236, W2237, W2238, W3771, W1424, W331, W1422, W1590, W3479, W1587, W1760, W74, W1757, W3481, W71, W70, W69, W3482, W66, W79, W3566, W3565, W3564, W3562, W1770, W1769, W77, W993, W1766, W3550, W1598, W3483, W59, W3551, W1597, W1734, W3548, W65, W996, W1594, W1595, W83, W64, W63, W62, W1742, W3574, W1020, W1806, W1019, W105, W1803, W3474, W3471, W6237, W6241, W102, W987, W3463, W1571, W1820, W3586, W986, W1578, W1814, W3581, W6223, W1782, W1786, W1581, W1784, W1783, W91, W88, W1781, W1780, W86, W1778, W3567, W1796, W100, W1795, W1793, W1792, W3569, W1788, W94, W93, W1580, W20, W1670, W18, W1669, W1667, W17, W16, W1012, W3520, W3497, W23, W1004, W3498, W3526, W3499, W1007, W3524, W1674, W3500, W3522, W1647, W7, W3504, W1632, W1010, W1635, W1636, W1662, W3502, W12, W1658, W1682, W1655, W3515, W1653, W1717, W3546, W1604, W3486, W44, W43, W1724, W1715, W41, W1714, W1712, W38, W52, W1601, W1729, W1728, W1602, W53, W1708, W1603, W50, W49, W48, W1725, W46, W1003, W29, W3536, W1623, W3534, W1685, W3532, W1013, W26, W1614, W1612, W36, W1706, W1613, W34, W33, W3494, W31, W1618, W1002, W1619, W3654, W3421, W184, W183, W3422, W1959, W1964, W181, W1954, W1953, W1951, W188, W190, W1519, W3658, W189, W3646, W1521, W1038, W1037, W3419, W186, W1534, W6034, W1933, W170, W6039, W171, W1034, W166, W1927, W971, W1925, W3640, W3425, W179, W3428, W1941, W1939, W3430, W3431, W172, W5928, W2010, W2009, W3674, W2007, W3406, W3407, W2004, W5931, W205, W2003, W1507, W3671, W1509, W209, W2020, W3680, W3403, W3677, W3670, W2015, W3676, W2012, W191, W197, W3413, W1984, W1983, W3663, W1515, W1979, W3662, W3415, W1975, W1517, W1512, W201, W1510, W199, W1992, W3630, W198, W1989, W1987, W3666, W3605, W1867, W1554, W3607, W1862, W980, W1859, W1026, W1856, W3602, W1878, W3446, W1029, W132, W3610, W1871, W1869, W1567, W6186, W3597, W1838, W3457, W3458, W1827, W1826, W3456, W1852, W1850, W1849, W125, W1848, W1030, W981, W1843, W1563, W974, W1910, W155, W1539, W153, W1906, W3622, W6087, W3441, W1902, W163, W162, W1542, W160, W1538, W1915, W1912, W1883, W1545, W1889, W1546, W143, W146, W140, W139, W1882, W137, W136, W1894, W1900, W1899, W1898, W1896, W1544, W3402, W6101, W1892, W147, W1236, W4567, W1235, W2854, W4579, W4582, W3177, W4584, W680, W4549, W833, W834, W2868, W4555, W681, W2849, W3174, W4560, W1233, W2862, W662, W4605, W1240, W2836, W2835, W4609, W3180, W2838, W661, W4617, W2832, W660, W1126, W4586, W669, W2846, W4593, W2843, W4548, W4596, W4597, W4598, W4051, W2840, W2839, W1219, W4079, W4497, W4499, W4501, W4492, W4077, W4505, W701, W4509, W700, W4484, W2908, W2907, W4478, W704, W4482, W3166, W1217, W4486, W1218, W2903, W690, W830, W2883, W4537, W691, W4067, W684, W3169, W3170, W2873, W3172, W4074, W699, W1222, W2895, W4518, W4519, W696, W4073, W1223, W1224, W4526, W2889, W2888, W2763, W2766, W626, W2765, W4726, W624, W4015, W4732, W2760, W4014, W620, W4019, W2775, W631, W2773, W630, W2772, W2771, W847, W1118, W4712, W4713, W3201, W609, W2744, W1116, W4758, W612, W2742, W610, W2746, W4765, W607, W1271, W605, W604, W4006, W1273, W2755, W2754, W3203, W4744, W4745, W2776, W2750, W1269, W615, W4753, W842, W4037, W1251, W4646, W843, W4648, W4641, W645, W4655, W4656, W4032, W1120, W839, W4624, W1242, W3183, W4628, W4044, W2824, W1255, W4042, W2821, W1125, W1124, W2818, W4638, W1246, W4682, W638, W637, W2785, W4689, W634, W2783, W2782, W2779, W3198, W4697, W2798, W3192, W1256, W3194, W1257, W2909, W4024, W2788, W4677, W4023, W3038, W1170, W767, W4271, W4272, W3127, W4135, W4275, W4277, W4279, W766, W3037, W1171, W3035, W1172, W4257, W3054, W4249, W4251, W773, W3051, W4255, W4256, W3128, W4258, W4259, W4140, W3125, W3046, W3044, W4266, W4312, W4303, W1180, W1181, W1184, W807, W809, W4315, W3014, W4124, W4319, W4123, W4294, W3129, W805, W762, W3130, W4291, W4292, W760, W1177, W759, W4297, W3131, W4299, W3024, W758, W789, W4187, W4188, W4190, W796, W4162, W4195, W3086, W4198, W4204, W3097, W3102, W1148, W4171, W1151, W3099, W3098, W4175, W4164, W4179, W4180, W1153, W1142, W4227, W1144, W3068, W4233, W4234, W800, W4241, W3061, W3059, W3058, W3057, W4206, W4209, W785, W4212, W3008, W782, W3079, W3077, W4221, W3075, W721, W4092, W3157, W4427, W2950, W2939, W4431, W1210, W2936, W3150, W2960, W4098, W4402, W727, W4406, W2957, W2956, W4410, W817, W2954, W2953, W1202, W725, W825, W2919, W2917, W710, W2916, W4082, W2914, W1215, W709, W708, W2912, W706, W2910, W705, W2925, W1211, W1212, W4441, W3159, W4447, W728, W2924, W716, W4085, W823, W3162, W4352, W747, W1134, W2992, W4113, W2995, W4353, W2988, W4355, W2987, W1193, W751, W1136, W3138, W4327, W3004, W4330, W4331, W4333, W4334, W1190, W1191, W814, W4379, W2972, W4104, W2967, W815, W4393, W4395, W4396, W4397, W1132, W4111, W740, W1194, W4366, W4367, W2981, W4369, W2979, W2978, W3144, W2975, W4376, W4377, W5175, W3894, W5168, W2492, W893, W467, W5180, W465, W5182, W3890, W2501, W5149, W477, W5156, W3888, W475, W474, W1342, W3897, W3264, W2495, W5204, W3881, W895, W2469, W3883, W2466, W5215, W2465, W2464, W3269, W3887, W2485, W2484, W1350, W3267, W2481, W5148, W2478, W3270, W2476, W2475, W1352, W498, W2541, W885, W2538, W884, W5100, W2535, W2533, W3913, W3912, W2530, W1330, W2551, W2548, W501, W5080, W2529, W5084, W3921, W883, W5135, W889, W3903, W1338, W5139, W890, W3260, W480, W479, W3898, W492, W3911, W3257, W2524, W3907, W489, W1334, W1337, W3273, W5122, W2515, W2514, W485, W5127, W5327, W908, W3848, W1081, W1382, W411, W910, W418, W2410, W423, W2407, W422, W905, W420, W1372, W417, W2404, W3852, W1375, W5314, W1083, W2372, W5357, W1385, W3834, W403, W402, W3297, W401, W400, W2367, W2379, W1080, W2381, W2380, W5345, W2411, W1383, W2377, W1079, W2375, W1384, W1365, W1359, W1361, W2444, W901, W445, W1366, W2438, W441, W2436, W2434, W5224, W3874, W897, W2456, W449, W2432, W3275, W1088, W448, W1087, W5280, W2419, W2417, W2420, W2414, W427, W5290, W2413, W425, W3860, W1367, W2428, W2427, W3283, W904, W434, W3286, W433, W5275, W432, W3986, W4868, W3985, W2684, W4865, W1111, W4877, W1290, W4880, W858, W4883, W4856, W580, W3213, W1286, W4852, W2693, W578, W2692, W4859, W4861, W575, W1296, W4904, W863, W864, W563, W4908, W4909, W2661, W4902, W2658, W4915, W558, W3969, W2656, W2655, W3975, W1292, W3221, W566, W2672, W3225, W2670, W3976, W581, W4895, W4897, W2665, W2723, W852, W2727, W4001, W2725, W2724, W4791, W593, W4803, W4000, W3999, W1279, W597, W601, W600, W599, W851, W1274, W4004, W4786, W4787, W1275, W3208, W585, W3211, W583, W1284, W4840, W2697, W2696, W2718, W4812, W2715, W2713, W2712, W865, W2705, W2704, W586, W1320, W2590, W2589, W3942, W1318, W2583, W1316, W2578, W2577, W5029, W518, W875, W3937, W516, W2598, W1313, W871, W1314, W5001, W5002, W1104, W1103, W528, W5009, W5010, W2593, W2592, W2558, W5055, W879, W5057, W1097, W1099, W1328, W0, W5066, W3924, W506, W3936, W1325, W876, W2569, W5043, W2568, W2566, W878, W5049, W2564, W510, W868, W2635, W4945, W2633, W4953, W549, W2629, W2653, W1298, W3967, W2647, W2645, W1307, W2642, W1303, W3964, W3231, W552, W537, W3952, W540, W2610, W2609, W2608, W4986, W3950, W870, W4959, W2627, W1308, W869, W2621, W2620, W4968, W1105, W2618, W3956, W4973;

  NOR2X1 G0 (.A1(W726), .A2(W403), .ZN(W3276));
  NOR2X1 G1 (.A1(W1253), .A2(I64), .ZN(W3244));
  NOR2X1 G2 (.A1(W825), .A2(W1671), .ZN(W3245));
  NOR2X1 G3 (.A1(W1232), .A2(W760), .ZN(W3246));
  NOR2X1 G4 (.A1(W1486), .A2(W1314), .ZN(W3247));
  NOR2X1 G5 (.A1(W2629), .A2(W1970), .ZN(O412));
  NOR2X1 G6 (.A1(W863), .A2(W1730), .ZN(O413));
  NOR2X1 G7 (.A1(I780), .A2(W245), .ZN(O415));
  NOR2X1 G8 (.A1(W425), .A2(W1010), .ZN(W3255));
  NOR2X1 G9 (.A1(I402), .A2(W595), .ZN(W3256));
  NOR2X1 G10 (.A1(W954), .A2(W249), .ZN(W3263));
  NOR2X1 G11 (.A1(W953), .A2(I266), .ZN(O418));
  NOR2X1 G12 (.A1(W1847), .A2(I268), .ZN(O419));
  NOR2X1 G13 (.A1(W3058), .A2(W1135), .ZN(O410));
  NOR2X1 G14 (.A1(W3069), .A2(W156), .ZN(W3278));
  NOR2X1 G15 (.A1(W705), .A2(I144), .ZN(W3279));
  NOR2X1 G16 (.A1(W1401), .A2(W3087), .ZN(W3284));
  NOR2X1 G17 (.A1(I701), .A2(W2079), .ZN(W3285));
  NOR2X1 G18 (.A1(W3087), .A2(W731), .ZN(O423));
  NOR2X1 G19 (.A1(W1823), .A2(W73), .ZN(W3291));
  NOR2X1 G20 (.A1(W783), .A2(I825), .ZN(W3294));
  NOR2X1 G21 (.A1(W2735), .A2(W20), .ZN(O425));
  NOR2X1 G22 (.A1(W1814), .A2(I140), .ZN(W3296));
  NOR2X1 G23 (.A1(W119), .A2(I310), .ZN(W3299));
  NOR2X1 G24 (.A1(W685), .A2(I665), .ZN(W3300));
  NOR2X1 G25 (.A1(W285), .A2(W2287), .ZN(W3301));
  NOR2X1 G26 (.A1(I799), .A2(I337), .ZN(W3210));
  NOR2X1 G27 (.A1(W46), .A2(I18), .ZN(W3181));
  NOR2X1 G28 (.A1(I937), .A2(W2847), .ZN(O393));
  NOR2X1 G29 (.A1(I902), .A2(W127), .ZN(W3185));
  NOR2X1 G30 (.A1(W2839), .A2(I469), .ZN(W3186));
  NOR2X1 G31 (.A1(W130), .A2(I862), .ZN(W3187));
  NOR2X1 G32 (.A1(W2795), .A2(W1723), .ZN(O394));
  NOR2X1 G33 (.A1(W1435), .A2(I898), .ZN(W3190));
  NOR2X1 G34 (.A1(W1643), .A2(W2521), .ZN(O397));
  NOR2X1 G35 (.A1(W1236), .A2(I202), .ZN(W3200));
  NOR2X1 G36 (.A1(W804), .A2(W630), .ZN(W3205));
  NOR2X1 G37 (.A1(W180), .A2(W485), .ZN(W3206));
  NOR2X1 G38 (.A1(W2109), .A2(W74), .ZN(W3209));
  NOR2X1 G39 (.A1(I870), .A2(W1621), .ZN(O426));
  NOR2X1 G40 (.A1(W1301), .A2(W1679), .ZN(W3215));
  NOR2X1 G41 (.A1(W1421), .A2(W3015), .ZN(W3216));
  NOR2X1 G42 (.A1(I264), .A2(W13), .ZN(W3217));
  NOR2X1 G43 (.A1(I266), .A2(W2653), .ZN(W3222));
  NOR2X1 G44 (.A1(W1297), .A2(W3007), .ZN(W3223));
  NOR2X1 G45 (.A1(W770), .A2(W1067), .ZN(W3224));
  NOR2X1 G46 (.A1(W2189), .A2(W2976), .ZN(W3229));
  NOR2X1 G47 (.A1(W2519), .A2(W1231), .ZN(W3232));
  NOR2X1 G48 (.A1(W2620), .A2(W322), .ZN(W3233));
  NOR2X1 G49 (.A1(W344), .A2(W151), .ZN(W3237));
  NOR2X1 G50 (.A1(W1353), .A2(W1673), .ZN(W3238));
  NOR2X1 G51 (.A1(W2715), .A2(W254), .ZN(W3239));
  NOR2X1 G52 (.A1(W2739), .A2(W1205), .ZN(O455));
  NOR2X1 G53 (.A1(W1592), .A2(W787), .ZN(W3381));
  NOR2X1 G54 (.A1(I629), .A2(W1978), .ZN(W3383));
  NOR2X1 G55 (.A1(W1561), .A2(W779), .ZN(W3389));
  NOR2X1 G56 (.A1(W1136), .A2(I682), .ZN(W3391));
  NOR2X1 G57 (.A1(I831), .A2(W2246), .ZN(O452));
  NOR2X1 G58 (.A1(I564), .A2(W2411), .ZN(W3398));
  NOR2X1 G59 (.A1(W667), .A2(W3238), .ZN(W3399));
  NOR2X1 G60 (.A1(W2536), .A2(W1951), .ZN(W3401));
  NOR2X1 G61 (.A1(W1978), .A2(I423), .ZN(W3404));
  NOR2X1 G62 (.A1(I980), .A2(W3058), .ZN(W3409));
  NOR2X1 G63 (.A1(W1406), .A2(W242), .ZN(W3412));
  NOR2X1 G64 (.A1(W1802), .A2(W3296), .ZN(W3417));
  NOR2X1 G65 (.A1(W2122), .A2(W2709), .ZN(W3379));
  NOR2X1 G66 (.A1(I289), .A2(I464), .ZN(W3423));
  NOR2X1 G67 (.A1(W2469), .A2(I163), .ZN(W3426));
  NOR2X1 G68 (.A1(W3308), .A2(W2733), .ZN(O460));
  NOR2X1 G69 (.A1(W1910), .A2(W3183), .ZN(O461));
  NOR2X1 G70 (.A1(W3018), .A2(W3391), .ZN(O463));
  NOR2X1 G71 (.A1(W2975), .A2(W1230), .ZN(W3438));
  NOR2X1 G72 (.A1(W2466), .A2(W458), .ZN(O467));
  NOR2X1 G73 (.A1(W1671), .A2(W1375), .ZN(O468));
  NOR2X1 G74 (.A1(W3383), .A2(W2903), .ZN(O469));
  NOR2X1 G75 (.A1(I441), .A2(W101), .ZN(W3450));
  NOR2X1 G76 (.A1(W3360), .A2(W376), .ZN(W3452));
  NOR2X1 G77 (.A1(I289), .A2(W5), .ZN(W3454));
  NOR2X1 G78 (.A1(W3061), .A2(W860), .ZN(O434));
  NOR2X1 G79 (.A1(W2629), .A2(W1644), .ZN(W3308));
  NOR2X1 G80 (.A1(W1382), .A2(W1628), .ZN(W3310));
  NOR2X1 G81 (.A1(W1915), .A2(W752), .ZN(O427));
  NOR2X1 G82 (.A1(W2169), .A2(I135), .ZN(W3316));
  NOR2X1 G83 (.A1(I834), .A2(W2001), .ZN(O430));
  NOR2X1 G84 (.A1(W275), .A2(W152), .ZN(W3325));
  NOR2X1 G85 (.A1(W22), .A2(I857), .ZN(O433));
  NOR2X1 G86 (.A1(W2235), .A2(W1200), .ZN(W3335));
  NOR2X1 G87 (.A1(W2902), .A2(I355), .ZN(W3336));
  NOR2X1 G88 (.A1(W1563), .A2(W36), .ZN(W3337));
  NOR2X1 G89 (.A1(W852), .A2(W2353), .ZN(W3338));
  NOR2X1 G90 (.A1(W238), .A2(I346), .ZN(W3339));
  NOR2X1 G91 (.A1(I262), .A2(W870), .ZN(O392));
  NOR2X1 G92 (.A1(W813), .A2(I118), .ZN(W3344));
  NOR2X1 G93 (.A1(W2374), .A2(W3345), .ZN(W3351));
  NOR2X1 G94 (.A1(W530), .A2(I250), .ZN(O439));
  NOR2X1 G95 (.A1(W2981), .A2(W2275), .ZN(W3362));
  NOR2X1 G96 (.A1(W3331), .A2(I248), .ZN(O440));
  NOR2X1 G97 (.A1(W1168), .A2(W510), .ZN(O441));
  NOR2X1 G98 (.A1(W2295), .A2(W1551), .ZN(O444));
  NOR2X1 G99 (.A1(W3081), .A2(W2980), .ZN(O445));
  NOR2X1 G100 (.A1(W272), .A2(W1697), .ZN(W3374));
  NOR2X1 G101 (.A1(W974), .A2(I879), .ZN(W3376));
  NOR2X1 G102 (.A1(W360), .A2(W1929), .ZN(W3378));
  NOR2X1 G103 (.A1(W2608), .A2(W453), .ZN(W2996));
  NOR2X1 G104 (.A1(W16), .A2(W1955), .ZN(W2949));
  NOR2X1 G105 (.A1(W1361), .A2(I350), .ZN(W2952));
  NOR2X1 G106 (.A1(W239), .A2(W2461), .ZN(W2955));
  NOR2X1 G107 (.A1(W1470), .A2(W1406), .ZN(W2961));
  NOR2X1 G108 (.A1(W1239), .A2(W2814), .ZN(W2963));
  NOR2X1 G109 (.A1(W1983), .A2(I550), .ZN(W2969));
  NOR2X1 G110 (.A1(W2883), .A2(W1865), .ZN(W2970));
  NOR2X1 G111 (.A1(W1796), .A2(W734), .ZN(W2974));
  NOR2X1 G112 (.A1(W451), .A2(W2487), .ZN(W2977));
  NOR2X1 G113 (.A1(W829), .A2(W850), .ZN(W2982));
  NOR2X1 G114 (.A1(W1814), .A2(I860), .ZN(W2986));
  NOR2X1 G115 (.A1(W140), .A2(W923), .ZN(W2989));
  NOR2X1 G116 (.A1(W22), .A2(W795), .ZN(O333));
  NOR2X1 G117 (.A1(I610), .A2(W2172), .ZN(O342));
  NOR2X1 G118 (.A1(W651), .A2(W1150), .ZN(W3002));
  NOR2X1 G119 (.A1(W325), .A2(W1221), .ZN(W3003));
  NOR2X1 G120 (.A1(W410), .A2(W856), .ZN(W3007));
  NOR2X1 G121 (.A1(W1697), .A2(W2699), .ZN(W3013));
  NOR2X1 G122 (.A1(I564), .A2(W2310), .ZN(W3015));
  NOR2X1 G123 (.A1(W2840), .A2(I344), .ZN(W3017));
  NOR2X1 G124 (.A1(I460), .A2(W1477), .ZN(W3018));
  NOR2X1 G125 (.A1(I780), .A2(W195), .ZN(W3019));
  NOR2X1 G126 (.A1(W2898), .A2(W1756), .ZN(W3020));
  NOR2X1 G127 (.A1(W1693), .A2(W2396), .ZN(O346));
  NOR2X1 G128 (.A1(W472), .A2(W2388), .ZN(W3022));
  NOR2X1 G129 (.A1(I727), .A2(W603), .ZN(W2911));
  NOR2X1 G130 (.A1(W2110), .A2(W1689), .ZN(W2875));
  NOR2X1 G131 (.A1(W1776), .A2(W1676), .ZN(W2877));
  NOR2X1 G132 (.A1(W1810), .A2(W2212), .ZN(W2878));
  NOR2X1 G133 (.A1(W1234), .A2(W2417), .ZN(W2886));
  NOR2X1 G134 (.A1(I648), .A2(W1390), .ZN(O318));
  NOR2X1 G135 (.A1(W692), .A2(I415), .ZN(W2891));
  NOR2X1 G136 (.A1(W2793), .A2(I457), .ZN(O319));
  NOR2X1 G137 (.A1(W656), .A2(I848), .ZN(W2898));
  NOR2X1 G138 (.A1(I51), .A2(W2), .ZN(W2899));
  NOR2X1 G139 (.A1(W2220), .A2(W1561), .ZN(W2900));
  NOR2X1 G140 (.A1(W1444), .A2(W1871), .ZN(O321));
  NOR2X1 G141 (.A1(W1054), .A2(I2), .ZN(W2905));
  NOR2X1 G142 (.A1(W308), .A2(W2147), .ZN(W3026));
  NOR2X1 G143 (.A1(W1651), .A2(I355), .ZN(O325));
  NOR2X1 G144 (.A1(W2724), .A2(W1093), .ZN(W2927));
  NOR2X1 G145 (.A1(I958), .A2(W2682), .ZN(W2928));
  NOR2X1 G146 (.A1(W1088), .A2(W1203), .ZN(O329));
  NOR2X1 G147 (.A1(W2324), .A2(W2751), .ZN(W2934));
  NOR2X1 G148 (.A1(W1378), .A2(W1540), .ZN(W2937));
  NOR2X1 G149 (.A1(W1571), .A2(W1545), .ZN(W2940));
  NOR2X1 G150 (.A1(I987), .A2(W2236), .ZN(W2942));
  NOR2X1 G151 (.A1(I910), .A2(I534), .ZN(W2944));
  NOR2X1 G152 (.A1(I335), .A2(I756), .ZN(W2945));
  NOR2X1 G153 (.A1(W1468), .A2(W1209), .ZN(W2946));
  NOR2X1 G154 (.A1(W200), .A2(W1214), .ZN(O371));
  NOR2X1 G155 (.A1(W1130), .A2(W2030), .ZN(O365));
  NOR2X1 G156 (.A1(W2055), .A2(I58), .ZN(W3100));
  NOR2X1 G157 (.A1(W1571), .A2(W389), .ZN(O367));
  NOR2X1 G158 (.A1(W2169), .A2(W1989), .ZN(W3104));
  NOR2X1 G159 (.A1(W2466), .A2(I138), .ZN(W3105));
  NOR2X1 G160 (.A1(W2867), .A2(W2913), .ZN(W3107));
  NOR2X1 G161 (.A1(W2959), .A2(W1107), .ZN(W3111));
  NOR2X1 G162 (.A1(W709), .A2(W2823), .ZN(W3113));
  NOR2X1 G163 (.A1(I665), .A2(W2352), .ZN(W3117));
  NOR2X1 G164 (.A1(W2162), .A2(W2221), .ZN(W3118));
  NOR2X1 G165 (.A1(I92), .A2(W1531), .ZN(W3119));
  NOR2X1 G166 (.A1(W1649), .A2(I622), .ZN(W3122));
  NOR2X1 G167 (.A1(I126), .A2(W1358), .ZN(W3093));
  NOR2X1 G168 (.A1(W2347), .A2(W1061), .ZN(O372));
  NOR2X1 G169 (.A1(W92), .A2(W765), .ZN(O373));
  NOR2X1 G170 (.A1(W1731), .A2(W502), .ZN(W3134));
  NOR2X1 G171 (.A1(I582), .A2(W527), .ZN(W3135));
  NOR2X1 G172 (.A1(W385), .A2(W92), .ZN(O376));
  NOR2X1 G173 (.A1(I408), .A2(I659), .ZN(W3141));
  NOR2X1 G174 (.A1(W311), .A2(W2328), .ZN(W3142));
  NOR2X1 G175 (.A1(W2871), .A2(I347), .ZN(O378));
  NOR2X1 G176 (.A1(W2950), .A2(W2574), .ZN(O381));
  NOR2X1 G177 (.A1(W769), .A2(I44), .ZN(O384));
  NOR2X1 G178 (.A1(W2624), .A2(I98), .ZN(W3154));
  NOR2X1 G179 (.A1(W2833), .A2(W810), .ZN(W3171));
  NOR2X1 G180 (.A1(I8), .A2(I104), .ZN(W3062));
  NOR2X1 G181 (.A1(W1120), .A2(W128), .ZN(W3027));
  NOR2X1 G182 (.A1(I428), .A2(I75), .ZN(W3029));
  NOR2X1 G183 (.A1(I817), .A2(I371), .ZN(W3030));
  NOR2X1 G184 (.A1(I732), .A2(W284), .ZN(O347));
  NOR2X1 G185 (.A1(W1992), .A2(W1886), .ZN(O348));
  NOR2X1 G186 (.A1(I772), .A2(W485), .ZN(O349));
  NOR2X1 G187 (.A1(W1870), .A2(W1947), .ZN(W3036));
  NOR2X1 G188 (.A1(W2535), .A2(W1318), .ZN(W3041));
  NOR2X1 G189 (.A1(W2463), .A2(W1760), .ZN(W3047));
  NOR2X1 G190 (.A1(W638), .A2(W2117), .ZN(O352));
  NOR2X1 G191 (.A1(W560), .A2(W520), .ZN(O353));
  NOR2X1 G192 (.A1(I82), .A2(W1870), .ZN(W3056));
  NOR2X1 G193 (.A1(W2181), .A2(W1376), .ZN(O472));
  NOR2X1 G194 (.A1(W343), .A2(W894), .ZN(W3063));
  NOR2X1 G195 (.A1(W2624), .A2(W920), .ZN(W3064));
  NOR2X1 G196 (.A1(W3016), .A2(W28), .ZN(O355));
  NOR2X1 G197 (.A1(W1742), .A2(W1865), .ZN(W3067));
  NOR2X1 G198 (.A1(W2169), .A2(I303), .ZN(W3070));
  NOR2X1 G199 (.A1(W2724), .A2(W86), .ZN(W3071));
  NOR2X1 G200 (.A1(I524), .A2(W1756), .ZN(W3078));
  NOR2X1 G201 (.A1(W1346), .A2(W959), .ZN(W3081));
  NOR2X1 G202 (.A1(W2177), .A2(W1630), .ZN(W3084));
  NOR2X1 G203 (.A1(I284), .A2(W2759), .ZN(W3088));
  NOR2X1 G204 (.A1(W2498), .A2(W904), .ZN(W3090));
  NOR2X1 G205 (.A1(I521), .A2(W1023), .ZN(O644));
  NOR2X1 G206 (.A1(W346), .A2(W3024), .ZN(W3880));
  NOR2X1 G207 (.A1(W764), .A2(W2995), .ZN(W3891));
  NOR2X1 G208 (.A1(W971), .A2(W240), .ZN(O636));
  NOR2X1 G209 (.A1(W201), .A2(W3464), .ZN(O638));
  NOR2X1 G210 (.A1(W3810), .A2(W592), .ZN(W3901));
  NOR2X1 G211 (.A1(W812), .A2(W2263), .ZN(W3902));
  NOR2X1 G212 (.A1(W3278), .A2(W292), .ZN(O639));
  NOR2X1 G213 (.A1(W1090), .A2(I684), .ZN(O641));
  NOR2X1 G214 (.A1(W705), .A2(W2964), .ZN(W3910));
  NOR2X1 G215 (.A1(W736), .A2(W1441), .ZN(W3914));
  NOR2X1 G216 (.A1(W2620), .A2(W345), .ZN(W3917));
  NOR2X1 G217 (.A1(W1551), .A2(W1968), .ZN(W3918));
  NOR2X1 G218 (.A1(W3054), .A2(W3792), .ZN(W3877));
  NOR2X1 G219 (.A1(W2441), .A2(W158), .ZN(O648));
  NOR2X1 G220 (.A1(W1604), .A2(W2777), .ZN(O649));
  NOR2X1 G221 (.A1(W3549), .A2(W2607), .ZN(W3929));
  NOR2X1 G222 (.A1(W237), .A2(W658), .ZN(O651));
  NOR2X1 G223 (.A1(W3255), .A2(W492), .ZN(W3932));
  NOR2X1 G224 (.A1(W3580), .A2(W811), .ZN(W3933));
  NOR2X1 G225 (.A1(W3361), .A2(W632), .ZN(O653));
  NOR2X1 G226 (.A1(W2796), .A2(W1343), .ZN(O655));
  NOR2X1 G227 (.A1(W2712), .A2(W1730), .ZN(O656));
  NOR2X1 G228 (.A1(W2992), .A2(W2294), .ZN(W3945));
  NOR2X1 G229 (.A1(W3298), .A2(W1462), .ZN(W3946));
  NOR2X1 G230 (.A1(W2287), .A2(W522), .ZN(W3947));
  NOR2X1 G231 (.A1(I676), .A2(W163), .ZN(O610));
  NOR2X1 G232 (.A1(W709), .A2(W3413), .ZN(W3813));
  NOR2X1 G233 (.A1(I490), .A2(W525), .ZN(W3816));
  NOR2X1 G234 (.A1(W2949), .A2(W2584), .ZN(O602));
  NOR2X1 G235 (.A1(W2905), .A2(W20), .ZN(W3820));
  NOR2X1 G236 (.A1(I385), .A2(W1878), .ZN(O603));
  NOR2X1 G237 (.A1(W3170), .A2(W3110), .ZN(W3826));
  NOR2X1 G238 (.A1(I760), .A2(W1444), .ZN(W3827));
  NOR2X1 G239 (.A1(W3374), .A2(W870), .ZN(W3830));
  NOR2X1 G240 (.A1(W1848), .A2(W30), .ZN(W3831));
  NOR2X1 G241 (.A1(W3069), .A2(W1830), .ZN(W3832));
  NOR2X1 G242 (.A1(W3438), .A2(W3690), .ZN(O609));
  NOR2X1 G243 (.A1(W1850), .A2(W3625), .ZN(W3838));
  NOR2X1 G244 (.A1(I811), .A2(W2969), .ZN(O662));
  NOR2X1 G245 (.A1(W3523), .A2(W2032), .ZN(W3844));
  NOR2X1 G246 (.A1(W2116), .A2(W3759), .ZN(O612));
  NOR2X1 G247 (.A1(I776), .A2(W141), .ZN(O614));
  NOR2X1 G248 (.A1(W3210), .A2(W1860), .ZN(O616));
  NOR2X1 G249 (.A1(W2026), .A2(W2692), .ZN(O621));
  NOR2X1 G250 (.A1(W2023), .A2(W3658), .ZN(O622));
  NOR2X1 G251 (.A1(W2838), .A2(W2040), .ZN(W3862));
  NOR2X1 G252 (.A1(W1799), .A2(W1029), .ZN(W3863));
  NOR2X1 G253 (.A1(W637), .A2(W2934), .ZN(O624));
  NOR2X1 G254 (.A1(W3286), .A2(W159), .ZN(W3865));
  NOR2X1 G255 (.A1(W1922), .A2(W605), .ZN(W3870));
  NOR2X1 G256 (.A1(W371), .A2(W1233), .ZN(O629));
  NOR2X1 G257 (.A1(W960), .A2(W4061), .ZN(W4064));
  NOR2X1 G258 (.A1(W925), .A2(W1822), .ZN(O697));
  NOR2X1 G259 (.A1(W3075), .A2(I389), .ZN(W4036));
  NOR2X1 G260 (.A1(W1555), .A2(W3333), .ZN(O702));
  NOR2X1 G261 (.A1(W3731), .A2(W126), .ZN(O703));
  NOR2X1 G262 (.A1(W16), .A2(W2750), .ZN(O704));
  NOR2X1 G263 (.A1(W3239), .A2(I222), .ZN(O705));
  NOR2X1 G264 (.A1(W1423), .A2(W2425), .ZN(W4047));
  NOR2X1 G265 (.A1(W1736), .A2(W2361), .ZN(O708));
  NOR2X1 G266 (.A1(I693), .A2(W2782), .ZN(W4054));
  NOR2X1 G267 (.A1(W1497), .A2(W7), .ZN(O710));
  NOR2X1 G268 (.A1(W3409), .A2(W697), .ZN(O716));
  NOR2X1 G269 (.A1(W857), .A2(W2005), .ZN(W4063));
  NOR2X1 G270 (.A1(W568), .A2(W2469), .ZN(W4025));
  NOR2X1 G271 (.A1(W693), .A2(W2714), .ZN(O717));
  NOR2X1 G272 (.A1(W1805), .A2(W2936), .ZN(O719));
  NOR2X1 G273 (.A1(W2054), .A2(W3336), .ZN(O722));
  NOR2X1 G274 (.A1(I925), .A2(W573), .ZN(O723));
  NOR2X1 G275 (.A1(I447), .A2(I839), .ZN(O724));
  NOR2X1 G276 (.A1(W1535), .A2(W610), .ZN(W4078));
  NOR2X1 G277 (.A1(W296), .A2(W3950), .ZN(W4081));
  NOR2X1 G278 (.A1(W1937), .A2(W3160), .ZN(O725));
  NOR2X1 G279 (.A1(W3), .A2(I420), .ZN(W4084));
  NOR2X1 G280 (.A1(W506), .A2(W3638), .ZN(O726));
  NOR2X1 G281 (.A1(W356), .A2(I481), .ZN(O727));
  NOR2X1 G282 (.A1(W1024), .A2(W588), .ZN(O729));
  NOR2X1 G283 (.A1(W1256), .A2(W2369), .ZN(O678));
  NOR2X1 G284 (.A1(W2086), .A2(W3054), .ZN(O667));
  NOR2X1 G285 (.A1(W454), .A2(I898), .ZN(W3960));
  NOR2X1 G286 (.A1(W362), .A2(W2699), .ZN(W3963));
  NOR2X1 G287 (.A1(W2474), .A2(W1183), .ZN(W3966));
  NOR2X1 G288 (.A1(W3344), .A2(I28), .ZN(W3968));
  NOR2X1 G289 (.A1(W3704), .A2(W1295), .ZN(O671));
  NOR2X1 G290 (.A1(W3749), .A2(W2234), .ZN(O672));
  NOR2X1 G291 (.A1(W2750), .A2(I518), .ZN(O673));
  NOR2X1 G292 (.A1(W1297), .A2(W3067), .ZN(W3974));
  NOR2X1 G293 (.A1(W985), .A2(W2188), .ZN(O674));
  NOR2X1 G294 (.A1(W3059), .A2(W3588), .ZN(W3979));
  NOR2X1 G295 (.A1(I235), .A2(W3601), .ZN(W3980));
  NOR2X1 G296 (.A1(W3689), .A2(W2597), .ZN(W3812));
  NOR2X1 G297 (.A1(W3791), .A2(W3874), .ZN(O679));
  NOR2X1 G298 (.A1(I495), .A2(W3183), .ZN(O681));
  NOR2X1 G299 (.A1(W1113), .A2(W730), .ZN(W3991));
  NOR2X1 G300 (.A1(W358), .A2(W509), .ZN(O686));
  NOR2X1 G301 (.A1(W3897), .A2(W1096), .ZN(O688));
  NOR2X1 G302 (.A1(W1782), .A2(I665), .ZN(O689));
  NOR2X1 G303 (.A1(W3554), .A2(W3302), .ZN(W4007));
  NOR2X1 G304 (.A1(W1527), .A2(W2781), .ZN(W4008));
  NOR2X1 G305 (.A1(W1290), .A2(I292), .ZN(W4012));
  NOR2X1 G306 (.A1(W1718), .A2(I913), .ZN(O691));
  NOR2X1 G307 (.A1(I870), .A2(I879), .ZN(O694));
  NOR2X1 G308 (.A1(W2730), .A2(W105), .ZN(O510));
  NOR2X1 G309 (.A1(W1807), .A2(W2354), .ZN(O500));
  NOR2X1 G310 (.A1(W3076), .A2(W2635), .ZN(W3549));
  NOR2X1 G311 (.A1(W1129), .A2(W517), .ZN(W3554));
  NOR2X1 G312 (.A1(W2513), .A2(W3415), .ZN(W3556));
  NOR2X1 G313 (.A1(W640), .A2(I138), .ZN(W3560));
  NOR2X1 G314 (.A1(W1586), .A2(W1667), .ZN(O506));
  NOR2X1 G315 (.A1(I289), .A2(W1103), .ZN(O507));
  NOR2X1 G316 (.A1(W1081), .A2(W2086), .ZN(W3575));
  NOR2X1 G317 (.A1(W2952), .A2(W460), .ZN(W3577));
  NOR2X1 G318 (.A1(W3199), .A2(W1776), .ZN(W3580));
  NOR2X1 G319 (.A1(W877), .A2(W2412), .ZN(W3582));
  NOR2X1 G320 (.A1(W616), .A2(W2273), .ZN(W3583));
  NOR2X1 G321 (.A1(W3414), .A2(W55), .ZN(W3544));
  NOR2X1 G322 (.A1(W1666), .A2(W2523), .ZN(O512));
  NOR2X1 G323 (.A1(I822), .A2(W731), .ZN(O514));
  NOR2X1 G324 (.A1(W2183), .A2(W1748), .ZN(O515));
  NOR2X1 G325 (.A1(W1552), .A2(I459), .ZN(W3594));
  NOR2X1 G326 (.A1(W3198), .A2(W777), .ZN(W3599));
  NOR2X1 G327 (.A1(W1729), .A2(W1114), .ZN(W3606));
  NOR2X1 G328 (.A1(W1843), .A2(W1845), .ZN(W3609));
  NOR2X1 G329 (.A1(W3196), .A2(W1477), .ZN(O522));
  NOR2X1 G330 (.A1(W1206), .A2(W510), .ZN(O524));
  NOR2X1 G331 (.A1(I785), .A2(W206), .ZN(O528));
  NOR2X1 G332 (.A1(W875), .A2(W266), .ZN(W3623));
  NOR2X1 G333 (.A1(W1425), .A2(W14), .ZN(W3624));
  NOR2X1 G334 (.A1(W1839), .A2(I270), .ZN(W3503));
  NOR2X1 G335 (.A1(W3152), .A2(W2289), .ZN(O473));
  NOR2X1 G336 (.A1(W2577), .A2(W523), .ZN(W3461));
  NOR2X1 G337 (.A1(I462), .A2(W2526), .ZN(W3464));
  NOR2X1 G338 (.A1(I820), .A2(W843), .ZN(W3472));
  NOR2X1 G339 (.A1(W1599), .A2(W93), .ZN(W3473));
  NOR2X1 G340 (.A1(W2873), .A2(W382), .ZN(W3480));
  NOR2X1 G341 (.A1(W2730), .A2(W3093), .ZN(O485));
  NOR2X1 G342 (.A1(W2322), .A2(W426), .ZN(W3489));
  NOR2X1 G343 (.A1(W253), .A2(W2622), .ZN(W3490));
  NOR2X1 G344 (.A1(W799), .A2(W1747), .ZN(O487));
  NOR2X1 G345 (.A1(W1755), .A2(W497), .ZN(W3496));
  NOR2X1 G346 (.A1(W1459), .A2(W2752), .ZN(O489));
  NOR2X1 G347 (.A1(I198), .A2(W261), .ZN(O530));
  NOR2X1 G348 (.A1(W713), .A2(I767), .ZN(W3505));
  NOR2X1 G349 (.A1(W3329), .A2(W2388), .ZN(W3509));
  NOR2X1 G350 (.A1(W1834), .A2(W1269), .ZN(W3511));
  NOR2X1 G351 (.A1(W2942), .A2(W2731), .ZN(W3519));
  NOR2X1 G352 (.A1(I213), .A2(W3130), .ZN(W3523));
  NOR2X1 G353 (.A1(W2281), .A2(W2086), .ZN(W3525));
  NOR2X1 G354 (.A1(W2993), .A2(W1428), .ZN(W3528));
  NOR2X1 G355 (.A1(I637), .A2(W1203), .ZN(W3533));
  NOR2X1 G356 (.A1(I471), .A2(W645), .ZN(W3538));
  NOR2X1 G357 (.A1(W98), .A2(W2246), .ZN(W3542));
  NOR2X1 G358 (.A1(W926), .A2(W1904), .ZN(W3543));
  NOR2X1 G359 (.A1(W1314), .A2(W3688), .ZN(O581));
  NOR2X1 G360 (.A1(W788), .A2(W1514), .ZN(W3722));
  NOR2X1 G361 (.A1(I234), .A2(I203), .ZN(O566));
  NOR2X1 G362 (.A1(W1191), .A2(I444), .ZN(O568));
  NOR2X1 G363 (.A1(I552), .A2(W2377), .ZN(W3734));
  NOR2X1 G364 (.A1(W179), .A2(W1133), .ZN(W3735));
  NOR2X1 G365 (.A1(W2256), .A2(I911), .ZN(W3736));
  NOR2X1 G366 (.A1(W3629), .A2(W3179), .ZN(W3744));
  NOR2X1 G367 (.A1(W3654), .A2(W2871), .ZN(W3749));
  NOR2X1 G368 (.A1(W2994), .A2(W3315), .ZN(W3750));
  NOR2X1 G369 (.A1(W2118), .A2(W2220), .ZN(O575));
  NOR2X1 G370 (.A1(W1823), .A2(W1827), .ZN(O576));
  NOR2X1 G371 (.A1(I417), .A2(W1203), .ZN(O579));
  NOR2X1 G372 (.A1(W1178), .A2(W3355), .ZN(W3709));
  NOR2X1 G373 (.A1(W2818), .A2(W2111), .ZN(W3761));
  NOR2X1 G374 (.A1(W1009), .A2(W3699), .ZN(W3764));
  NOR2X1 G375 (.A1(I194), .A2(W804), .ZN(O583));
  NOR2X1 G376 (.A1(W659), .A2(W2687), .ZN(W3769));
  NOR2X1 G377 (.A1(W1103), .A2(W2329), .ZN(W3780));
  NOR2X1 G378 (.A1(W1509), .A2(I626), .ZN(O589));
  NOR2X1 G379 (.A1(W604), .A2(W3386), .ZN(O590));
  NOR2X1 G380 (.A1(I799), .A2(W3540), .ZN(O593));
  NOR2X1 G381 (.A1(W2347), .A2(W3720), .ZN(W3793));
  NOR2X1 G382 (.A1(W2129), .A2(W2157), .ZN(O599));
  NOR2X1 G383 (.A1(W3334), .A2(W3765), .ZN(O600));
  NOR2X1 G384 (.A1(W2332), .A2(W1381), .ZN(W3811));
  NOR2X1 G385 (.A1(W3378), .A2(W3346), .ZN(O550));
  NOR2X1 G386 (.A1(I527), .A2(W1468), .ZN(O532));
  NOR2X1 G387 (.A1(W2388), .A2(W1514), .ZN(O533));
  NOR2X1 G388 (.A1(W2849), .A2(W1032), .ZN(O535));
  NOR2X1 G389 (.A1(W2578), .A2(W2395), .ZN(W3636));
  NOR2X1 G390 (.A1(W1505), .A2(W1016), .ZN(W3639));
  NOR2X1 G391 (.A1(I110), .A2(W2100), .ZN(W3642));
  NOR2X1 G392 (.A1(W2174), .A2(W953), .ZN(O542));
  NOR2X1 G393 (.A1(W1521), .A2(W2193), .ZN(W3659));
  NOR2X1 G394 (.A1(W230), .A2(W638), .ZN(W3661));
  NOR2X1 G395 (.A1(W1634), .A2(W137), .ZN(W3664));
  NOR2X1 G396 (.A1(W2066), .A2(W929), .ZN(O547));
  NOR2X1 G397 (.A1(I781), .A2(W2228), .ZN(W3672));
  NOR2X1 G398 (.A1(W2041), .A2(W1878), .ZN(W2874));
  NOR2X1 G399 (.A1(W738), .A2(W3535), .ZN(W3683));
  NOR2X1 G400 (.A1(W2056), .A2(W1132), .ZN(W3687));
  NOR2X1 G401 (.A1(W2233), .A2(W2401), .ZN(W3690));
  NOR2X1 G402 (.A1(I226), .A2(W3260), .ZN(W3691));
  NOR2X1 G403 (.A1(W2419), .A2(W2298), .ZN(O557));
  NOR2X1 G404 (.A1(W2059), .A2(W2842), .ZN(W3695));
  NOR2X1 G405 (.A1(I433), .A2(W910), .ZN(W3697));
  NOR2X1 G406 (.A1(I420), .A2(W2392), .ZN(W3698));
  NOR2X1 G407 (.A1(I6), .A2(W2119), .ZN(O560));
  NOR2X1 G408 (.A1(I348), .A2(W2286), .ZN(W3705));
  NOR2X1 G409 (.A1(W3664), .A2(W967), .ZN(W3708));
  NOR2X1 G410 (.A1(W509), .A2(W582), .ZN(W2047));
  NOR2X1 G411 (.A1(W431), .A2(W1451), .ZN(W1999));
  NOR2X1 G412 (.A1(W1953), .A2(W35), .ZN(W2000));
  NOR2X1 G413 (.A1(W1068), .A2(W450), .ZN(W2002));
  NOR2X1 G414 (.A1(W1150), .A2(I479), .ZN(W2006));
  NOR2X1 G415 (.A1(W216), .A2(I288), .ZN(W2014));
  NOR2X1 G416 (.A1(I66), .A2(W1563), .ZN(O137));
  NOR2X1 G417 (.A1(I262), .A2(W117), .ZN(W2029));
  NOR2X1 G418 (.A1(W747), .A2(W632), .ZN(O139));
  NOR2X1 G419 (.A1(W1155), .A2(I548), .ZN(W2040));
  NOR2X1 G420 (.A1(W864), .A2(W1324), .ZN(O140));
  NOR2X1 G421 (.A1(W1282), .A2(I175), .ZN(W2044));
  NOR2X1 G422 (.A1(I488), .A2(W1070), .ZN(W2046));
  NOR2X1 G423 (.A1(I909), .A2(W601), .ZN(O135));
  NOR2X1 G424 (.A1(W1167), .A2(I648), .ZN(W2048));
  NOR2X1 G425 (.A1(I9), .A2(W1415), .ZN(W2051));
  NOR2X1 G426 (.A1(W1949), .A2(W1301), .ZN(W2054));
  NOR2X1 G427 (.A1(W1952), .A2(W1126), .ZN(W2055));
  NOR2X1 G428 (.A1(W972), .A2(W274), .ZN(W2057));
  NOR2X1 G429 (.A1(W218), .A2(W155), .ZN(W2058));
  NOR2X1 G430 (.A1(W755), .A2(W802), .ZN(W2062));
  NOR2X1 G431 (.A1(W1679), .A2(I270), .ZN(W2063));
  NOR2X1 G432 (.A1(W1856), .A2(W1075), .ZN(O143));
  NOR2X1 G433 (.A1(W1224), .A2(W819), .ZN(W2068));
  NOR2X1 G434 (.A1(I436), .A2(W1654), .ZN(W2070));
  NOR2X1 G435 (.A1(I857), .A2(I339), .ZN(O145));
  NOR2X1 G436 (.A1(I330), .A2(W84), .ZN(W1963));
  NOR2X1 G437 (.A1(W22), .A2(I720), .ZN(W1928));
  NOR2X1 G438 (.A1(W922), .A2(I654), .ZN(W1931));
  NOR2X1 G439 (.A1(W822), .A2(W270), .ZN(W1932));
  NOR2X1 G440 (.A1(W987), .A2(W1630), .ZN(W1938));
  NOR2X1 G441 (.A1(W761), .A2(W478), .ZN(W1942));
  NOR2X1 G442 (.A1(I634), .A2(I524), .ZN(W1944));
  NOR2X1 G443 (.A1(W1783), .A2(W1748), .ZN(W1945));
  NOR2X1 G444 (.A1(W1490), .A2(I44), .ZN(W1947));
  NOR2X1 G445 (.A1(I256), .A2(W655), .ZN(W1949));
  NOR2X1 G446 (.A1(W1776), .A2(W111), .ZN(W1950));
  NOR2X1 G447 (.A1(I849), .A2(I416), .ZN(W1955));
  NOR2X1 G448 (.A1(W1949), .A2(W660), .ZN(W1956));
  NOR2X1 G449 (.A1(W2072), .A2(W334), .ZN(W2076));
  NOR2X1 G450 (.A1(W671), .A2(W194), .ZN(W1966));
  NOR2X1 G451 (.A1(I212), .A2(W1256), .ZN(W1968));
  NOR2X1 G452 (.A1(W1631), .A2(W1929), .ZN(W1969));
  NOR2X1 G453 (.A1(I600), .A2(W1244), .ZN(W1970));
  NOR2X1 G454 (.A1(I21), .A2(W1207), .ZN(O133));
  NOR2X1 G455 (.A1(W1546), .A2(W704), .ZN(W1974));
  NOR2X1 G456 (.A1(I832), .A2(W1849), .ZN(O134));
  NOR2X1 G457 (.A1(W1782), .A2(W1774), .ZN(W1980));
  NOR2X1 G458 (.A1(W831), .A2(I130), .ZN(W1988));
  NOR2X1 G459 (.A1(W619), .A2(W1959), .ZN(W1990));
  NOR2X1 G460 (.A1(W1811), .A2(W949), .ZN(W1991));
  NOR2X1 G461 (.A1(W133), .A2(W61), .ZN(W1993));
  NOR2X1 G462 (.A1(W556), .A2(W1080), .ZN(W2172));
  NOR2X1 G463 (.A1(W791), .A2(W1728), .ZN(O161));
  NOR2X1 G464 (.A1(W1054), .A2(I232), .ZN(W2147));
  NOR2X1 G465 (.A1(I446), .A2(I928), .ZN(W2150));
  NOR2X1 G466 (.A1(W1259), .A2(W105), .ZN(W2155));
  NOR2X1 G467 (.A1(I52), .A2(W1639), .ZN(W2158));
  NOR2X1 G468 (.A1(I576), .A2(W2053), .ZN(W2159));
  NOR2X1 G469 (.A1(W26), .A2(W1907), .ZN(W2160));
  NOR2X1 G470 (.A1(W213), .A2(W1148), .ZN(W2161));
  NOR2X1 G471 (.A1(I940), .A2(W528), .ZN(W2162));
  NOR2X1 G472 (.A1(I522), .A2(W1190), .ZN(W2164));
  NOR2X1 G473 (.A1(W73), .A2(I468), .ZN(W2168));
  NOR2X1 G474 (.A1(W502), .A2(I572), .ZN(W2169));
  NOR2X1 G475 (.A1(W1456), .A2(W1318), .ZN(O160));
  NOR2X1 G476 (.A1(I829), .A2(W1006), .ZN(W2178));
  NOR2X1 G477 (.A1(I612), .A2(I765), .ZN(W2180));
  NOR2X1 G478 (.A1(I392), .A2(W542), .ZN(W2185));
  NOR2X1 G479 (.A1(I40), .A2(W39), .ZN(O169));
  NOR2X1 G480 (.A1(W2126), .A2(I828), .ZN(W2188));
  NOR2X1 G481 (.A1(W1748), .A2(W1855), .ZN(W2190));
  NOR2X1 G482 (.A1(I491), .A2(W375), .ZN(W2192));
  NOR2X1 G483 (.A1(W1295), .A2(I921), .ZN(W2193));
  NOR2X1 G484 (.A1(W305), .A2(W2080), .ZN(W2195));
  NOR2X1 G485 (.A1(W1579), .A2(W158), .ZN(O170));
  NOR2X1 G486 (.A1(W1240), .A2(W319), .ZN(O173));
  NOR2X1 G487 (.A1(W1240), .A2(W218), .ZN(O175));
  NOR2X1 G488 (.A1(I137), .A2(W1695), .ZN(O155));
  NOR2X1 G489 (.A1(W1209), .A2(I905), .ZN(W2078));
  NOR2X1 G490 (.A1(W152), .A2(I468), .ZN(W2080));
  NOR2X1 G491 (.A1(I6), .A2(I241), .ZN(W2082));
  NOR2X1 G492 (.A1(W870), .A2(W889), .ZN(O146));
  NOR2X1 G493 (.A1(W1841), .A2(W1815), .ZN(W2085));
  NOR2X1 G494 (.A1(I278), .A2(W366), .ZN(W2088));
  NOR2X1 G495 (.A1(I725), .A2(W760), .ZN(W2089));
  NOR2X1 G496 (.A1(W1680), .A2(W674), .ZN(W2093));
  NOR2X1 G497 (.A1(W1737), .A2(W859), .ZN(O150));
  NOR2X1 G498 (.A1(I508), .A2(W1695), .ZN(O151));
  NOR2X1 G499 (.A1(I460), .A2(W1434), .ZN(W2099));
  NOR2X1 G500 (.A1(W71), .A2(W229), .ZN(W2106));
  NOR2X1 G501 (.A1(W1324), .A2(W1690), .ZN(W1922));
  NOR2X1 G502 (.A1(I641), .A2(W688), .ZN(W2111));
  NOR2X1 G503 (.A1(W1009), .A2(W1884), .ZN(W2116));
  NOR2X1 G504 (.A1(W792), .A2(W173), .ZN(W2122));
  NOR2X1 G505 (.A1(W1750), .A2(W1729), .ZN(W2128));
  NOR2X1 G506 (.A1(W1819), .A2(W698), .ZN(W2130));
  NOR2X1 G507 (.A1(W2018), .A2(W132), .ZN(W2131));
  NOR2X1 G508 (.A1(W273), .A2(W748), .ZN(W2133));
  NOR2X1 G509 (.A1(I452), .A2(I870), .ZN(O159));
  NOR2X1 G510 (.A1(I868), .A2(W253), .ZN(W2138));
  NOR2X1 G511 (.A1(W421), .A2(I122), .ZN(W2140));
  NOR2X1 G512 (.A1(I539), .A2(W1949), .ZN(W2141));
  NOR2X1 G513 (.A1(W617), .A2(W761), .ZN(W1735));
  NOR2X1 G514 (.A1(W1236), .A2(W1310), .ZN(W1707));
  NOR2X1 G515 (.A1(W1697), .A2(W813), .ZN(W1709));
  NOR2X1 G516 (.A1(W1594), .A2(W1383), .ZN(O97));
  NOR2X1 G517 (.A1(I730), .A2(I614), .ZN(W1711));
  NOR2X1 G518 (.A1(W965), .A2(W352), .ZN(O98));
  NOR2X1 G519 (.A1(W1029), .A2(I648), .ZN(O99));
  NOR2X1 G520 (.A1(I953), .A2(I469), .ZN(W1720));
  NOR2X1 G521 (.A1(I927), .A2(W1444), .ZN(W1721));
  NOR2X1 G522 (.A1(I745), .A2(I629), .ZN(W1722));
  NOR2X1 G523 (.A1(W74), .A2(W368), .ZN(O100));
  NOR2X1 G524 (.A1(W637), .A2(I684), .ZN(O101));
  NOR2X1 G525 (.A1(W1580), .A2(W1099), .ZN(W1731));
  NOR2X1 G526 (.A1(W1423), .A2(I12), .ZN(W1705));
  NOR2X1 G527 (.A1(W1111), .A2(W875), .ZN(W1737));
  NOR2X1 G528 (.A1(W346), .A2(I285), .ZN(W1740));
  NOR2X1 G529 (.A1(I102), .A2(W104), .ZN(W1741));
  NOR2X1 G530 (.A1(W937), .A2(I618), .ZN(W1743));
  NOR2X1 G531 (.A1(W566), .A2(I677), .ZN(W1744));
  NOR2X1 G532 (.A1(I879), .A2(W929), .ZN(W1745));
  NOR2X1 G533 (.A1(W574), .A2(I594), .ZN(W1746));
  NOR2X1 G534 (.A1(I50), .A2(W1307), .ZN(W1748));
  NOR2X1 G535 (.A1(I413), .A2(W692), .ZN(W1749));
  NOR2X1 G536 (.A1(W100), .A2(I118), .ZN(W1752));
  NOR2X1 G537 (.A1(W1519), .A2(W1462), .ZN(W1755));
  NOR2X1 G538 (.A1(W1474), .A2(W970), .ZN(W1756));
  NOR2X1 G539 (.A1(W1318), .A2(I781), .ZN(W1673));
  NOR2X1 G540 (.A1(W752), .A2(W1400), .ZN(W1640));
  NOR2X1 G541 (.A1(W1457), .A2(W853), .ZN(W1642));
  NOR2X1 G542 (.A1(I219), .A2(I737), .ZN(W1643));
  NOR2X1 G543 (.A1(W95), .A2(W1329), .ZN(W1645));
  NOR2X1 G544 (.A1(I934), .A2(W1516), .ZN(W1648));
  NOR2X1 G545 (.A1(W1516), .A2(W1067), .ZN(W1651));
  NOR2X1 G546 (.A1(W197), .A2(W1295), .ZN(W1652));
  NOR2X1 G547 (.A1(W146), .A2(W689), .ZN(W1659));
  NOR2X1 G548 (.A1(W210), .A2(W661), .ZN(W1661));
  NOR2X1 G549 (.A1(I927), .A2(W1504), .ZN(W1665));
  NOR2X1 G550 (.A1(I230), .A2(W1602), .ZN(W1668));
  NOR2X1 G551 (.A1(W148), .A2(W931), .ZN(W1672));
  NOR2X1 G552 (.A1(W1226), .A2(W492), .ZN(W1761));
  NOR2X1 G553 (.A1(W258), .A2(I318), .ZN(W1680));
  NOR2X1 G554 (.A1(I928), .A2(I743), .ZN(W1689));
  NOR2X1 G555 (.A1(W1418), .A2(I163), .ZN(W1691));
  NOR2X1 G556 (.A1(I338), .A2(W605), .ZN(W1692));
  NOR2X1 G557 (.A1(W1258), .A2(I151), .ZN(W1693));
  NOR2X1 G558 (.A1(W1211), .A2(W679), .ZN(W1695));
  NOR2X1 G559 (.A1(I371), .A2(W1541), .ZN(W1697));
  NOR2X1 G560 (.A1(W768), .A2(W270), .ZN(O95));
  NOR2X1 G561 (.A1(I707), .A2(I892), .ZN(W1699));
  NOR2X1 G562 (.A1(W1291), .A2(W486), .ZN(W1701));
  NOR2X1 G563 (.A1(I564), .A2(I181), .ZN(W1702));
  NOR2X1 G564 (.A1(W870), .A2(W1078), .ZN(W1884));
  NOR2X1 G565 (.A1(W1701), .A2(W562), .ZN(W1845));
  NOR2X1 G566 (.A1(W1019), .A2(W955), .ZN(W1846));
  NOR2X1 G567 (.A1(W109), .A2(I968), .ZN(W1851));
  NOR2X1 G568 (.A1(W1635), .A2(W961), .ZN(W1853));
  NOR2X1 G569 (.A1(W697), .A2(W1216), .ZN(W1854));
  NOR2X1 G570 (.A1(W1075), .A2(W1326), .ZN(W1860));
  NOR2X1 G571 (.A1(I42), .A2(W598), .ZN(W1865));
  NOR2X1 G572 (.A1(I542), .A2(I741), .ZN(W1866));
  NOR2X1 G573 (.A1(W1191), .A2(I213), .ZN(O117));
  NOR2X1 G574 (.A1(I243), .A2(I894), .ZN(W1873));
  NOR2X1 G575 (.A1(W297), .A2(I103), .ZN(W1876));
  NOR2X1 G576 (.A1(W1461), .A2(I895), .ZN(W1881));
  NOR2X1 G577 (.A1(W1005), .A2(I511), .ZN(W1844));
  NOR2X1 G578 (.A1(W1617), .A2(W11), .ZN(W1886));
  NOR2X1 G579 (.A1(W639), .A2(I20), .ZN(W1887));
  NOR2X1 G580 (.A1(W1327), .A2(W134), .ZN(O120));
  NOR2X1 G581 (.A1(W316), .A2(W1163), .ZN(W1890));
  NOR2X1 G582 (.A1(W1788), .A2(W1662), .ZN(W1895));
  NOR2X1 G583 (.A1(I124), .A2(W1189), .ZN(W1897));
  NOR2X1 G584 (.A1(W1589), .A2(I626), .ZN(O122));
  NOR2X1 G585 (.A1(W942), .A2(W1), .ZN(O123));
  NOR2X1 G586 (.A1(W184), .A2(W1688), .ZN(W1907));
  NOR2X1 G587 (.A1(W643), .A2(I542), .ZN(W1909));
  NOR2X1 G588 (.A1(W1166), .A2(W857), .ZN(W1916));
  NOR2X1 G589 (.A1(W90), .A2(W1451), .ZN(W1919));
  NOR2X1 G590 (.A1(W1697), .A2(W1257), .ZN(W1811));
  NOR2X1 G591 (.A1(W1086), .A2(W718), .ZN(W1762));
  NOR2X1 G592 (.A1(I328), .A2(I452), .ZN(W1763));
  NOR2X1 G593 (.A1(W839), .A2(I222), .ZN(W1764));
  NOR2X1 G594 (.A1(W1326), .A2(I23), .ZN(O104));
  NOR2X1 G595 (.A1(W34), .A2(I621), .ZN(W1779));
  NOR2X1 G596 (.A1(W1206), .A2(W151), .ZN(W1785));
  NOR2X1 G597 (.A1(W947), .A2(W475), .ZN(O107));
  NOR2X1 G598 (.A1(W741), .A2(W838), .ZN(W1789));
  NOR2X1 G599 (.A1(I655), .A2(W256), .ZN(W1797));
  NOR2X1 G600 (.A1(W430), .A2(W642), .ZN(W1801));
  NOR2X1 G601 (.A1(W567), .A2(W1074), .ZN(W1804));
  NOR2X1 G602 (.A1(W130), .A2(W1003), .ZN(O111));
  NOR2X1 G603 (.A1(I696), .A2(W1219), .ZN(W2214));
  NOR2X1 G604 (.A1(I833), .A2(W1382), .ZN(W1813));
  NOR2X1 G605 (.A1(W261), .A2(W938), .ZN(W1819));
  NOR2X1 G606 (.A1(W944), .A2(I290), .ZN(W1821));
  NOR2X1 G607 (.A1(W477), .A2(I228), .ZN(W1824));
  NOR2X1 G608 (.A1(W246), .A2(W1543), .ZN(W1825));
  NOR2X1 G609 (.A1(W283), .A2(W400), .ZN(O113));
  NOR2X1 G610 (.A1(W1588), .A2(W1023), .ZN(W1832));
  NOR2X1 G611 (.A1(W1334), .A2(I753), .ZN(W1834));
  NOR2X1 G612 (.A1(W1778), .A2(W1278), .ZN(W1835));
  NOR2X1 G613 (.A1(I153), .A2(W513), .ZN(W1841));
  NOR2X1 G614 (.A1(W91), .A2(W1563), .ZN(W1842));
  NOR2X1 G615 (.A1(W1927), .A2(W1863), .ZN(O259));
  NOR2X1 G616 (.A1(I748), .A2(W1424), .ZN(W2632));
  NOR2X1 G617 (.A1(I29), .A2(W2487), .ZN(O250));
  NOR2X1 G618 (.A1(W1702), .A2(W2089), .ZN(W2640));
  NOR2X1 G619 (.A1(W1630), .A2(W1636), .ZN(W2641));
  NOR2X1 G620 (.A1(W1346), .A2(W1941), .ZN(W2646));
  NOR2X1 G621 (.A1(W356), .A2(W12), .ZN(O252));
  NOR2X1 G622 (.A1(W1322), .A2(W2157), .ZN(O253));
  NOR2X1 G623 (.A1(W779), .A2(W967), .ZN(W2652));
  NOR2X1 G624 (.A1(W1878), .A2(W501), .ZN(O255));
  NOR2X1 G625 (.A1(W647), .A2(W1488), .ZN(W2659));
  NOR2X1 G626 (.A1(W1819), .A2(W2026), .ZN(W2660));
  NOR2X1 G627 (.A1(W2492), .A2(W2567), .ZN(O257));
  NOR2X1 G628 (.A1(I710), .A2(I62), .ZN(W2630));
  NOR2X1 G629 (.A1(W331), .A2(W2579), .ZN(W2674));
  NOR2X1 G630 (.A1(W1613), .A2(I684), .ZN(W2675));
  NOR2X1 G631 (.A1(W1205), .A2(W2263), .ZN(W2680));
  NOR2X1 G632 (.A1(W569), .A2(W488), .ZN(W2682));
  NOR2X1 G633 (.A1(W2434), .A2(I228), .ZN(O263));
  NOR2X1 G634 (.A1(W2496), .A2(W2660), .ZN(W2687));
  NOR2X1 G635 (.A1(W2070), .A2(W1094), .ZN(W2694));
  NOR2X1 G636 (.A1(W2033), .A2(W1448), .ZN(O268));
  NOR2X1 G637 (.A1(W668), .A2(I849), .ZN(W2703));
  NOR2X1 G638 (.A1(W73), .A2(W1963), .ZN(W2708));
  NOR2X1 G639 (.A1(W952), .A2(W429), .ZN(W2710));
  NOR2X1 G640 (.A1(W1852), .A2(I660), .ZN(W2714));
  NOR2X1 G641 (.A1(I257), .A2(I680), .ZN(W2584));
  NOR2X1 G642 (.A1(I556), .A2(I551), .ZN(O230));
  NOR2X1 G643 (.A1(I620), .A2(W240), .ZN(O232));
  NOR2X1 G644 (.A1(W832), .A2(W60), .ZN(W2556));
  NOR2X1 G645 (.A1(I882), .A2(W881), .ZN(W2562));
  NOR2X1 G646 (.A1(I953), .A2(I660), .ZN(W2567));
  NOR2X1 G647 (.A1(W1066), .A2(W2413), .ZN(W2571));
  NOR2X1 G648 (.A1(I550), .A2(W1246), .ZN(W2572));
  NOR2X1 G649 (.A1(W2170), .A2(W334), .ZN(W2573));
  NOR2X1 G650 (.A1(W1439), .A2(W663), .ZN(W2574));
  NOR2X1 G651 (.A1(W463), .A2(W1152), .ZN(W2575));
  NOR2X1 G652 (.A1(W65), .A2(W1251), .ZN(W2579));
  NOR2X1 G653 (.A1(W2277), .A2(W1629), .ZN(W2582));
  NOR2X1 G654 (.A1(I489), .A2(W1187), .ZN(W2716));
  NOR2X1 G655 (.A1(W1570), .A2(W2029), .ZN(W2588));
  NOR2X1 G656 (.A1(W2399), .A2(W752), .ZN(W2591));
  NOR2X1 G657 (.A1(W741), .A2(W940), .ZN(W2595));
  NOR2X1 G658 (.A1(W2265), .A2(W716), .ZN(W2599));
  NOR2X1 G659 (.A1(W2568), .A2(W286), .ZN(W2601));
  NOR2X1 G660 (.A1(W2526), .A2(W295), .ZN(O245));
  NOR2X1 G661 (.A1(I540), .A2(W648), .ZN(W2622));
  NOR2X1 G662 (.A1(W2146), .A2(I988), .ZN(W2624));
  NOR2X1 G663 (.A1(W470), .A2(I314), .ZN(W2625));
  NOR2X1 G664 (.A1(W2320), .A2(I976), .ZN(O248));
  NOR2X1 G665 (.A1(W1360), .A2(W1135), .ZN(O249));
  NOR2X1 G666 (.A1(W1836), .A2(I632), .ZN(W2829));
  NOR2X1 G667 (.A1(W2111), .A2(W1392), .ZN(W2804));
  NOR2X1 G668 (.A1(W2676), .A2(W137), .ZN(W2805));
  NOR2X1 G669 (.A1(W774), .A2(W2568), .ZN(W2807));
  NOR2X1 G670 (.A1(W2637), .A2(W672), .ZN(O291));
  NOR2X1 G671 (.A1(W1611), .A2(W2447), .ZN(O293));
  NOR2X1 G672 (.A1(I447), .A2(W198), .ZN(W2812));
  NOR2X1 G673 (.A1(W1685), .A2(W2328), .ZN(O294));
  NOR2X1 G674 (.A1(W357), .A2(W2781), .ZN(W2815));
  NOR2X1 G675 (.A1(W128), .A2(I936), .ZN(W2816));
  NOR2X1 G676 (.A1(W2814), .A2(W2276), .ZN(W2817));
  NOR2X1 G677 (.A1(W2653), .A2(W1587), .ZN(O295));
  NOR2X1 G678 (.A1(I110), .A2(W690), .ZN(O297));
  NOR2X1 G679 (.A1(I652), .A2(W1291), .ZN(W2801));
  NOR2X1 G680 (.A1(W618), .A2(W135), .ZN(W2834));
  NOR2X1 G681 (.A1(W741), .A2(W933), .ZN(O301));
  NOR2X1 G682 (.A1(W2255), .A2(W2357), .ZN(W2845));
  NOR2X1 G683 (.A1(I164), .A2(W757), .ZN(W2847));
  NOR2X1 G684 (.A1(W1338), .A2(W1688), .ZN(O305));
  NOR2X1 G685 (.A1(W1477), .A2(I252), .ZN(W2856));
  NOR2X1 G686 (.A1(W541), .A2(I990), .ZN(O309));
  NOR2X1 G687 (.A1(W799), .A2(I581), .ZN(W2859));
  NOR2X1 G688 (.A1(W579), .A2(W1279), .ZN(W2863));
  NOR2X1 G689 (.A1(W1917), .A2(W2642), .ZN(W2864));
  NOR2X1 G690 (.A1(W166), .A2(I347), .ZN(W2871));
  NOR2X1 G691 (.A1(I996), .A2(I987), .ZN(W2872));
  NOR2X1 G692 (.A1(W1912), .A2(W765), .ZN(W2751));
  NOR2X1 G693 (.A1(I61), .A2(W1455), .ZN(W2720));
  NOR2X1 G694 (.A1(W646), .A2(W2575), .ZN(W2721));
  NOR2X1 G695 (.A1(W1026), .A2(W2515), .ZN(W2729));
  NOR2X1 G696 (.A1(I797), .A2(W288), .ZN(W2730));
  NOR2X1 G697 (.A1(W2190), .A2(I975), .ZN(W2731));
  NOR2X1 G698 (.A1(W201), .A2(I799), .ZN(O273));
  NOR2X1 G699 (.A1(W1695), .A2(W2194), .ZN(W2736));
  NOR2X1 G700 (.A1(W2414), .A2(W1394), .ZN(W2737));
  NOR2X1 G701 (.A1(W724), .A2(W2496), .ZN(W2739));
  NOR2X1 G702 (.A1(W551), .A2(W2549), .ZN(O277));
  NOR2X1 G703 (.A1(I98), .A2(W2295), .ZN(O278));
  NOR2X1 G704 (.A1(I506), .A2(W1510), .ZN(W2749));
  NOR2X1 G705 (.A1(I248), .A2(W1303), .ZN(W2536));
  NOR2X1 G706 (.A1(W2683), .A2(W2304), .ZN(O280));
  NOR2X1 G707 (.A1(W1115), .A2(W2158), .ZN(W2758));
  NOR2X1 G708 (.A1(I175), .A2(W568), .ZN(W2759));
  NOR2X1 G709 (.A1(W539), .A2(W1573), .ZN(O284));
  NOR2X1 G710 (.A1(W522), .A2(W1789), .ZN(W2769));
  NOR2X1 G711 (.A1(W587), .A2(W1113), .ZN(W2774));
  NOR2X1 G712 (.A1(W1045), .A2(W1075), .ZN(W2777));
  NOR2X1 G713 (.A1(W1823), .A2(W2718), .ZN(W2781));
  NOR2X1 G714 (.A1(W5), .A2(W1321), .ZN(W2789));
  NOR2X1 G715 (.A1(W82), .A2(W2011), .ZN(W2793));
  NOR2X1 G716 (.A1(W1084), .A2(W506), .ZN(W2795));
  NOR2X1 G717 (.A1(W1858), .A2(W1203), .ZN(O195));
  NOR2X1 G718 (.A1(I888), .A2(W1799), .ZN(W2290));
  NOR2X1 G719 (.A1(I643), .A2(W1496), .ZN(W2291));
  NOR2X1 G720 (.A1(W107), .A2(W187), .ZN(O188));
  NOR2X1 G721 (.A1(W1052), .A2(I424), .ZN(W2293));
  NOR2X1 G722 (.A1(I361), .A2(I444), .ZN(W2296));
  NOR2X1 G723 (.A1(W541), .A2(W826), .ZN(O189));
  NOR2X1 G724 (.A1(W2125), .A2(W1486), .ZN(O190));
  NOR2X1 G725 (.A1(W776), .A2(W84), .ZN(W2308));
  NOR2X1 G726 (.A1(W868), .A2(W2044), .ZN(W2310));
  NOR2X1 G727 (.A1(W2177), .A2(W2147), .ZN(W2314));
  NOR2X1 G728 (.A1(W1459), .A2(W2279), .ZN(W2324));
  NOR2X1 G729 (.A1(I554), .A2(I494), .ZN(W2325));
  NOR2X1 G730 (.A1(I998), .A2(I26), .ZN(W2289));
  NOR2X1 G731 (.A1(W972), .A2(I467), .ZN(W2337));
  NOR2X1 G732 (.A1(W2041), .A2(W122), .ZN(W2338));
  NOR2X1 G733 (.A1(W313), .A2(W270), .ZN(O196));
  NOR2X1 G734 (.A1(W798), .A2(W1004), .ZN(W2347));
  NOR2X1 G735 (.A1(I574), .A2(I626), .ZN(W2350));
  NOR2X1 G736 (.A1(W1989), .A2(W1012), .ZN(W2351));
  NOR2X1 G737 (.A1(I925), .A2(I462), .ZN(W2354));
  NOR2X1 G738 (.A1(I458), .A2(I495), .ZN(W2357));
  NOR2X1 G739 (.A1(W1741), .A2(I871), .ZN(W2358));
  NOR2X1 G740 (.A1(W1141), .A2(I530), .ZN(W2371));
  NOR2X1 G741 (.A1(I969), .A2(W175), .ZN(W2374));
  NOR2X1 G742 (.A1(W1085), .A2(I503), .ZN(W2378));
  NOR2X1 G743 (.A1(W51), .A2(W804), .ZN(W2259));
  NOR2X1 G744 (.A1(I864), .A2(W434), .ZN(W2216));
  NOR2X1 G745 (.A1(I235), .A2(W1562), .ZN(W2222));
  NOR2X1 G746 (.A1(I157), .A2(I96), .ZN(W2223));
  NOR2X1 G747 (.A1(W984), .A2(W113), .ZN(W2225));
  NOR2X1 G748 (.A1(W1392), .A2(W1933), .ZN(W2233));
  NOR2X1 G749 (.A1(W2171), .A2(I540), .ZN(W2234));
  NOR2X1 G750 (.A1(W31), .A2(W1025), .ZN(W2239));
  NOR2X1 G751 (.A1(I584), .A2(W74), .ZN(W2241));
  NOR2X1 G752 (.A1(W389), .A2(I100), .ZN(O179));
  NOR2X1 G753 (.A1(W726), .A2(I153), .ZN(W2243));
  NOR2X1 G754 (.A1(W2081), .A2(I970), .ZN(O180));
  NOR2X1 G755 (.A1(W257), .A2(W1489), .ZN(O183));
  NOR2X1 G756 (.A1(W773), .A2(I269), .ZN(W2385));
  NOR2X1 G757 (.A1(I542), .A2(W1666), .ZN(W2260));
  NOR2X1 G758 (.A1(W2026), .A2(W1387), .ZN(W2265));
  NOR2X1 G759 (.A1(I905), .A2(W195), .ZN(W2266));
  NOR2X1 G760 (.A1(W1824), .A2(W1773), .ZN(W2268));
  NOR2X1 G761 (.A1(I380), .A2(I150), .ZN(W2270));
  NOR2X1 G762 (.A1(I184), .A2(W1486), .ZN(W2273));
  NOR2X1 G763 (.A1(W582), .A2(W2087), .ZN(W2275));
  NOR2X1 G764 (.A1(W797), .A2(I792), .ZN(W2276));
  NOR2X1 G765 (.A1(W312), .A2(W973), .ZN(W2278));
  NOR2X1 G766 (.A1(W1513), .A2(W2046), .ZN(W2279));
  NOR2X1 G767 (.A1(W2067), .A2(W1881), .ZN(W2281));
  NOR2X1 G768 (.A1(I939), .A2(W1786), .ZN(W2498));
  NOR2X1 G769 (.A1(W1019), .A2(W2104), .ZN(W2463));
  NOR2X1 G770 (.A1(I544), .A2(W312), .ZN(W2467));
  NOR2X1 G771 (.A1(W2350), .A2(W173), .ZN(W2468));
  NOR2X1 G772 (.A1(W1421), .A2(W1865), .ZN(W2470));
  NOR2X1 G773 (.A1(W1171), .A2(W993), .ZN(W2474));
  NOR2X1 G774 (.A1(W1610), .A2(W2239), .ZN(W2479));
  NOR2X1 G775 (.A1(W1683), .A2(W283), .ZN(W2483));
  NOR2X1 G776 (.A1(W692), .A2(W2275), .ZN(W2486));
  NOR2X1 G777 (.A1(W2102), .A2(I724), .ZN(W2490));
  NOR2X1 G778 (.A1(W1898), .A2(W1734), .ZN(O218));
  NOR2X1 G779 (.A1(W1006), .A2(W496), .ZN(W2494));
  NOR2X1 G780 (.A1(I701), .A2(I546), .ZN(W2496));
  NOR2X1 G781 (.A1(I257), .A2(W1459), .ZN(W2455));
  NOR2X1 G782 (.A1(W2273), .A2(W1255), .ZN(O220));
  NOR2X1 G783 (.A1(I718), .A2(W430), .ZN(O221));
  NOR2X1 G784 (.A1(W923), .A2(I0), .ZN(W2506));
  NOR2X1 G785 (.A1(W1452), .A2(W2285), .ZN(W2508));
  NOR2X1 G786 (.A1(W2382), .A2(W1453), .ZN(W2512));
  NOR2X1 G787 (.A1(I0), .A2(I262), .ZN(W2513));
  NOR2X1 G788 (.A1(W2472), .A2(W2161), .ZN(O225));
  NOR2X1 G789 (.A1(W746), .A2(W2172), .ZN(W2519));
  NOR2X1 G790 (.A1(I912), .A2(W2206), .ZN(W2520));
  NOR2X1 G791 (.A1(W123), .A2(I121), .ZN(W2521));
  NOR2X1 G792 (.A1(W2120), .A2(I592), .ZN(O227));
  NOR2X1 G793 (.A1(W173), .A2(W335), .ZN(W2534));
  NOR2X1 G794 (.A1(W1191), .A2(I79), .ZN(W2424));
  NOR2X1 G795 (.A1(W1631), .A2(I272), .ZN(W2388));
  NOR2X1 G796 (.A1(W2251), .A2(I731), .ZN(W2393));
  NOR2X1 G797 (.A1(W2140), .A2(I410), .ZN(W2394));
  NOR2X1 G798 (.A1(W1160), .A2(W238), .ZN(W2395));
  NOR2X1 G799 (.A1(W987), .A2(W1429), .ZN(W2396));
  NOR2X1 G800 (.A1(W1071), .A2(W1250), .ZN(W2399));
  NOR2X1 G801 (.A1(I620), .A2(W305), .ZN(W2400));
  NOR2X1 G802 (.A1(I153), .A2(I904), .ZN(W2402));
  NOR2X1 G803 (.A1(W1097), .A2(I830), .ZN(W2403));
  NOR2X1 G804 (.A1(W1855), .A2(I976), .ZN(W2405));
  NOR2X1 G805 (.A1(W1792), .A2(I993), .ZN(W2408));
  NOR2X1 G806 (.A1(W1369), .A2(W898), .ZN(W2415));
  NOR2X1 G807 (.A1(W3680), .A2(W4082), .ZN(O731));
  NOR2X1 G808 (.A1(W2195), .A2(W1616), .ZN(W2425));
  NOR2X1 G809 (.A1(W34), .A2(W544), .ZN(W2430));
  NOR2X1 G810 (.A1(I772), .A2(W521), .ZN(W2439));
  NOR2X1 G811 (.A1(I639), .A2(W400), .ZN(O214));
  NOR2X1 G812 (.A1(W465), .A2(W1104), .ZN(W2441));
  NOR2X1 G813 (.A1(W132), .A2(I916), .ZN(W2442));
  NOR2X1 G814 (.A1(W1419), .A2(I538), .ZN(O215));
  NOR2X1 G815 (.A1(W817), .A2(W1952), .ZN(W2446));
  NOR2X1 G816 (.A1(I148), .A2(W104), .ZN(W2447));
  NOR2X1 G817 (.A1(W1878), .A2(W60), .ZN(W2448));
  NOR2X1 G818 (.A1(W197), .A2(W109), .ZN(W2452));
  NOR2X1 G819 (.A1(I826), .A2(W1813), .ZN(O1731));
  NOR2X1 G820 (.A1(W734), .A2(W39), .ZN(O1712));
  NOR2X1 G821 (.A1(W3909), .A2(W3594), .ZN(O1716));
  NOR2X1 G822 (.A1(W244), .A2(W1781), .ZN(O1718));
  NOR2X1 G823 (.A1(W537), .A2(W4916), .ZN(W5710));
  NOR2X1 G824 (.A1(W4322), .A2(W259), .ZN(O1719));
  NOR2X1 G825 (.A1(W834), .A2(W4715), .ZN(O1720));
  NOR2X1 G826 (.A1(W2597), .A2(W1810), .ZN(O1722));
  NOR2X1 G827 (.A1(W5698), .A2(W601), .ZN(O1723));
  NOR2X1 G828 (.A1(W3814), .A2(I741), .ZN(O1725));
  NOR2X1 G829 (.A1(W5111), .A2(W5653), .ZN(O1726));
  NOR2X1 G830 (.A1(W24), .A2(W4168), .ZN(O1727));
  NOR2X1 G831 (.A1(W2484), .A2(W2910), .ZN(O1730));
  NOR2X1 G832 (.A1(W3366), .A2(W1210), .ZN(O1708));
  NOR2X1 G833 (.A1(W265), .A2(W1549), .ZN(O1732));
  NOR2X1 G834 (.A1(W3812), .A2(I705), .ZN(O1737));
  NOR2X1 G835 (.A1(W95), .A2(W1742), .ZN(O1738));
  NOR2X1 G836 (.A1(W5436), .A2(W123), .ZN(W5737));
  NOR2X1 G837 (.A1(W28), .A2(W5442), .ZN(O1744));
  NOR2X1 G838 (.A1(W5354), .A2(W891), .ZN(O1747));
  NOR2X1 G839 (.A1(W422), .A2(W1682), .ZN(O1748));
  NOR2X1 G840 (.A1(W2735), .A2(W2992), .ZN(O1750));
  NOR2X1 G841 (.A1(W2512), .A2(W5273), .ZN(O1751));
  NOR2X1 G842 (.A1(W2412), .A2(W532), .ZN(O1754));
  NOR2X1 G843 (.A1(W2201), .A2(W397), .ZN(O1760));
  NOR2X1 G844 (.A1(W1734), .A2(I450), .ZN(O1766));
  NOR2X1 G845 (.A1(W3162), .A2(I224), .ZN(O1682));
  NOR2X1 G846 (.A1(W1661), .A2(W496), .ZN(O1660));
  NOR2X1 G847 (.A1(W3368), .A2(I210), .ZN(O1661));
  NOR2X1 G848 (.A1(W923), .A2(W4130), .ZN(W5637));
  NOR2X1 G849 (.A1(I661), .A2(W4362), .ZN(W5638));
  NOR2X1 G850 (.A1(W2758), .A2(W4852), .ZN(O1662));
  NOR2X1 G851 (.A1(I862), .A2(W1232), .ZN(O1668));
  NOR2X1 G852 (.A1(W2361), .A2(W829), .ZN(O1672));
  NOR2X1 G853 (.A1(W4298), .A2(W1205), .ZN(O1677));
  NOR2X1 G854 (.A1(W3422), .A2(W1513), .ZN(O1678));
  NOR2X1 G855 (.A1(I697), .A2(W745), .ZN(W5658));
  NOR2X1 G856 (.A1(W2539), .A2(W5288), .ZN(W5659));
  NOR2X1 G857 (.A1(W1820), .A2(W4147), .ZN(O1681));
  NOR2X1 G858 (.A1(W4501), .A2(W3738), .ZN(W5763));
  NOR2X1 G859 (.A1(W3250), .A2(W5056), .ZN(O1688));
  NOR2X1 G860 (.A1(W1989), .A2(W700), .ZN(W5674));
  NOR2X1 G861 (.A1(W4047), .A2(W4304), .ZN(O1690));
  NOR2X1 G862 (.A1(I405), .A2(W4755), .ZN(O1691));
  NOR2X1 G863 (.A1(W1018), .A2(W1664), .ZN(W5679));
  NOR2X1 G864 (.A1(W5665), .A2(W1788), .ZN(W5680));
  NOR2X1 G865 (.A1(W125), .A2(W4294), .ZN(O1694));
  NOR2X1 G866 (.A1(W3605), .A2(W1718), .ZN(O1696));
  NOR2X1 G867 (.A1(W5547), .A2(W3640), .ZN(O1697));
  NOR2X1 G868 (.A1(W694), .A2(I91), .ZN(O1701));
  NOR2X1 G869 (.A1(W1598), .A2(W1389), .ZN(O1703));
  NOR2X1 G870 (.A1(I655), .A2(W194), .ZN(O1704));
  NOR2X1 G871 (.A1(W1004), .A2(W3844), .ZN(O1872));
  NOR2X1 G872 (.A1(W68), .A2(W1745), .ZN(W5852));
  NOR2X1 G873 (.A1(W2720), .A2(I357), .ZN(O1845));
  NOR2X1 G874 (.A1(W1970), .A2(W4590), .ZN(O1848));
  NOR2X1 G875 (.A1(W4313), .A2(W234), .ZN(O1849));
  NOR2X1 G876 (.A1(I288), .A2(W2490), .ZN(O1851));
  NOR2X1 G877 (.A1(W4868), .A2(W2489), .ZN(O1853));
  NOR2X1 G878 (.A1(W1919), .A2(W1048), .ZN(O1855));
  NOR2X1 G879 (.A1(W1899), .A2(W5009), .ZN(O1858));
  NOR2X1 G880 (.A1(W3607), .A2(W1145), .ZN(O1861));
  NOR2X1 G881 (.A1(W1713), .A2(W2751), .ZN(O1866));
  NOR2X1 G882 (.A1(W376), .A2(W1538), .ZN(O1869));
  NOR2X1 G883 (.A1(W1962), .A2(W525), .ZN(O1871));
  NOR2X1 G884 (.A1(I288), .A2(W409), .ZN(W5848));
  NOR2X1 G885 (.A1(W1571), .A2(W1408), .ZN(O1873));
  NOR2X1 G886 (.A1(W958), .A2(W699), .ZN(O1877));
  NOR2X1 G887 (.A1(W5453), .A2(W2927), .ZN(O1879));
  NOR2X1 G888 (.A1(W1198), .A2(W2747), .ZN(O1880));
  NOR2X1 G889 (.A1(W5519), .A2(W3346), .ZN(O1881));
  NOR2X1 G890 (.A1(W3222), .A2(W2160), .ZN(O1884));
  NOR2X1 G891 (.A1(W3852), .A2(I494), .ZN(O1886));
  NOR2X1 G892 (.A1(W4564), .A2(I192), .ZN(O1890));
  NOR2X1 G893 (.A1(W5127), .A2(W2789), .ZN(O1893));
  NOR2X1 G894 (.A1(W4997), .A2(W4124), .ZN(O1898));
  NOR2X1 G895 (.A1(W5118), .A2(W4178), .ZN(O1905));
  NOR2X1 G896 (.A1(W3913), .A2(W693), .ZN(O1907));
  NOR2X1 G897 (.A1(W3406), .A2(W3652), .ZN(W5807));
  NOR2X1 G898 (.A1(W565), .A2(W2640), .ZN(O1771));
  NOR2X1 G899 (.A1(W2485), .A2(W1266), .ZN(O1775));
  NOR2X1 G900 (.A1(W3518), .A2(W3463), .ZN(O1776));
  NOR2X1 G901 (.A1(W3328), .A2(W3536), .ZN(O1777));
  NOR2X1 G902 (.A1(W4638), .A2(W3670), .ZN(O1788));
  NOR2X1 G903 (.A1(W1493), .A2(W3610), .ZN(W5788));
  NOR2X1 G904 (.A1(W109), .A2(W5074), .ZN(O1789));
  NOR2X1 G905 (.A1(W480), .A2(I541), .ZN(O1790));
  NOR2X1 G906 (.A1(W5558), .A2(W2081), .ZN(O1791));
  NOR2X1 G907 (.A1(W1167), .A2(W1324), .ZN(O1794));
  NOR2X1 G908 (.A1(W3542), .A2(W2447), .ZN(O1797));
  NOR2X1 G909 (.A1(W4463), .A2(W2370), .ZN(O1803));
  NOR2X1 G910 (.A1(W1941), .A2(W5622), .ZN(O1657));
  NOR2X1 G911 (.A1(W4519), .A2(W4264), .ZN(O1809));
  NOR2X1 G912 (.A1(W5031), .A2(W797), .ZN(O1813));
  NOR2X1 G913 (.A1(W1227), .A2(W4828), .ZN(O1814));
  NOR2X1 G914 (.A1(W4032), .A2(W903), .ZN(O1817));
  NOR2X1 G915 (.A1(W2322), .A2(W102), .ZN(O1818));
  NOR2X1 G916 (.A1(W3059), .A2(I339), .ZN(O1819));
  NOR2X1 G917 (.A1(W4236), .A2(W5062), .ZN(W5824));
  NOR2X1 G918 (.A1(W5090), .A2(W3957), .ZN(O1820));
  NOR2X1 G919 (.A1(W2060), .A2(W4484), .ZN(O1823));
  NOR2X1 G920 (.A1(W4881), .A2(I750), .ZN(O1828));
  NOR2X1 G921 (.A1(W1601), .A2(W1880), .ZN(W5836));
  NOR2X1 G922 (.A1(W5037), .A2(W2690), .ZN(W5454));
  NOR2X1 G923 (.A1(W3560), .A2(I376), .ZN(O1503));
  NOR2X1 G924 (.A1(W2198), .A2(W2225), .ZN(O1511));
  NOR2X1 G925 (.A1(W4973), .A2(W4754), .ZN(W5436));
  NOR2X1 G926 (.A1(I210), .A2(W2727), .ZN(W5437));
  NOR2X1 G927 (.A1(W4869), .A2(W327), .ZN(O1514));
  NOR2X1 G928 (.A1(W5135), .A2(W4514), .ZN(O1515));
  NOR2X1 G929 (.A1(W1577), .A2(W3276), .ZN(O1516));
  NOR2X1 G930 (.A1(W3225), .A2(W1649), .ZN(W5442));
  NOR2X1 G931 (.A1(W4547), .A2(W2383), .ZN(O1521));
  NOR2X1 G932 (.A1(W3969), .A2(W1320), .ZN(O1522));
  NOR2X1 G933 (.A1(W1261), .A2(W1802), .ZN(O1524));
  NOR2X1 G934 (.A1(W2483), .A2(I986), .ZN(W5452));
  NOR2X1 G935 (.A1(W1665), .A2(W796), .ZN(O1500));
  NOR2X1 G936 (.A1(W3736), .A2(W2241), .ZN(O1526));
  NOR2X1 G937 (.A1(W193), .A2(W4023), .ZN(O1527));
  NOR2X1 G938 (.A1(I714), .A2(W2950), .ZN(O1528));
  NOR2X1 G939 (.A1(W1782), .A2(W780), .ZN(O1529));
  NOR2X1 G940 (.A1(W2162), .A2(W2318), .ZN(O1530));
  NOR2X1 G941 (.A1(W3683), .A2(I533), .ZN(W5468));
  NOR2X1 G942 (.A1(W1119), .A2(W479), .ZN(W5470));
  NOR2X1 G943 (.A1(W4959), .A2(W3251), .ZN(O1538));
  NOR2X1 G944 (.A1(W5307), .A2(W3563), .ZN(O1540));
  NOR2X1 G945 (.A1(I85), .A2(W3796), .ZN(O1541));
  NOR2X1 G946 (.A1(W669), .A2(W2055), .ZN(W5483));
  NOR2X1 G947 (.A1(W4906), .A2(W3834), .ZN(O1547));
  NOR2X1 G948 (.A1(W1692), .A2(W4939), .ZN(O1465));
  NOR2X1 G949 (.A1(W1093), .A2(W4537), .ZN(W5348));
  NOR2X1 G950 (.A1(W2824), .A2(W2370), .ZN(O1445));
  NOR2X1 G951 (.A1(W2814), .A2(W4275), .ZN(W5351));
  NOR2X1 G952 (.A1(W284), .A2(W1118), .ZN(O1448));
  NOR2X1 G953 (.A1(W4851), .A2(W4964), .ZN(W5354));
  NOR2X1 G954 (.A1(W5300), .A2(W4290), .ZN(O1451));
  NOR2X1 G955 (.A1(W3232), .A2(W4170), .ZN(O1453));
  NOR2X1 G956 (.A1(W4080), .A2(W733), .ZN(W5363));
  NOR2X1 G957 (.A1(W2144), .A2(W197), .ZN(O1458));
  NOR2X1 G958 (.A1(W1714), .A2(W3319), .ZN(O1461));
  NOR2X1 G959 (.A1(W4382), .A2(W4364), .ZN(W5371));
  NOR2X1 G960 (.A1(W3023), .A2(W1993), .ZN(O1464));
  NOR2X1 G961 (.A1(W5175), .A2(W1651), .ZN(O1552));
  NOR2X1 G962 (.A1(W967), .A2(I376), .ZN(O1469));
  NOR2X1 G963 (.A1(W4209), .A2(W2142), .ZN(O1470));
  NOR2X1 G964 (.A1(W1408), .A2(W1607), .ZN(O1476));
  NOR2X1 G965 (.A1(W1376), .A2(W1730), .ZN(O1477));
  NOR2X1 G966 (.A1(W983), .A2(W4608), .ZN(O1481));
  NOR2X1 G967 (.A1(W4808), .A2(W4686), .ZN(W5400));
  NOR2X1 G968 (.A1(W4046), .A2(W3903), .ZN(O1486));
  NOR2X1 G969 (.A1(W1302), .A2(W4438), .ZN(W5408));
  NOR2X1 G970 (.A1(W2538), .A2(W2565), .ZN(W5409));
  NOR2X1 G971 (.A1(W1720), .A2(W3398), .ZN(O1492));
  NOR2X1 G972 (.A1(W504), .A2(W1117), .ZN(O1494));
  NOR2X1 G973 (.A1(W22), .A2(I944), .ZN(O1625));
  NOR2X1 G974 (.A1(W4810), .A2(I227), .ZN(W5564));
  NOR2X1 G975 (.A1(W97), .A2(W3776), .ZN(W5567));
  NOR2X1 G976 (.A1(W4598), .A2(W556), .ZN(O1609));
  NOR2X1 G977 (.A1(W1917), .A2(W3419), .ZN(O1610));
  NOR2X1 G978 (.A1(W2255), .A2(I743), .ZN(O1611));
  NOR2X1 G979 (.A1(I360), .A2(W5414), .ZN(O1613));
  NOR2X1 G980 (.A1(W143), .A2(W1492), .ZN(O1618));
  NOR2X1 G981 (.A1(W4928), .A2(W1736), .ZN(O1620));
  NOR2X1 G982 (.A1(W3395), .A2(W3185), .ZN(O1622));
  NOR2X1 G983 (.A1(W1497), .A2(W3947), .ZN(O1623));
  NOR2X1 G984 (.A1(W4402), .A2(W5452), .ZN(W5588));
  NOR2X1 G985 (.A1(W3839), .A2(W645), .ZN(O1624));
  NOR2X1 G986 (.A1(I19), .A2(W2706), .ZN(O1606));
  NOR2X1 G987 (.A1(W4889), .A2(I629), .ZN(O1627));
  NOR2X1 G988 (.A1(W460), .A2(W3474), .ZN(O1629));
  NOR2X1 G989 (.A1(W2970), .A2(W1198), .ZN(O1630));
  NOR2X1 G990 (.A1(I614), .A2(W3911), .ZN(O1634));
  NOR2X1 G991 (.A1(W3423), .A2(W4188), .ZN(O1639));
  NOR2X1 G992 (.A1(W5191), .A2(W2187), .ZN(O1641));
  NOR2X1 G993 (.A1(W3963), .A2(W4515), .ZN(O1646));
  NOR2X1 G994 (.A1(W5510), .A2(W808), .ZN(W5616));
  NOR2X1 G995 (.A1(W4567), .A2(W1029), .ZN(O1647));
  NOR2X1 G996 (.A1(W3547), .A2(W5182), .ZN(O1650));
  NOR2X1 G997 (.A1(W2454), .A2(W2894), .ZN(O1651));
  NOR2X1 G998 (.A1(W3748), .A2(W4600), .ZN(O1655));
  NOR2X1 G999 (.A1(W3594), .A2(W620), .ZN(O1572));
  NOR2X1 G1000 (.A1(W4118), .A2(W3556), .ZN(W5494));
  NOR2X1 G1001 (.A1(W970), .A2(W3945), .ZN(O1555));
  NOR2X1 G1002 (.A1(W3190), .A2(W3194), .ZN(O1557));
  NOR2X1 G1003 (.A1(W1638), .A2(W4006), .ZN(O1558));
  NOR2X1 G1004 (.A1(W2391), .A2(W1577), .ZN(O1563));
  NOR2X1 G1005 (.A1(W4204), .A2(W5371), .ZN(O1564));
  NOR2X1 G1006 (.A1(W5176), .A2(W1785), .ZN(O1565));
  NOR2X1 G1007 (.A1(W5448), .A2(W692), .ZN(W5511));
  NOR2X1 G1008 (.A1(W3778), .A2(I261), .ZN(O1568));
  NOR2X1 G1009 (.A1(W3105), .A2(W2361), .ZN(O1569));
  NOR2X1 G1010 (.A1(W789), .A2(I42), .ZN(O1570));
  NOR2X1 G1011 (.A1(W404), .A2(W4949), .ZN(O1571));
  NOR2X1 G1012 (.A1(I530), .A2(W4572), .ZN(O1912));
  NOR2X1 G1013 (.A1(W3877), .A2(W747), .ZN(O1573));
  NOR2X1 G1014 (.A1(W3980), .A2(W4123), .ZN(O1574));
  NOR2X1 G1015 (.A1(I423), .A2(W998), .ZN(W5529));
  NOR2X1 G1016 (.A1(W5494), .A2(W3891), .ZN(O1580));
  NOR2X1 G1017 (.A1(W2200), .A2(W5515), .ZN(O1584));
  NOR2X1 G1018 (.A1(I882), .A2(W3271), .ZN(O1586));
  NOR2X1 G1019 (.A1(W4588), .A2(W3618), .ZN(W5547));
  NOR2X1 G1020 (.A1(W948), .A2(W4378), .ZN(O1597));
  NOR2X1 G1021 (.A1(W5224), .A2(W4978), .ZN(O1599));
  NOR2X1 G1022 (.A1(W3937), .A2(W4918), .ZN(O1601));
  NOR2X1 G1023 (.A1(W3748), .A2(W419), .ZN(O1605));
  NOR2X1 G1024 (.A1(W3985), .A2(W4149), .ZN(W6329));
  NOR2X1 G1025 (.A1(W2487), .A2(I390), .ZN(O2247));
  NOR2X1 G1026 (.A1(W3495), .A2(I779), .ZN(O2250));
  NOR2X1 G1027 (.A1(W4969), .A2(W3163), .ZN(O2253));
  NOR2X1 G1028 (.A1(W5468), .A2(W5067), .ZN(O2254));
  NOR2X1 G1029 (.A1(I79), .A2(W371), .ZN(O2257));
  NOR2X1 G1030 (.A1(W3238), .A2(W3102), .ZN(O2260));
  NOR2X1 G1031 (.A1(W750), .A2(W2945), .ZN(O2261));
  NOR2X1 G1032 (.A1(W6186), .A2(W4041), .ZN(O2263));
  NOR2X1 G1033 (.A1(W4296), .A2(W457), .ZN(O2264));
  NOR2X1 G1034 (.A1(I516), .A2(W1044), .ZN(O2265));
  NOR2X1 G1035 (.A1(W5470), .A2(W2311), .ZN(O2266));
  NOR2X1 G1036 (.A1(W4732), .A2(W1735), .ZN(O2269));
  NOR2X1 G1037 (.A1(W5286), .A2(I72), .ZN(O2244));
  NOR2X1 G1038 (.A1(W3003), .A2(I223), .ZN(O2279));
  NOR2X1 G1039 (.A1(W6022), .A2(I791), .ZN(O2280));
  NOR2X1 G1040 (.A1(W2772), .A2(W4697), .ZN(W6334));
  NOR2X1 G1041 (.A1(W3026), .A2(W2704), .ZN(O2286));
  NOR2X1 G1042 (.A1(W676), .A2(W4393), .ZN(O2289));
  NOR2X1 G1043 (.A1(W6334), .A2(I906), .ZN(O2296));
  NOR2X1 G1044 (.A1(W5638), .A2(W5424), .ZN(O2303));
  NOR2X1 G1045 (.A1(I937), .A2(I631), .ZN(O2304));
  NOR2X1 G1046 (.A1(W412), .A2(W5404), .ZN(O2307));
  NOR2X1 G1047 (.A1(W4840), .A2(W4697), .ZN(O2309));
  NOR2X1 G1048 (.A1(W1935), .A2(I257), .ZN(O2311));
  NOR2X1 G1049 (.A1(W4437), .A2(W5806), .ZN(O2312));
  NOR2X1 G1050 (.A1(W6101), .A2(I300), .ZN(W6267));
  NOR2X1 G1051 (.A1(W5841), .A2(W5191), .ZN(O2195));
  NOR2X1 G1052 (.A1(W3421), .A2(W5931), .ZN(O2197));
  NOR2X1 G1053 (.A1(W1367), .A2(W319), .ZN(O2198));
  NOR2X1 G1054 (.A1(W4572), .A2(W4343), .ZN(O2199));
  NOR2X1 G1055 (.A1(W5964), .A2(W2747), .ZN(O2202));
  NOR2X1 G1056 (.A1(W3425), .A2(W1998), .ZN(O2203));
  NOR2X1 G1057 (.A1(W4935), .A2(W540), .ZN(O2205));
  NOR2X1 G1058 (.A1(W6009), .A2(W4953), .ZN(O2209));
  NOR2X1 G1059 (.A1(W2841), .A2(W2232), .ZN(O2210));
  NOR2X1 G1060 (.A1(W54), .A2(I507), .ZN(O2211));
  NOR2X1 G1061 (.A1(W213), .A2(I870), .ZN(O2212));
  NOR2X1 G1062 (.A1(W873), .A2(W4073), .ZN(W6262));
  NOR2X1 G1063 (.A1(W88), .A2(I650), .ZN(O2313));
  NOR2X1 G1064 (.A1(W3786), .A2(I424), .ZN(O2220));
  NOR2X1 G1065 (.A1(W5206), .A2(W3345), .ZN(O2224));
  NOR2X1 G1066 (.A1(W1507), .A2(W1137), .ZN(O2225));
  NOR2X1 G1067 (.A1(W3269), .A2(W5616), .ZN(O2227));
  NOR2X1 G1068 (.A1(W4150), .A2(I227), .ZN(O2228));
  NOR2X1 G1069 (.A1(W4276), .A2(W3704), .ZN(O2229));
  NOR2X1 G1070 (.A1(W3870), .A2(I802), .ZN(O2231));
  NOR2X1 G1071 (.A1(W4272), .A2(W4482), .ZN(O2237));
  NOR2X1 G1072 (.A1(W5657), .A2(W5619), .ZN(O2238));
  NOR2X1 G1073 (.A1(W777), .A2(W1474), .ZN(O2239));
  NOR2X1 G1074 (.A1(W1189), .A2(W111), .ZN(O2240));
  NOR2X1 G1075 (.A1(W2792), .A2(W3071), .ZN(O2243));
  NOR2X1 G1076 (.A1(W1756), .A2(W1515), .ZN(O2416));
  NOR2X1 G1077 (.A1(W5587), .A2(W544), .ZN(O2377));
  NOR2X1 G1078 (.A1(W2937), .A2(W2960), .ZN(O2378));
  NOR2X1 G1079 (.A1(W6015), .A2(W5848), .ZN(O2381));
  NOR2X1 G1080 (.A1(W2443), .A2(W4064), .ZN(O2385));
  NOR2X1 G1081 (.A1(W854), .A2(W4608), .ZN(O2391));
  NOR2X1 G1082 (.A1(W3205), .A2(I613), .ZN(O2397));
  NOR2X1 G1083 (.A1(W487), .A2(W708), .ZN(O2399));
  NOR2X1 G1084 (.A1(W879), .A2(W3840), .ZN(O2400));
  NOR2X1 G1085 (.A1(W2506), .A2(I320), .ZN(O2405));
  NOR2X1 G1086 (.A1(W5858), .A2(W5843), .ZN(O2407));
  NOR2X1 G1087 (.A1(I890), .A2(W5543), .ZN(O2408));
  NOR2X1 G1088 (.A1(W5001), .A2(W1750), .ZN(O2413));
  NOR2X1 G1089 (.A1(W4816), .A2(I929), .ZN(O2375));
  NOR2X1 G1090 (.A1(W996), .A2(W3230), .ZN(O2418));
  NOR2X1 G1091 (.A1(W1357), .A2(W3122), .ZN(O2421));
  NOR2X1 G1092 (.A1(W958), .A2(W2807), .ZN(O2425));
  NOR2X1 G1093 (.A1(I913), .A2(W25), .ZN(O2426));
  NOR2X1 G1094 (.A1(W334), .A2(W5002), .ZN(O2428));
  NOR2X1 G1095 (.A1(W156), .A2(W6237), .ZN(O2432));
  NOR2X1 G1096 (.A1(W2573), .A2(W2862), .ZN(O2437));
  NOR2X1 G1097 (.A1(W2835), .A2(W3676), .ZN(O2440));
  NOR2X1 G1098 (.A1(W571), .A2(W399), .ZN(O2441));
  NOR2X1 G1099 (.A1(W2037), .A2(W5149), .ZN(O2444));
  NOR2X1 G1100 (.A1(W1469), .A2(W3642), .ZN(O2445));
  NOR2X1 G1101 (.A1(W4655), .A2(O2337), .ZN(O2448));
  NOR2X1 G1102 (.A1(W932), .A2(W3519), .ZN(O2339));
  NOR2X1 G1103 (.A1(W1128), .A2(W5788), .ZN(O2314));
  NOR2X1 G1104 (.A1(W5841), .A2(W2598), .ZN(O2315));
  NOR2X1 G1105 (.A1(W3298), .A2(W2175), .ZN(O2317));
  NOR2X1 G1106 (.A1(W1619), .A2(W751), .ZN(O2318));
  NOR2X1 G1107 (.A1(I862), .A2(I218), .ZN(O2319));
  NOR2X1 G1108 (.A1(W3246), .A2(W941), .ZN(O2320));
  NOR2X1 G1109 (.A1(I810), .A2(W1056), .ZN(O2325));
  NOR2X1 G1110 (.A1(W3298), .A2(W1597), .ZN(O2327));
  NOR2X1 G1111 (.A1(W1447), .A2(I793), .ZN(O2329));
  NOR2X1 G1112 (.A1(W3830), .A2(W2343), .ZN(O2333));
  NOR2X1 G1113 (.A1(W1168), .A2(W2934), .ZN(O2335));
  NOR2X1 G1114 (.A1(W4262), .A2(I610), .ZN(O2337));
  NOR2X1 G1115 (.A1(W1118), .A2(W4135), .ZN(O2194));
  NOR2X1 G1116 (.A1(W4447), .A2(W2179), .ZN(O2340));
  NOR2X1 G1117 (.A1(W3015), .A2(I819), .ZN(O2343));
  NOR2X1 G1118 (.A1(W3769), .A2(W383), .ZN(O2344));
  NOR2X1 G1119 (.A1(W3504), .A2(W518), .ZN(O2346));
  NOR2X1 G1120 (.A1(W4468), .A2(I986), .ZN(O2350));
  NOR2X1 G1121 (.A1(W294), .A2(W5002), .ZN(O2352));
  NOR2X1 G1122 (.A1(W4588), .A2(W611), .ZN(O2353));
  NOR2X1 G1123 (.A1(W6082), .A2(W645), .ZN(O2357));
  NOR2X1 G1124 (.A1(W3409), .A2(W6133), .ZN(O2360));
  NOR2X1 G1125 (.A1(W3947), .A2(W2974), .ZN(O2361));
  NOR2X1 G1126 (.A1(W3569), .A2(W1910), .ZN(O2370));
  NOR2X1 G1127 (.A1(W214), .A2(W4640), .ZN(O2011));
  NOR2X1 G1128 (.A1(I660), .A2(I422), .ZN(O1988));
  NOR2X1 G1129 (.A1(W1173), .A2(W4369), .ZN(O1992));
  NOR2X1 G1130 (.A1(I740), .A2(W2677), .ZN(W6022));
  NOR2X1 G1131 (.A1(I434), .A2(W3004), .ZN(O1994));
  NOR2X1 G1132 (.A1(W1083), .A2(W3263), .ZN(O1996));
  NOR2X1 G1133 (.A1(W947), .A2(W1558), .ZN(O1998));
  NOR2X1 G1134 (.A1(W3896), .A2(W3716), .ZN(O2000));
  NOR2X1 G1135 (.A1(W932), .A2(W5239), .ZN(O2001));
  NOR2X1 G1136 (.A1(W4724), .A2(W2078), .ZN(O2003));
  NOR2X1 G1137 (.A1(W842), .A2(I815), .ZN(O2005));
  NOR2X1 G1138 (.A1(I162), .A2(W1364), .ZN(O2008));
  NOR2X1 G1139 (.A1(W1036), .A2(W5588), .ZN(O2010));
  NOR2X1 G1140 (.A1(W5595), .A2(W4431), .ZN(W6015));
  NOR2X1 G1141 (.A1(W1786), .A2(W4811), .ZN(O2012));
  NOR2X1 G1142 (.A1(W4283), .A2(W3818), .ZN(O2014));
  NOR2X1 G1143 (.A1(W304), .A2(W4801), .ZN(W6055));
  NOR2X1 G1144 (.A1(W5144), .A2(W2099), .ZN(O2024));
  NOR2X1 G1145 (.A1(W2169), .A2(W4528), .ZN(O2025));
  NOR2X1 G1146 (.A1(W1408), .A2(W4395), .ZN(O2026));
  NOR2X1 G1147 (.A1(W3497), .A2(W4579), .ZN(O2029));
  NOR2X1 G1148 (.A1(W1708), .A2(I361), .ZN(O2030));
  NOR2X1 G1149 (.A1(W2474), .A2(W4669), .ZN(O2033));
  NOR2X1 G1150 (.A1(W5623), .A2(W1042), .ZN(O2035));
  NOR2X1 G1151 (.A1(W4191), .A2(W3810), .ZN(O2039));
  NOR2X1 G1152 (.A1(W314), .A2(W2474), .ZN(W6075));
  NOR2X1 G1153 (.A1(W121), .A2(W2832), .ZN(O1942));
  NOR2X1 G1154 (.A1(W3522), .A2(I944), .ZN(O1914));
  NOR2X1 G1155 (.A1(W3577), .A2(W2496), .ZN(W5936));
  NOR2X1 G1156 (.A1(W1383), .A2(W4508), .ZN(O1916));
  NOR2X1 G1157 (.A1(I829), .A2(W3827), .ZN(W5938));
  NOR2X1 G1158 (.A1(I817), .A2(W724), .ZN(O1920));
  NOR2X1 G1159 (.A1(W1603), .A2(W4447), .ZN(O1922));
  NOR2X1 G1160 (.A1(I443), .A2(W5357), .ZN(O1928));
  NOR2X1 G1161 (.A1(W4266), .A2(W5855), .ZN(O1936));
  NOR2X1 G1162 (.A1(W2339), .A2(W177), .ZN(O1937));
  NOR2X1 G1163 (.A1(W2792), .A2(W24), .ZN(O1939));
  NOR2X1 G1164 (.A1(W1223), .A2(W1073), .ZN(O1941));
  NOR2X1 G1165 (.A1(W3258), .A2(I595), .ZN(W5964));
  NOR2X1 G1166 (.A1(W1577), .A2(W2346), .ZN(O2045));
  NOR2X1 G1167 (.A1(W607), .A2(W2484), .ZN(O1944));
  NOR2X1 G1168 (.A1(W479), .A2(W3983), .ZN(O1956));
  NOR2X1 G1169 (.A1(W1898), .A2(W5891), .ZN(O1959));
  NOR2X1 G1170 (.A1(W1439), .A2(W204), .ZN(W5985));
  NOR2X1 G1171 (.A1(W3312), .A2(W2185), .ZN(O1961));
  NOR2X1 G1172 (.A1(W443), .A2(W469), .ZN(O1966));
  NOR2X1 G1173 (.A1(W5700), .A2(W2764), .ZN(O1968));
  NOR2X1 G1174 (.A1(W2540), .A2(W4949), .ZN(O1974));
  NOR2X1 G1175 (.A1(W2551), .A2(W1894), .ZN(O1975));
  NOR2X1 G1176 (.A1(W5591), .A2(W894), .ZN(O1979));
  NOR2X1 G1177 (.A1(W5725), .A2(W1171), .ZN(W6009));
  NOR2X1 G1178 (.A1(W5253), .A2(W3125), .ZN(O2157));
  NOR2X1 G1179 (.A1(W4520), .A2(W3099), .ZN(O2126));
  NOR2X1 G1180 (.A1(W3674), .A2(I674), .ZN(O2128));
  NOR2X1 G1181 (.A1(I416), .A2(W1853), .ZN(O2131));
  NOR2X1 G1182 (.A1(W4978), .A2(W3409), .ZN(O2132));
  NOR2X1 G1183 (.A1(W3603), .A2(W2153), .ZN(O2135));
  NOR2X1 G1184 (.A1(W4586), .A2(W978), .ZN(O2137));
  NOR2X1 G1185 (.A1(W292), .A2(I495), .ZN(O2138));
  NOR2X1 G1186 (.A1(W4007), .A2(I722), .ZN(O2145));
  NOR2X1 G1187 (.A1(W1613), .A2(W2508), .ZN(O2147));
  NOR2X1 G1188 (.A1(W2280), .A2(W3565), .ZN(O2148));
  NOR2X1 G1189 (.A1(W4006), .A2(W3484), .ZN(O2150));
  NOR2X1 G1190 (.A1(W3866), .A2(W3556), .ZN(O2152));
  NOR2X1 G1191 (.A1(W4783), .A2(W1991), .ZN(O2117));
  NOR2X1 G1192 (.A1(W3532), .A2(W2028), .ZN(O2159));
  NOR2X1 G1193 (.A1(W353), .A2(W4259), .ZN(O2165));
  NOR2X1 G1194 (.A1(W1), .A2(W5680), .ZN(O2167));
  NOR2X1 G1195 (.A1(I464), .A2(W969), .ZN(O2170));
  NOR2X1 G1196 (.A1(W1163), .A2(I999), .ZN(O2172));
  NOR2X1 G1197 (.A1(I477), .A2(I647), .ZN(O2173));
  NOR2X1 G1198 (.A1(W4632), .A2(W3544), .ZN(O2174));
  NOR2X1 G1199 (.A1(W3614), .A2(I196), .ZN(O2179));
  NOR2X1 G1200 (.A1(W674), .A2(I116), .ZN(O2180));
  NOR2X1 G1201 (.A1(W3734), .A2(W5186), .ZN(O2185));
  NOR2X1 G1202 (.A1(W3511), .A2(W5457), .ZN(W6232));
  NOR2X1 G1203 (.A1(W726), .A2(W6154), .ZN(O2191));
  NOR2X1 G1204 (.A1(W4103), .A2(W237), .ZN(O2080));
  NOR2X1 G1205 (.A1(W4398), .A2(W32), .ZN(W6082));
  NOR2X1 G1206 (.A1(W923), .A2(W2337), .ZN(O2048));
  NOR2X1 G1207 (.A1(W3390), .A2(W1150), .ZN(O2051));
  NOR2X1 G1208 (.A1(W2523), .A2(W4596), .ZN(O2054));
  NOR2X1 G1209 (.A1(W5666), .A2(W257), .ZN(O2061));
  NOR2X1 G1210 (.A1(W4663), .A2(W2364), .ZN(O2062));
  NOR2X1 G1211 (.A1(W3879), .A2(W604), .ZN(O2068));
  NOR2X1 G1212 (.A1(W91), .A2(W5191), .ZN(O2070));
  NOR2X1 G1213 (.A1(W5806), .A2(W1663), .ZN(O2072));
  NOR2X1 G1214 (.A1(W5029), .A2(W2653), .ZN(O2076));
  NOR2X1 G1215 (.A1(W4188), .A2(W4517), .ZN(O2077));
  NOR2X1 G1216 (.A1(W4803), .A2(W1220), .ZN(O2078));
  NOR2X1 G1217 (.A1(W4534), .A2(W3211), .ZN(O1435));
  NOR2X1 G1218 (.A1(W3210), .A2(W3820), .ZN(O2081));
  NOR2X1 G1219 (.A1(W1751), .A2(W5525), .ZN(O2082));
  NOR2X1 G1220 (.A1(W5191), .A2(W1956), .ZN(O2085));
  NOR2X1 G1221 (.A1(I407), .A2(W1393), .ZN(O2086));
  NOR2X1 G1222 (.A1(W4209), .A2(W727), .ZN(O2089));
  NOR2X1 G1223 (.A1(W2710), .A2(W6039), .ZN(W6133));
  NOR2X1 G1224 (.A1(I218), .A2(W2992), .ZN(O2095));
  NOR2X1 G1225 (.A1(W4000), .A2(W5436), .ZN(O2101));
  NOR2X1 G1226 (.A1(W1968), .A2(W157), .ZN(O2102));
  NOR2X1 G1227 (.A1(W1502), .A2(W3883), .ZN(O2112));
  NOR2X1 G1228 (.A1(W2786), .A2(W5527), .ZN(O2115));
  NOR2X1 G1229 (.A1(W1425), .A2(I527), .ZN(W4559));
  NOR2X1 G1230 (.A1(W3674), .A2(W1566), .ZN(O932));
  NOR2X1 G1231 (.A1(W1471), .A2(W3902), .ZN(O933));
  NOR2X1 G1232 (.A1(W822), .A2(I84), .ZN(O934));
  NOR2X1 G1233 (.A1(W307), .A2(W768), .ZN(W4535));
  NOR2X1 G1234 (.A1(W751), .A2(I626), .ZN(O935));
  NOR2X1 G1235 (.A1(W2788), .A2(W4067), .ZN(O936));
  NOR2X1 G1236 (.A1(W3102), .A2(W620), .ZN(W4542));
  NOR2X1 G1237 (.A1(W2736), .A2(W2942), .ZN(O942));
  NOR2X1 G1238 (.A1(I209), .A2(W1583), .ZN(O944));
  NOR2X1 G1239 (.A1(W1605), .A2(W2375), .ZN(O947));
  NOR2X1 G1240 (.A1(W905), .A2(W4526), .ZN(O948));
  NOR2X1 G1241 (.A1(W1335), .A2(W3030), .ZN(W4558));
  NOR2X1 G1242 (.A1(W1977), .A2(W4518), .ZN(O931));
  NOR2X1 G1243 (.A1(W2583), .A2(W1886), .ZN(O950));
  NOR2X1 G1244 (.A1(W3256), .A2(I247), .ZN(W4569));
  NOR2X1 G1245 (.A1(W559), .A2(W1577), .ZN(O959));
  NOR2X1 G1246 (.A1(W4348), .A2(I326), .ZN(W4578));
  NOR2X1 G1247 (.A1(W1953), .A2(W2842), .ZN(O961));
  NOR2X1 G1248 (.A1(W3411), .A2(W765), .ZN(O962));
  NOR2X1 G1249 (.A1(W3806), .A2(W4136), .ZN(W4585));
  NOR2X1 G1250 (.A1(I882), .A2(W285), .ZN(W4588));
  NOR2X1 G1251 (.A1(W2946), .A2(I923), .ZN(W4589));
  NOR2X1 G1252 (.A1(W3343), .A2(W2246), .ZN(W4602));
  NOR2X1 G1253 (.A1(W345), .A2(W3722), .ZN(O970));
  NOR2X1 G1254 (.A1(W867), .A2(I530), .ZN(W4604));
  NOR2X1 G1255 (.A1(W2983), .A2(W1598), .ZN(W4480));
  NOR2X1 G1256 (.A1(W3130), .A2(W1494), .ZN(W4452));
  NOR2X1 G1257 (.A1(W3963), .A2(W2592), .ZN(O889));
  NOR2X1 G1258 (.A1(W3320), .A2(W1278), .ZN(W4454));
  NOR2X1 G1259 (.A1(W405), .A2(W2425), .ZN(O890));
  NOR2X1 G1260 (.A1(W1144), .A2(W2102), .ZN(O892));
  NOR2X1 G1261 (.A1(W3666), .A2(W702), .ZN(O893));
  NOR2X1 G1262 (.A1(W2747), .A2(W581), .ZN(O895));
  NOR2X1 G1263 (.A1(I908), .A2(W1277), .ZN(O899));
  NOR2X1 G1264 (.A1(W348), .A2(W526), .ZN(W4467));
  NOR2X1 G1265 (.A1(I163), .A2(I622), .ZN(O900));
  NOR2X1 G1266 (.A1(W243), .A2(W1565), .ZN(O902));
  NOR2X1 G1267 (.A1(W144), .A2(I649), .ZN(O905));
  NOR2X1 G1268 (.A1(I296), .A2(I38), .ZN(W4607));
  NOR2X1 G1269 (.A1(W2693), .A2(W1219), .ZN(O914));
  NOR2X1 G1270 (.A1(W3534), .A2(W1581), .ZN(W4491));
  NOR2X1 G1271 (.A1(W2908), .A2(W3304), .ZN(W4506));
  NOR2X1 G1272 (.A1(W853), .A2(W50), .ZN(O923));
  NOR2X1 G1273 (.A1(W321), .A2(W2461), .ZN(W4514));
  NOR2X1 G1274 (.A1(W1847), .A2(W2789), .ZN(W4515));
  NOR2X1 G1275 (.A1(W3568), .A2(W841), .ZN(W4517));
  NOR2X1 G1276 (.A1(W1701), .A2(W2282), .ZN(W4520));
  NOR2X1 G1277 (.A1(W2423), .A2(W3127), .ZN(W4521));
  NOR2X1 G1278 (.A1(W700), .A2(W993), .ZN(W4522));
  NOR2X1 G1279 (.A1(W2682), .A2(I730), .ZN(O927));
  NOR2X1 G1280 (.A1(W43), .A2(W580), .ZN(W4527));
  NOR2X1 G1281 (.A1(W1260), .A2(I407), .ZN(O1034));
  NOR2X1 G1282 (.A1(W449), .A2(W990), .ZN(O1004));
  NOR2X1 G1283 (.A1(W576), .A2(W4319), .ZN(W4684));
  NOR2X1 G1284 (.A1(I354), .A2(W1790), .ZN(O1010));
  NOR2X1 G1285 (.A1(W4184), .A2(W2423), .ZN(W4686));
  NOR2X1 G1286 (.A1(W2386), .A2(W4509), .ZN(O1011));
  NOR2X1 G1287 (.A1(W711), .A2(W1999), .ZN(O1013));
  NOR2X1 G1288 (.A1(W2193), .A2(W2996), .ZN(O1015));
  NOR2X1 G1289 (.A1(W3813), .A2(W817), .ZN(W4695));
  NOR2X1 G1290 (.A1(W2255), .A2(W4042), .ZN(O1020));
  NOR2X1 G1291 (.A1(W1273), .A2(W4), .ZN(O1023));
  NOR2X1 G1292 (.A1(W2606), .A2(W3128), .ZN(W4707));
  NOR2X1 G1293 (.A1(W3396), .A2(W1524), .ZN(O1024));
  NOR2X1 G1294 (.A1(W937), .A2(W3911), .ZN(W4675));
  NOR2X1 G1295 (.A1(W516), .A2(W340), .ZN(W4723));
  NOR2X1 G1296 (.A1(W2917), .A2(W4364), .ZN(W4725));
  NOR2X1 G1297 (.A1(W3344), .A2(W3608), .ZN(O1036));
  NOR2X1 G1298 (.A1(W4102), .A2(W3670), .ZN(O1037));
  NOR2X1 G1299 (.A1(W633), .A2(W1919), .ZN(O1038));
  NOR2X1 G1300 (.A1(W1349), .A2(W1924), .ZN(O1043));
  NOR2X1 G1301 (.A1(W4548), .A2(W471), .ZN(W4736));
  NOR2X1 G1302 (.A1(W1558), .A2(W4602), .ZN(O1046));
  NOR2X1 G1303 (.A1(W4014), .A2(W4088), .ZN(O1047));
  NOR2X1 G1304 (.A1(W192), .A2(W1583), .ZN(W4748));
  NOR2X1 G1305 (.A1(W278), .A2(W3422), .ZN(W4749));
  NOR2X1 G1306 (.A1(W4585), .A2(W754), .ZN(O1052));
  NOR2X1 G1307 (.A1(W4292), .A2(W1276), .ZN(O986));
  NOR2X1 G1308 (.A1(W2856), .A2(I116), .ZN(W4608));
  NOR2X1 G1309 (.A1(W4221), .A2(W679), .ZN(O972));
  NOR2X1 G1310 (.A1(W4609), .A2(I463), .ZN(W4613));
  NOR2X1 G1311 (.A1(I548), .A2(W3374), .ZN(W4615));
  NOR2X1 G1312 (.A1(W2668), .A2(W3022), .ZN(O979));
  NOR2X1 G1313 (.A1(W2614), .A2(W1406), .ZN(W4622));
  NOR2X1 G1314 (.A1(W1468), .A2(I451), .ZN(O981));
  NOR2X1 G1315 (.A1(W3721), .A2(W2967), .ZN(O982));
  NOR2X1 G1316 (.A1(W335), .A2(W4506), .ZN(W4627));
  NOR2X1 G1317 (.A1(I764), .A2(W3155), .ZN(W4630));
  NOR2X1 G1318 (.A1(I402), .A2(W883), .ZN(O983));
  NOR2X1 G1319 (.A1(W2934), .A2(W4333), .ZN(O985));
  NOR2X1 G1320 (.A1(W155), .A2(W559), .ZN(O881));
  NOR2X1 G1321 (.A1(W3189), .A2(W4452), .ZN(W4640));
  NOR2X1 G1322 (.A1(W3662), .A2(I615), .ZN(O987));
  NOR2X1 G1323 (.A1(W2497), .A2(W2209), .ZN(O988));
  NOR2X1 G1324 (.A1(W417), .A2(W1804), .ZN(O989));
  NOR2X1 G1325 (.A1(W4053), .A2(W1540), .ZN(W4647));
  NOR2X1 G1326 (.A1(I672), .A2(I214), .ZN(W4653));
  NOR2X1 G1327 (.A1(W1876), .A2(W642), .ZN(O993));
  NOR2X1 G1328 (.A1(W692), .A2(W3014), .ZN(W4657));
  NOR2X1 G1329 (.A1(W1777), .A2(W2511), .ZN(W4659));
  NOR2X1 G1330 (.A1(W3100), .A2(W721), .ZN(W4669));
  NOR2X1 G1331 (.A1(W2579), .A2(I587), .ZN(O1003));
  NOR2X1 G1332 (.A1(I346), .A2(W3206), .ZN(O789));
  NOR2X1 G1333 (.A1(W2422), .A2(W818), .ZN(W4170));
  NOR2X1 G1334 (.A1(W1198), .A2(W883), .ZN(W4174));
  NOR2X1 G1335 (.A1(W3698), .A2(W2131), .ZN(W4176));
  NOR2X1 G1336 (.A1(W573), .A2(W4088), .ZN(W4177));
  NOR2X1 G1337 (.A1(W1169), .A2(W1034), .ZN(O768));
  NOR2X1 G1338 (.A1(W1033), .A2(W1048), .ZN(W4194));
  NOR2X1 G1339 (.A1(W1728), .A2(W995), .ZN(O773));
  NOR2X1 G1340 (.A1(I75), .A2(W2574), .ZN(W4203));
  NOR2X1 G1341 (.A1(W2227), .A2(I623), .ZN(O783));
  NOR2X1 G1342 (.A1(W2467), .A2(W1343), .ZN(O784));
  NOR2X1 G1343 (.A1(W2593), .A2(W3376), .ZN(W4215));
  NOR2X1 G1344 (.A1(W211), .A2(W2150), .ZN(W4216));
  NOR2X1 G1345 (.A1(W1969), .A2(W3523), .ZN(W4168));
  NOR2X1 G1346 (.A1(W3881), .A2(W3764), .ZN(O796));
  NOR2X1 G1347 (.A1(W2118), .A2(W60), .ZN(W4236));
  NOR2X1 G1348 (.A1(W249), .A2(W83), .ZN(O804));
  NOR2X1 G1349 (.A1(I486), .A2(W19), .ZN(W4245));
  NOR2X1 G1350 (.A1(W1311), .A2(W3246), .ZN(O805));
  NOR2X1 G1351 (.A1(W327), .A2(W2742), .ZN(O806));
  NOR2X1 G1352 (.A1(W538), .A2(I519), .ZN(W4250));
  NOR2X1 G1353 (.A1(W282), .A2(W1350), .ZN(O807));
  NOR2X1 G1354 (.A1(I704), .A2(W2971), .ZN(W4253));
  NOR2X1 G1355 (.A1(I502), .A2(W2072), .ZN(O808));
  NOR2X1 G1356 (.A1(W114), .A2(W1377), .ZN(W4262));
  NOR2X1 G1357 (.A1(W2714), .A2(W1165), .ZN(W4264));
  NOR2X1 G1358 (.A1(W694), .A2(W1689), .ZN(W4131));
  NOR2X1 G1359 (.A1(W1388), .A2(W2713), .ZN(W4094));
  NOR2X1 G1360 (.A1(I632), .A2(W3551), .ZN(O733));
  NOR2X1 G1361 (.A1(I728), .A2(I777), .ZN(W4099));
  NOR2X1 G1362 (.A1(W2856), .A2(W4077), .ZN(W4100));
  NOR2X1 G1363 (.A1(W2133), .A2(W3461), .ZN(W4102));
  NOR2X1 G1364 (.A1(I80), .A2(W3887), .ZN(W4103));
  NOR2X1 G1365 (.A1(W2362), .A2(W2403), .ZN(O735));
  NOR2X1 G1366 (.A1(W3111), .A2(W289), .ZN(W4106));
  NOR2X1 G1367 (.A1(W3907), .A2(I962), .ZN(W4120));
  NOR2X1 G1368 (.A1(W2063), .A2(W306), .ZN(O745));
  NOR2X1 G1369 (.A1(W2629), .A2(W623), .ZN(W4128));
  NOR2X1 G1370 (.A1(W2216), .A2(W687), .ZN(O747));
  NOR2X1 G1371 (.A1(I20), .A2(W3691), .ZN(W4267));
  NOR2X1 G1372 (.A1(W4024), .A2(W2316), .ZN(W4132));
  NOR2X1 G1373 (.A1(W3562), .A2(I406), .ZN(O748));
  NOR2X1 G1374 (.A1(I132), .A2(W3509), .ZN(O750));
  NOR2X1 G1375 (.A1(W3017), .A2(W2865), .ZN(O751));
  NOR2X1 G1376 (.A1(W48), .A2(W2008), .ZN(W4142));
  NOR2X1 G1377 (.A1(W1127), .A2(W3001), .ZN(O753));
  NOR2X1 G1378 (.A1(W3708), .A2(I162), .ZN(W4146));
  NOR2X1 G1379 (.A1(W1917), .A2(W1558), .ZN(W4147));
  NOR2X1 G1380 (.A1(W1363), .A2(W1396), .ZN(W4157));
  NOR2X1 G1381 (.A1(W1583), .A2(W2088), .ZN(O761));
  NOR2X1 G1382 (.A1(W645), .A2(W2226), .ZN(O763));
  NOR2X1 G1383 (.A1(W3663), .A2(W3490), .ZN(W4390));
  NOR2X1 G1384 (.A1(W2364), .A2(W1237), .ZN(W4357));
  NOR2X1 G1385 (.A1(W921), .A2(W2793), .ZN(W4359));
  NOR2X1 G1386 (.A1(I925), .A2(W3441), .ZN(W4364));
  NOR2X1 G1387 (.A1(W4100), .A2(W1594), .ZN(O846));
  NOR2X1 G1388 (.A1(W3119), .A2(W1342), .ZN(W4371));
  NOR2X1 G1389 (.A1(W2240), .A2(W3112), .ZN(O849));
  NOR2X1 G1390 (.A1(W774), .A2(I880), .ZN(W4380));
  NOR2X1 G1391 (.A1(W1293), .A2(W3200), .ZN(W4381));
  NOR2X1 G1392 (.A1(W38), .A2(W3774), .ZN(W4382));
  NOR2X1 G1393 (.A1(W851), .A2(I885), .ZN(W4383));
  NOR2X1 G1394 (.A1(W4299), .A2(W1211), .ZN(W4386));
  NOR2X1 G1395 (.A1(W3508), .A2(W17), .ZN(W4389));
  NOR2X1 G1396 (.A1(W2465), .A2(W883), .ZN(O843));
  NOR2X1 G1397 (.A1(I664), .A2(W2871), .ZN(W4392));
  NOR2X1 G1398 (.A1(W1027), .A2(W1450), .ZN(W4398));
  NOR2X1 G1399 (.A1(W3552), .A2(W2112), .ZN(W4405));
  NOR2X1 G1400 (.A1(W139), .A2(W2278), .ZN(W4413));
  NOR2X1 G1401 (.A1(W132), .A2(W1897), .ZN(O866));
  NOR2X1 G1402 (.A1(W2173), .A2(W3624), .ZN(O867));
  NOR2X1 G1403 (.A1(W948), .A2(W885), .ZN(O869));
  NOR2X1 G1404 (.A1(W3115), .A2(I508), .ZN(O871));
  NOR2X1 G1405 (.A1(W1223), .A2(W3763), .ZN(W4423));
  NOR2X1 G1406 (.A1(W972), .A2(W3009), .ZN(O873));
  NOR2X1 G1407 (.A1(W64), .A2(I752), .ZN(O878));
  NOR2X1 G1408 (.A1(W4078), .A2(W3862), .ZN(O879));
  NOR2X1 G1409 (.A1(I864), .A2(W3431), .ZN(O819));
  NOR2X1 G1410 (.A1(W405), .A2(W448), .ZN(W4270));
  NOR2X1 G1411 (.A1(W3186), .A2(W2583), .ZN(W4280));
  NOR2X1 G1412 (.A1(W1219), .A2(W635), .ZN(W4281));
  NOR2X1 G1413 (.A1(W3735), .A2(W443), .ZN(O814));
  NOR2X1 G1414 (.A1(W3138), .A2(W131), .ZN(O817));
  NOR2X1 G1415 (.A1(W3816), .A2(I596), .ZN(O818));
  NOR2X1 G1416 (.A1(I296), .A2(W2575), .ZN(W4290));
  NOR2X1 G1417 (.A1(W1047), .A2(W359), .ZN(W4293));
  NOR2X1 G1418 (.A1(W1994), .A2(W2007), .ZN(W4296));
  NOR2X1 G1419 (.A1(W1964), .A2(W2263), .ZN(W4301));
  NOR2X1 G1420 (.A1(W2268), .A2(W1002), .ZN(W4302));
  NOR2X1 G1421 (.A1(W1482), .A2(W3246), .ZN(W4304));
  NOR2X1 G1422 (.A1(W4028), .A2(W3231), .ZN(W4755));
  NOR2X1 G1423 (.A1(W2736), .A2(W2963), .ZN(O820));
  NOR2X1 G1424 (.A1(W2954), .A2(W56), .ZN(O823));
  NOR2X1 G1425 (.A1(W2859), .A2(W3575), .ZN(W4313));
  NOR2X1 G1426 (.A1(W2424), .A2(W2928), .ZN(O832));
  NOR2X1 G1427 (.A1(I849), .A2(W1095), .ZN(W4336));
  NOR2X1 G1428 (.A1(W3986), .A2(I499), .ZN(W4337));
  NOR2X1 G1429 (.A1(W1556), .A2(W564), .ZN(O835));
  NOR2X1 G1430 (.A1(W723), .A2(W3105), .ZN(W4343));
  NOR2X1 G1431 (.A1(W2201), .A2(W2627), .ZN(O838));
  NOR2X1 G1432 (.A1(W3899), .A2(W1235), .ZN(W4346));
  NOR2X1 G1433 (.A1(I38), .A2(I954), .ZN(O840));
  NOR2X1 G1434 (.A1(W4495), .A2(W4864), .ZN(O1310));
  NOR2X1 G1435 (.A1(I84), .A2(W3421), .ZN(O1287));
  NOR2X1 G1436 (.A1(W1815), .A2(W4194), .ZN(O1288));
  NOR2X1 G1437 (.A1(I907), .A2(W3172), .ZN(O1291));
  NOR2X1 G1438 (.A1(W3447), .A2(W3156), .ZN(W5136));
  NOR2X1 G1439 (.A1(W699), .A2(W3483), .ZN(O1296));
  NOR2X1 G1440 (.A1(I578), .A2(W3517), .ZN(W5141));
  NOR2X1 G1441 (.A1(W3056), .A2(I302), .ZN(W5143));
  NOR2X1 G1442 (.A1(W991), .A2(W3910), .ZN(W5144));
  NOR2X1 G1443 (.A1(W541), .A2(W2866), .ZN(O1299));
  NOR2X1 G1444 (.A1(W1651), .A2(W162), .ZN(O1304));
  NOR2X1 G1445 (.A1(W1743), .A2(W1019), .ZN(O1308));
  NOR2X1 G1446 (.A1(I909), .A2(W3970), .ZN(O1309));
  NOR2X1 G1447 (.A1(W2623), .A2(I210), .ZN(O1284));
  NOR2X1 G1448 (.A1(W2917), .A2(W2330), .ZN(O1311));
  NOR2X1 G1449 (.A1(W2891), .A2(I225), .ZN(O1313));
  NOR2X1 G1450 (.A1(W2210), .A2(W2815), .ZN(W5165));
  NOR2X1 G1451 (.A1(W3415), .A2(W848), .ZN(O1318));
  NOR2X1 G1452 (.A1(W3353), .A2(W4753), .ZN(O1321));
  NOR2X1 G1453 (.A1(W4410), .A2(W57), .ZN(O1322));
  NOR2X1 G1454 (.A1(W4977), .A2(W1741), .ZN(W5176));
  NOR2X1 G1455 (.A1(I11), .A2(W3499), .ZN(O1323));
  NOR2X1 G1456 (.A1(W1247), .A2(I960), .ZN(W5181));
  NOR2X1 G1457 (.A1(I118), .A2(W1068), .ZN(W5183));
  NOR2X1 G1458 (.A1(W4707), .A2(W1792), .ZN(W5186));
  NOR2X1 G1459 (.A1(W3605), .A2(W201), .ZN(O1329));
  NOR2X1 G1460 (.A1(W1906), .A2(W4765), .ZN(W5090));
  NOR2X1 G1461 (.A1(W492), .A2(W1605), .ZN(O1235));
  NOR2X1 G1462 (.A1(W2426), .A2(I753), .ZN(O1238));
  NOR2X1 G1463 (.A1(I430), .A2(W746), .ZN(W5062));
  NOR2X1 G1464 (.A1(W4357), .A2(W1675), .ZN(O1247));
  NOR2X1 G1465 (.A1(W3054), .A2(W1909), .ZN(W5067));
  NOR2X1 G1466 (.A1(I650), .A2(W2325), .ZN(O1251));
  NOR2X1 G1467 (.A1(W4909), .A2(W306), .ZN(W5072));
  NOR2X1 G1468 (.A1(W2854), .A2(I966), .ZN(O1253));
  NOR2X1 G1469 (.A1(W4373), .A2(W4092), .ZN(W5075));
  NOR2X1 G1470 (.A1(I391), .A2(W3086), .ZN(W5076));
  NOR2X1 G1471 (.A1(W3910), .A2(W686), .ZN(O1256));
  NOR2X1 G1472 (.A1(W2076), .A2(W629), .ZN(W5085));
  NOR2X1 G1473 (.A1(W705), .A2(W1017), .ZN(O1330));
  NOR2X1 G1474 (.A1(W2690), .A2(W1752), .ZN(O1263));
  NOR2X1 G1475 (.A1(W929), .A2(I459), .ZN(O1265));
  NOR2X1 G1476 (.A1(W1677), .A2(W3733), .ZN(O1267));
  NOR2X1 G1477 (.A1(W4797), .A2(W2334), .ZN(W5101));
  NOR2X1 G1478 (.A1(I198), .A2(W163), .ZN(O1270));
  NOR2X1 G1479 (.A1(W2624), .A2(W3747), .ZN(O1273));
  NOR2X1 G1480 (.A1(W3364), .A2(W1761), .ZN(O1278));
  NOR2X1 G1481 (.A1(W3706), .A2(W4054), .ZN(O1279));
  NOR2X1 G1482 (.A1(W2773), .A2(W2808), .ZN(O1280));
  NOR2X1 G1483 (.A1(W2295), .A2(W2127), .ZN(O1283));
  NOR2X1 G1484 (.A1(W717), .A2(W1807), .ZN(W5118));
  NOR2X1 G1485 (.A1(W3825), .A2(W1149), .ZN(O1406));
  NOR2X1 G1486 (.A1(W470), .A2(W375), .ZN(O1388));
  NOR2X1 G1487 (.A1(I508), .A2(W2630), .ZN(O1389));
  NOR2X1 G1488 (.A1(W3870), .A2(W805), .ZN(W5274));
  NOR2X1 G1489 (.A1(W2326), .A2(W1245), .ZN(O1391));
  NOR2X1 G1490 (.A1(W1045), .A2(W2529), .ZN(W5282));
  NOR2X1 G1491 (.A1(W4605), .A2(W2395), .ZN(W5283));
  NOR2X1 G1492 (.A1(W132), .A2(W319), .ZN(O1397));
  NOR2X1 G1493 (.A1(W3401), .A2(W229), .ZN(W5286));
  NOR2X1 G1494 (.A1(W1848), .A2(W3202), .ZN(O1399));
  NOR2X1 G1495 (.A1(W3773), .A2(W2760), .ZN(O1401));
  NOR2X1 G1496 (.A1(W3682), .A2(W1072), .ZN(O1404));
  NOR2X1 G1497 (.A1(W3985), .A2(W1210), .ZN(W5296));
  NOR2X1 G1498 (.A1(W2727), .A2(W2789), .ZN(O1387));
  NOR2X1 G1499 (.A1(W3588), .A2(W1057), .ZN(W5301));
  NOR2X1 G1500 (.A1(W1395), .A2(I247), .ZN(W5302));
  NOR2X1 G1501 (.A1(W3304), .A2(W1232), .ZN(O1407));
  NOR2X1 G1502 (.A1(W4144), .A2(W1691), .ZN(O1408));
  NOR2X1 G1503 (.A1(W3818), .A2(W627), .ZN(O1409));
  NOR2X1 G1504 (.A1(W962), .A2(I534), .ZN(O1410));
  NOR2X1 G1505 (.A1(W3550), .A2(I940), .ZN(O1416));
  NOR2X1 G1506 (.A1(W1316), .A2(W3814), .ZN(O1424));
  NOR2X1 G1507 (.A1(W2931), .A2(W5047), .ZN(O1427));
  NOR2X1 G1508 (.A1(W4247), .A2(W3474), .ZN(O1432));
  NOR2X1 G1509 (.A1(W1736), .A2(W3339), .ZN(O1433));
  NOR2X1 G1510 (.A1(W1834), .A2(W2241), .ZN(O1434));
  NOR2X1 G1511 (.A1(W337), .A2(W2116), .ZN(O1357));
  NOR2X1 G1512 (.A1(W3353), .A2(W151), .ZN(O1331));
  NOR2X1 G1513 (.A1(W1241), .A2(W3299), .ZN(O1333));
  NOR2X1 G1514 (.A1(W2869), .A2(W612), .ZN(O1336));
  NOR2X1 G1515 (.A1(W3077), .A2(W4454), .ZN(O1338));
  NOR2X1 G1516 (.A1(I656), .A2(W388), .ZN(O1339));
  NOR2X1 G1517 (.A1(W3947), .A2(W3544), .ZN(O1340));
  NOR2X1 G1518 (.A1(W2893), .A2(W2036), .ZN(W5206));
  NOR2X1 G1519 (.A1(W4429), .A2(W2180), .ZN(O1343));
  NOR2X1 G1520 (.A1(W1730), .A2(W3750), .ZN(W5208));
  NOR2X1 G1521 (.A1(W3847), .A2(W837), .ZN(W5218));
  NOR2X1 G1522 (.A1(W3544), .A2(W2612), .ZN(O1349));
  NOR2X1 G1523 (.A1(W54), .A2(W1919), .ZN(O1355));
  NOR2X1 G1524 (.A1(I894), .A2(W4883), .ZN(O1234));
  NOR2X1 G1525 (.A1(I904), .A2(W795), .ZN(O1359));
  NOR2X1 G1526 (.A1(I754), .A2(W4135), .ZN(O1361));
  NOR2X1 G1527 (.A1(I462), .A2(W2015), .ZN(O1362));
  NOR2X1 G1528 (.A1(W709), .A2(W2183), .ZN(O1368));
  NOR2X1 G1529 (.A1(W1470), .A2(I61), .ZN(W5250));
  NOR2X1 G1530 (.A1(I695), .A2(W994), .ZN(W5254));
  NOR2X1 G1531 (.A1(W3664), .A2(W1768), .ZN(O1374));
  NOR2X1 G1532 (.A1(W4136), .A2(W4112), .ZN(O1375));
  NOR2X1 G1533 (.A1(W1722), .A2(W2572), .ZN(O1380));
  NOR2X1 G1534 (.A1(W4630), .A2(W2803), .ZN(O1383));
  NOR2X1 G1535 (.A1(W29), .A2(W3747), .ZN(O1386));
  NOR2X1 G1536 (.A1(W207), .A2(W4368), .ZN(O1120));
  NOR2X1 G1537 (.A1(W711), .A2(W609), .ZN(O1096));
  NOR2X1 G1538 (.A1(I259), .A2(W2700), .ZN(W4824));
  NOR2X1 G1539 (.A1(W147), .A2(I81), .ZN(W4827));
  NOR2X1 G1540 (.A1(W192), .A2(I822), .ZN(W4830));
  NOR2X1 G1541 (.A1(W2616), .A2(W173), .ZN(W4833));
  NOR2X1 G1542 (.A1(I587), .A2(W2108), .ZN(O1104));
  NOR2X1 G1543 (.A1(W4184), .A2(W538), .ZN(O1110));
  NOR2X1 G1544 (.A1(W376), .A2(W348), .ZN(O1114));
  NOR2X1 G1545 (.A1(W3212), .A2(I625), .ZN(W4848));
  NOR2X1 G1546 (.A1(W2526), .A2(W3771), .ZN(W4851));
  NOR2X1 G1547 (.A1(W1335), .A2(W1869), .ZN(O1118));
  NOR2X1 G1548 (.A1(I879), .A2(W4321), .ZN(O1119));
  NOR2X1 G1549 (.A1(W457), .A2(W3129), .ZN(O1090));
  NOR2X1 G1550 (.A1(W121), .A2(W305), .ZN(O1121));
  NOR2X1 G1551 (.A1(I426), .A2(W1956), .ZN(O1122));
  NOR2X1 G1552 (.A1(W1367), .A2(W2198), .ZN(W4869));
  NOR2X1 G1553 (.A1(W2661), .A2(W178), .ZN(O1125));
  NOR2X1 G1554 (.A1(W1153), .A2(W1900), .ZN(O1129));
  NOR2X1 G1555 (.A1(W2496), .A2(W2700), .ZN(W4879));
  NOR2X1 G1556 (.A1(W2860), .A2(W1199), .ZN(W4881));
  NOR2X1 G1557 (.A1(W4745), .A2(W654), .ZN(O1132));
  NOR2X1 G1558 (.A1(W4621), .A2(I116), .ZN(O1133));
  NOR2X1 G1559 (.A1(W1110), .A2(W790), .ZN(W4889));
  NOR2X1 G1560 (.A1(W4848), .A2(W1289), .ZN(O1138));
  NOR2X1 G1561 (.A1(I690), .A2(W4624), .ZN(O1144));
  NOR2X1 G1562 (.A1(W3737), .A2(W1463), .ZN(O1068));
  NOR2X1 G1563 (.A1(W3497), .A2(W587), .ZN(O1054));
  NOR2X1 G1564 (.A1(W2706), .A2(W1668), .ZN(O1056));
  NOR2X1 G1565 (.A1(W2214), .A2(I239), .ZN(O1057));
  NOR2X1 G1566 (.A1(W1979), .A2(W1184), .ZN(W4762));
  NOR2X1 G1567 (.A1(W1067), .A2(W2284), .ZN(O1059));
  NOR2X1 G1568 (.A1(W160), .A2(W1682), .ZN(W4766));
  NOR2X1 G1569 (.A1(W1006), .A2(W9), .ZN(W4767));
  NOR2X1 G1570 (.A1(W4284), .A2(I742), .ZN(W4769));
  NOR2X1 G1571 (.A1(W2561), .A2(W4586), .ZN(O1061));
  NOR2X1 G1572 (.A1(W2893), .A2(W251), .ZN(O1062));
  NOR2X1 G1573 (.A1(I468), .A2(W3362), .ZN(O1063));
  NOR2X1 G1574 (.A1(W2793), .A2(W2567), .ZN(O1066));
  NOR2X1 G1575 (.A1(I193), .A2(W1833), .ZN(O1146));
  NOR2X1 G1576 (.A1(W227), .A2(W2004), .ZN(O1069));
  NOR2X1 G1577 (.A1(I659), .A2(W1550), .ZN(W4780));
  NOR2X1 G1578 (.A1(W371), .A2(W3484), .ZN(O1071));
  NOR2X1 G1579 (.A1(W2070), .A2(W4106), .ZN(W4783));
  NOR2X1 G1580 (.A1(I424), .A2(W1226), .ZN(W4789));
  NOR2X1 G1581 (.A1(W2666), .A2(W4131), .ZN(O1078));
  NOR2X1 G1582 (.A1(W582), .A2(W67), .ZN(W4800));
  NOR2X1 G1583 (.A1(W2785), .A2(W2891), .ZN(W4801));
  NOR2X1 G1584 (.A1(W3780), .A2(W2230), .ZN(O1086));
  NOR2X1 G1585 (.A1(W2639), .A2(W1035), .ZN(W4808));
  NOR2X1 G1586 (.A1(W2274), .A2(W3606), .ZN(W4810));
  NOR2X1 G1587 (.A1(W1145), .A2(W2272), .ZN(O1211));
  NOR2X1 G1588 (.A1(W4142), .A2(W2694), .ZN(W4985));
  NOR2X1 G1589 (.A1(W4187), .A2(W509), .ZN(O1195));
  NOR2X1 G1590 (.A1(W6), .A2(W3827), .ZN(O1196));
  NOR2X1 G1591 (.A1(W424), .A2(W3512), .ZN(O1198));
  NOR2X1 G1592 (.A1(W1827), .A2(W4631), .ZN(O1200));
  NOR2X1 G1593 (.A1(W1219), .A2(I894), .ZN(W4999));
  NOR2X1 G1594 (.A1(W1107), .A2(I558), .ZN(O1205));
  NOR2X1 G1595 (.A1(W4159), .A2(W2086), .ZN(W5005));
  NOR2X1 G1596 (.A1(W1206), .A2(W3237), .ZN(O1206));
  NOR2X1 G1597 (.A1(I294), .A2(W2777), .ZN(W5007));
  NOR2X1 G1598 (.A1(W767), .A2(I624), .ZN(W5011));
  NOR2X1 G1599 (.A1(W3581), .A2(W4377), .ZN(O1209));
  NOR2X1 G1600 (.A1(W2473), .A2(W4215), .ZN(O1193));
  NOR2X1 G1601 (.A1(W331), .A2(W1820), .ZN(O1212));
  NOR2X1 G1602 (.A1(W4394), .A2(W4243), .ZN(O1215));
  NOR2X1 G1603 (.A1(W3031), .A2(W1388), .ZN(O1216));
  NOR2X1 G1604 (.A1(W4390), .A2(W4816), .ZN(O1218));
  NOR2X1 G1605 (.A1(W3407), .A2(W4258), .ZN(O1220));
  NOR2X1 G1606 (.A1(W3534), .A2(W3074), .ZN(O1222));
  NOR2X1 G1607 (.A1(W4849), .A2(W349), .ZN(W5030));
  NOR2X1 G1608 (.A1(W2078), .A2(W2452), .ZN(W5031));
  NOR2X1 G1609 (.A1(W613), .A2(W3677), .ZN(O1224));
  NOR2X1 G1610 (.A1(W2684), .A2(W3894), .ZN(O1226));
  NOR2X1 G1611 (.A1(I436), .A2(W1086), .ZN(O1231));
  NOR2X1 G1612 (.A1(W1736), .A2(W1615), .ZN(O1232));
  NOR2X1 G1613 (.A1(W1287), .A2(I975), .ZN(O1166));
  NOR2X1 G1614 (.A1(W3879), .A2(W4140), .ZN(O1147));
  NOR2X1 G1615 (.A1(I546), .A2(W4423), .ZN(O1148));
  NOR2X1 G1616 (.A1(W2007), .A2(W723), .ZN(O1149));
  NOR2X1 G1617 (.A1(W689), .A2(W481), .ZN(O1150));
  NOR2X1 G1618 (.A1(I940), .A2(W1649), .ZN(W4916));
  NOR2X1 G1619 (.A1(W319), .A2(I38), .ZN(W4918));
  NOR2X1 G1620 (.A1(W3748), .A2(I27), .ZN(O1156));
  NOR2X1 G1621 (.A1(W4904), .A2(I815), .ZN(O1163));
  NOR2X1 G1622 (.A1(W214), .A2(W3068), .ZN(W4934));
  NOR2X1 G1623 (.A1(W3715), .A2(W1845), .ZN(W4935));
  NOR2X1 G1624 (.A1(I846), .A2(I682), .ZN(W4938));
  NOR2X1 G1625 (.A1(W2642), .A2(W1580), .ZN(W4939));
  NOR2X1 G1626 (.A1(W326), .A2(W2969), .ZN(W3251));
  NOR2X1 G1627 (.A1(W3812), .A2(I683), .ZN(O1175));
  NOR2X1 G1628 (.A1(W4271), .A2(W2100), .ZN(O1181));
  NOR2X1 G1629 (.A1(W1469), .A2(W2832), .ZN(W4962));
  NOR2X1 G1630 (.A1(I342), .A2(W2356), .ZN(W4964));
  NOR2X1 G1631 (.A1(W3776), .A2(W1984), .ZN(W4969));
  NOR2X1 G1632 (.A1(I572), .A2(W821), .ZN(O1185));
  NOR2X1 G1633 (.A1(W1670), .A2(W1718), .ZN(O1186));
  NOR2X1 G1634 (.A1(W3192), .A2(W3206), .ZN(O1189));
  NOR2X1 G1635 (.A1(W215), .A2(W4264), .ZN(W4977));
  NOR2X1 G1636 (.A1(W944), .A2(W624), .ZN(O1191));
  NOR2X1 G1637 (.A1(I716), .A2(W3100), .ZN(O1192));
  NOR2X1 G1638 (.A1(I34), .A2(W721), .ZN(W790));
  NOR2X1 G1639 (.A1(I315), .A2(W244), .ZN(W797));
  NOR2X1 G1640 (.A1(W1223), .A2(W1093), .ZN(W1427));
  NOR2X1 G1641 (.A1(W655), .A2(W491), .ZN(W1147));
  NOR2X1 G1642 (.A1(I152), .A2(W1104), .ZN(W1426));
  NOR2X1 G1643 (.A1(I658), .A2(I659), .ZN(W329));
  NOR2X1 G1644 (.A1(I12), .A2(W891), .ZN(W1149));
  NOR2X1 G1645 (.A1(I668), .A2(I669), .ZN(W334));
  NOR2X1 G1646 (.A1(I670), .A2(I671), .ZN(W335));
  NOR2X1 G1647 (.A1(I672), .A2(I673), .ZN(W336));
  NOR2X1 G1648 (.A1(I674), .A2(I675), .ZN(W337));
  NOR2X1 G1649 (.A1(I676), .A2(I677), .ZN(W338));
  NOR2X1 G1650 (.A1(I648), .A2(I649), .ZN(W324));
  NOR2X1 G1651 (.A1(I678), .A2(I679), .ZN(W339));
  NOR2X1 G1652 (.A1(W348), .A2(W1018), .ZN(O65));
  NOR2X1 G1653 (.A1(I680), .A2(I681), .ZN(W340));
  NOR2X1 G1654 (.A1(I682), .A2(I683), .ZN(W341));
  NOR2X1 G1655 (.A1(W754), .A2(W293), .ZN(W1418));
  NOR2X1 G1656 (.A1(I452), .A2(W958), .ZN(W1154));
  NOR2X1 G1657 (.A1(W267), .A2(W36), .ZN(W1416));
  NOR2X1 G1658 (.A1(I42), .A2(I759), .ZN(W788));
  NOR2X1 G1659 (.A1(W109), .A2(W745), .ZN(W787));
  NOR2X1 G1660 (.A1(W104), .A2(I414), .ZN(W1414));
  NOR2X1 G1661 (.A1(I694), .A2(I695), .ZN(W347));
  NOR2X1 G1662 (.A1(W1249), .A2(W62), .ZN(W1433));
  NOR2X1 G1663 (.A1(I614), .A2(I615), .ZN(W307));
  NOR2X1 G1664 (.A1(I618), .A2(I619), .ZN(W309));
  NOR2X1 G1665 (.A1(W1313), .A2(I217), .ZN(W1436));
  NOR2X1 G1666 (.A1(I620), .A2(I621), .ZN(W310));
  NOR2X1 G1667 (.A1(I624), .A2(I625), .ZN(W312));
  NOR2X1 G1668 (.A1(W457), .A2(W798), .ZN(W1434));
  NOR2X1 G1669 (.A1(I628), .A2(I629), .ZN(W314));
  NOR2X1 G1670 (.A1(W86), .A2(W362), .ZN(W801));
  NOR2X1 G1671 (.A1(I630), .A2(I631), .ZN(W315));
  NOR2X1 G1672 (.A1(I632), .A2(I633), .ZN(W316));
  NOR2X1 G1673 (.A1(I191), .A2(I206), .ZN(W799));
  NOR2X1 G1674 (.A1(W1134), .A2(W696), .ZN(W1411));
  NOR2X1 G1675 (.A1(W184), .A2(W200), .ZN(W798));
  NOR2X1 G1676 (.A1(W920), .A2(W375), .ZN(O66));
  NOR2X1 G1677 (.A1(I634), .A2(I635), .ZN(O4));
  NOR2X1 G1678 (.A1(W985), .A2(W364), .ZN(W1143));
  NOR2X1 G1679 (.A1(I636), .A2(I637), .ZN(W318));
  NOR2X1 G1680 (.A1(I638), .A2(I639), .ZN(W319));
  NOR2X1 G1681 (.A1(W774), .A2(W843), .ZN(W1430));
  NOR2X1 G1682 (.A1(I640), .A2(I641), .ZN(W320));
  NOR2X1 G1683 (.A1(W998), .A2(W273), .ZN(W1145));
  NOR2X1 G1684 (.A1(I646), .A2(I647), .ZN(W323));
  NOR2X1 G1685 (.A1(W396), .A2(W486), .ZN(W1392));
  NOR2X1 G1686 (.A1(I744), .A2(I745), .ZN(W372));
  NOR2X1 G1687 (.A1(W535), .A2(I106), .ZN(W772));
  NOR2X1 G1688 (.A1(W860), .A2(W305), .ZN(W1397));
  NOR2X1 G1689 (.A1(W1278), .A2(I490), .ZN(W1396));
  NOR2X1 G1690 (.A1(I752), .A2(I753), .ZN(W376));
  NOR2X1 G1691 (.A1(I996), .A2(W114), .ZN(W771));
  NOR2X1 G1692 (.A1(W1041), .A2(W50), .ZN(W1168));
  NOR2X1 G1693 (.A1(W41), .A2(I6), .ZN(W770));
  NOR2X1 G1694 (.A1(I764), .A2(I765), .ZN(W382));
  NOR2X1 G1695 (.A1(I766), .A2(I767), .ZN(W383));
  NOR2X1 G1696 (.A1(W489), .A2(W675), .ZN(W768));
  NOR2X1 G1697 (.A1(I247), .A2(I252), .ZN(W774));
  NOR2X1 G1698 (.A1(I776), .A2(I777), .ZN(W388));
  NOR2X1 G1699 (.A1(I778), .A2(I779), .ZN(W389));
  NOR2X1 G1700 (.A1(I780), .A2(I781), .ZN(W390));
  NOR2X1 G1701 (.A1(I898), .A2(W1387), .ZN(W1389));
  NOR2X1 G1702 (.A1(W208), .A2(I580), .ZN(W1173));
  NOR2X1 G1703 (.A1(I784), .A2(I785), .ZN(W392));
  NOR2X1 G1704 (.A1(I786), .A2(I787), .ZN(W393));
  NOR2X1 G1705 (.A1(I298), .A2(W597), .ZN(W1178));
  NOR2X1 G1706 (.A1(I790), .A2(I791), .ZN(W395));
  NOR2X1 G1707 (.A1(I792), .A2(I793), .ZN(W396));
  NOR2X1 G1708 (.A1(W393), .A2(I915), .ZN(W757));
  NOR2X1 G1709 (.A1(I525), .A2(W170), .ZN(W1401));
  NOR2X1 G1710 (.A1(W59), .A2(I754), .ZN(W1410));
  NOR2X1 G1711 (.A1(I700), .A2(I701), .ZN(W350));
  NOR2X1 G1712 (.A1(I705), .A2(W772), .ZN(W1409));
  NOR2X1 G1713 (.A1(W739), .A2(I890), .ZN(W784));
  NOR2X1 G1714 (.A1(I706), .A2(I707), .ZN(W353));
  NOR2X1 G1715 (.A1(W447), .A2(W556), .ZN(W781));
  NOR2X1 G1716 (.A1(I710), .A2(I711), .ZN(W355));
  NOR2X1 G1717 (.A1(I712), .A2(I713), .ZN(W356));
  NOR2X1 G1718 (.A1(I531), .A2(I711), .ZN(W1404));
  NOR2X1 G1719 (.A1(I7), .A2(W778), .ZN(W1159));
  NOR2X1 G1720 (.A1(W821), .A2(I160), .ZN(W1160));
  NOR2X1 G1721 (.A1(I612), .A2(I613), .ZN(W306));
  NOR2X1 G1722 (.A1(I722), .A2(I723), .ZN(W361));
  NOR2X1 G1723 (.A1(I126), .A2(W781), .ZN(W1163));
  NOR2X1 G1724 (.A1(I724), .A2(I725), .ZN(W362));
  NOR2X1 G1725 (.A1(I726), .A2(I727), .ZN(W363));
  NOR2X1 G1726 (.A1(I728), .A2(I729), .ZN(W364));
  NOR2X1 G1727 (.A1(I730), .A2(I731), .ZN(W365));
  NOR2X1 G1728 (.A1(I590), .A2(I92), .ZN(W778));
  NOR2X1 G1729 (.A1(W600), .A2(W478), .ZN(W777));
  NOR2X1 G1730 (.A1(W729), .A2(I391), .ZN(W1166));
  NOR2X1 G1731 (.A1(I736), .A2(I737), .ZN(W368));
  NOR2X1 G1732 (.A1(I744), .A2(W485), .ZN(W853));
  NOR2X1 G1733 (.A1(I134), .A2(I794), .ZN(O71));
  NOR2X1 G1734 (.A1(I598), .A2(W741), .ZN(W1109));
  NOR2X1 G1735 (.A1(I462), .A2(I463), .ZN(W231));
  NOR2X1 G1736 (.A1(I728), .A2(I640), .ZN(W1110));
  NOR2X1 G1737 (.A1(I134), .A2(I43), .ZN(W860));
  NOR2X1 G1738 (.A1(W659), .A2(I552), .ZN(W1488));
  NOR2X1 G1739 (.A1(I911), .A2(W203), .ZN(W1112));
  NOR2X1 G1740 (.A1(I466), .A2(I467), .ZN(W233));
  NOR2X1 G1741 (.A1(I451), .A2(W676), .ZN(W857));
  NOR2X1 G1742 (.A1(I468), .A2(I469), .ZN(W234));
  NOR2X1 G1743 (.A1(I219), .A2(W313), .ZN(W856));
  NOR2X1 G1744 (.A1(I537), .A2(I431), .ZN(W1108));
  NOR2X1 G1745 (.A1(W158), .A2(I460), .ZN(W850));
  NOR2X1 G1746 (.A1(W721), .A2(W447), .ZN(W1482));
  NOR2X1 G1747 (.A1(W1009), .A2(W781), .ZN(W1481));
  NOR2X1 G1748 (.A1(I480), .A2(I481), .ZN(W240));
  NOR2X1 G1749 (.A1(I170), .A2(I11), .ZN(O69));
  NOR2X1 G1750 (.A1(I484), .A2(I485), .ZN(W242));
  NOR2X1 G1751 (.A1(I685), .A2(W370), .ZN(O30));
  NOR2X1 G1752 (.A1(W506), .A2(I620), .ZN(W845));
  NOR2X1 G1753 (.A1(I661), .A2(I992), .ZN(W1119));
  NOR2X1 G1754 (.A1(I610), .A2(W886), .ZN(W1474));
  NOR2X1 G1755 (.A1(I492), .A2(I493), .ZN(W246));
  NOR2X1 G1756 (.A1(I444), .A2(I445), .ZN(W222));
  NOR2X1 G1757 (.A1(I646), .A2(I542), .ZN(W886));
  NOR2X1 G1758 (.A1(W170), .A2(I636), .ZN(W1505));
  NOR2X1 G1759 (.A1(I420), .A2(I421), .ZN(W210));
  NOR2X1 G1760 (.A1(W737), .A2(W1025), .ZN(W1096));
  NOR2X1 G1761 (.A1(W773), .A2(I64), .ZN(W1504));
  NOR2X1 G1762 (.A1(W692), .A2(W431), .ZN(W1098));
  NOR2X1 G1763 (.A1(I430), .A2(I431), .ZN(W215));
  NOR2X1 G1764 (.A1(W1391), .A2(I276), .ZN(W1503));
  NOR2X1 G1765 (.A1(I434), .A2(I435), .ZN(W217));
  NOR2X1 G1766 (.A1(I440), .A2(I441), .ZN(W220));
  NOR2X1 G1767 (.A1(I442), .A2(I443), .ZN(W221));
  NOR2X1 G1768 (.A1(I494), .A2(I495), .ZN(W247));
  NOR2X1 G1769 (.A1(I446), .A2(I447), .ZN(W223));
  NOR2X1 G1770 (.A1(I336), .A2(W319), .ZN(O45));
  NOR2X1 G1771 (.A1(I469), .A2(I111), .ZN(W867));
  NOR2X1 G1772 (.A1(I485), .A2(I511), .ZN(W1498));
  NOR2X1 G1773 (.A1(W1229), .A2(I605), .ZN(W1497));
  NOR2X1 G1774 (.A1(W1109), .A2(W1261), .ZN(W1496));
  NOR2X1 G1775 (.A1(I454), .A2(I455), .ZN(W227));
  NOR2X1 G1776 (.A1(W226), .A2(W188), .ZN(W1107));
  NOR2X1 G1777 (.A1(I206), .A2(I700), .ZN(W866));
  NOR2X1 G1778 (.A1(I458), .A2(I459), .ZN(W229));
  NOR2X1 G1779 (.A1(I64), .A2(I421), .ZN(O46));
  NOR2X1 G1780 (.A1(I558), .A2(I559), .ZN(W279));
  NOR2X1 G1781 (.A1(W16), .A2(W153), .ZN(W821));
  NOR2X1 G1782 (.A1(I562), .A2(I563), .ZN(W281));
  NOR2X1 G1783 (.A1(I566), .A2(I567), .ZN(W283));
  NOR2X1 G1784 (.A1(W402), .A2(I470), .ZN(W1129));
  NOR2X1 G1785 (.A1(W1118), .A2(I596), .ZN(W1130));
  NOR2X1 G1786 (.A1(W1361), .A2(I748), .ZN(W1449));
  NOR2X1 G1787 (.A1(I578), .A2(I579), .ZN(W289));
  NOR2X1 G1788 (.A1(I421), .A2(W736), .ZN(W1448));
  NOR2X1 G1789 (.A1(I631), .A2(I678), .ZN(W1447));
  NOR2X1 G1790 (.A1(I582), .A2(I583), .ZN(W291));
  NOR2X1 G1791 (.A1(I556), .A2(I557), .ZN(W278));
  NOR2X1 G1792 (.A1(I704), .A2(W486), .ZN(W811));
  NOR2X1 G1793 (.A1(W1116), .A2(I385), .ZN(W1445));
  NOR2X1 G1794 (.A1(I836), .A2(I147), .ZN(W1135));
  NOR2X1 G1795 (.A1(W94), .A2(I64), .ZN(W1442));
  NOR2X1 G1796 (.A1(W257), .A2(W1057), .ZN(W1137));
  NOR2X1 G1797 (.A1(W1028), .A2(W626), .ZN(W1441));
  NOR2X1 G1798 (.A1(W399), .A2(I697), .ZN(W808));
  NOR2X1 G1799 (.A1(I445), .A2(I80), .ZN(W806));
  NOR2X1 G1800 (.A1(I606), .A2(I607), .ZN(W303));
  NOR2X1 G1801 (.A1(W116), .A2(W188), .ZN(W804));
  NOR2X1 G1802 (.A1(I524), .A2(I525), .ZN(W262));
  NOR2X1 G1803 (.A1(W894), .A2(I866), .ZN(W1122));
  NOR2X1 G1804 (.A1(I252), .A2(W300), .ZN(W1123));
  NOR2X1 G1805 (.A1(I794), .A2(W472), .ZN(W838));
  NOR2X1 G1806 (.A1(I510), .A2(I511), .ZN(W255));
  NOR2X1 G1807 (.A1(W209), .A2(I963), .ZN(W837));
  NOR2X1 G1808 (.A1(I248), .A2(I196), .ZN(W835));
  NOR2X1 G1809 (.A1(I516), .A2(I517), .ZN(W258));
  NOR2X1 G1810 (.A1(W206), .A2(W506), .ZN(W1128));
  NOR2X1 G1811 (.A1(I518), .A2(I519), .ZN(W259));
  NOR2X1 G1812 (.A1(I930), .A2(I877), .ZN(O68));
  NOR2X1 G1813 (.A1(I520), .A2(I521), .ZN(W260));
  NOR2X1 G1814 (.A1(I808), .A2(I809), .ZN(W404));
  NOR2X1 G1815 (.A1(I526), .A2(I527), .ZN(W263));
  NOR2X1 G1816 (.A1(I530), .A2(I531), .ZN(W265));
  NOR2X1 G1817 (.A1(I538), .A2(I539), .ZN(W269));
  NOR2X1 G1818 (.A1(I819), .A2(I283), .ZN(W1460));
  NOR2X1 G1819 (.A1(I540), .A2(I541), .ZN(W270));
  NOR2X1 G1820 (.A1(I546), .A2(I547), .ZN(W273));
  NOR2X1 G1821 (.A1(W1256), .A2(W475), .ZN(W1458));
  NOR2X1 G1822 (.A1(I548), .A2(I549), .ZN(W274));
  NOR2X1 G1823 (.A1(I550), .A2(I551), .ZN(W275));
  NOR2X1 G1824 (.A1(I554), .A2(I555), .ZN(W277));
  NOR2X1 G1825 (.A1(I437), .A2(I815), .ZN(W665));
  NOR2X1 G1826 (.A1(W242), .A2(I517), .ZN(W542));
  NOR2X1 G1827 (.A1(W248), .A2(W441), .ZN(O56));
  NOR2X1 G1828 (.A1(I437), .A2(I443), .ZN(W1239));
  NOR2X1 G1829 (.A1(W548), .A2(W383), .ZN(W1311));
  NOR2X1 G1830 (.A1(I16), .A2(I863), .ZN(W546));
  NOR2X1 G1831 (.A1(I103), .A2(I568), .ZN(W668));
  NOR2X1 G1832 (.A1(W156), .A2(I124), .ZN(O61));
  NOR2X1 G1833 (.A1(I5), .A2(I27), .ZN(W547));
  NOR2X1 G1834 (.A1(I747), .A2(I209), .ZN(W548));
  NOR2X1 G1835 (.A1(W79), .A2(I735), .ZN(W667));
  NOR2X1 G1836 (.A1(W300), .A2(I120), .ZN(W666));
  NOR2X1 G1837 (.A1(W347), .A2(W235), .ZN(W541));
  NOR2X1 G1838 (.A1(W1255), .A2(W510), .ZN(W1305));
  NOR2X1 G1839 (.A1(W150), .A2(I108), .ZN(W664));
  NOR2X1 G1840 (.A1(W222), .A2(I243), .ZN(W663));
  NOR2X1 G1841 (.A1(W399), .A2(I14), .ZN(W550));
  NOR2X1 G1842 (.A1(I206), .A2(W1179), .ZN(W1302));
  NOR2X1 G1843 (.A1(W334), .A2(I923), .ZN(W657));
  NOR2X1 G1844 (.A1(W478), .A2(I423), .ZN(W655));
  NOR2X1 G1845 (.A1(I925), .A2(W325), .ZN(W1301));
  NOR2X1 G1846 (.A1(W835), .A2(W1233), .ZN(W1300));
  NOR2X1 G1847 (.A1(W732), .A2(I21), .ZN(W1299));
  NOR2X1 G1848 (.A1(I330), .A2(I495), .ZN(W653));
  NOR2X1 G1849 (.A1(I746), .A2(W269), .ZN(W527));
  NOR2X1 G1850 (.A1(W258), .A2(I811), .ZN(W515));
  NOR2X1 G1851 (.A1(W250), .A2(W678), .ZN(W1229));
  NOR2X1 G1852 (.A1(W1151), .A2(W511), .ZN(W1230));
  NOR2X1 G1853 (.A1(W443), .A2(W209), .ZN(W520));
  NOR2X1 G1854 (.A1(W320), .A2(W363), .ZN(W1319));
  NOR2X1 G1855 (.A1(I584), .A2(I416), .ZN(W521));
  NOR2X1 G1856 (.A1(I969), .A2(I305), .ZN(W523));
  NOR2X1 G1857 (.A1(I481), .A2(W2), .ZN(W524));
  NOR2X1 G1858 (.A1(I88), .A2(W182), .ZN(W525));
  NOR2X1 G1859 (.A1(I646), .A2(I679), .ZN(W678));
  NOR2X1 G1860 (.A1(I894), .A2(I842), .ZN(O21));
  NOR2X1 G1861 (.A1(I993), .A2(I356), .ZN(W652));
  NOR2X1 G1862 (.A1(W30), .A2(W582), .ZN(W676));
  NOR2X1 G1863 (.A1(W627), .A2(I919), .ZN(W1234));
  NOR2X1 G1864 (.A1(W450), .A2(I168), .ZN(W675));
  NOR2X1 G1865 (.A1(I584), .A2(I357), .ZN(W673));
  NOR2X1 G1866 (.A1(W349), .A2(I72), .ZN(W535));
  NOR2X1 G1867 (.A1(W765), .A2(I57), .ZN(W1237));
  NOR2X1 G1868 (.A1(I973), .A2(W180), .ZN(W672));
  NOR2X1 G1869 (.A1(W382), .A2(I814), .ZN(W538));
  NOR2X1 G1870 (.A1(I448), .A2(I260), .ZN(W539));
  NOR2X1 G1871 (.A1(I846), .A2(I250), .ZN(W670));
  NOR2X1 G1872 (.A1(W800), .A2(W1150), .ZN(W1280));
  NOR2X1 G1873 (.A1(W560), .A2(I470), .ZN(O17));
  NOR2X1 G1874 (.A1(I710), .A2(W169), .ZN(W642));
  NOR2X1 G1875 (.A1(I714), .A2(W371), .ZN(W641));
  NOR2X1 G1876 (.A1(W377), .A2(I200), .ZN(W582));
  NOR2X1 G1877 (.A1(I613), .A2(I168), .ZN(W639));
  NOR2X1 G1878 (.A1(I600), .A2(W39), .ZN(W633));
  NOR2X1 G1879 (.A1(W386), .A2(W481), .ZN(W1259));
  NOR2X1 G1880 (.A1(I686), .A2(I746), .ZN(W1283));
  NOR2X1 G1881 (.A1(I853), .A2(W225), .ZN(W632));
  NOR2X1 G1882 (.A1(W963), .A2(W1092), .ZN(W1281));
  NOR2X1 G1883 (.A1(I800), .A2(W1103), .ZN(W1261));
  NOR2X1 G1884 (.A1(W127), .A2(W136), .ZN(W574));
  NOR2X1 G1885 (.A1(W45), .A2(W580), .ZN(W590));
  NOR2X1 G1886 (.A1(W121), .A2(I967), .ZN(W591));
  NOR2X1 G1887 (.A1(W408), .A2(W103), .ZN(W623));
  NOR2X1 G1888 (.A1(W162), .A2(I157), .ZN(W622));
  NOR2X1 G1889 (.A1(I936), .A2(I152), .ZN(W596));
  NOR2X1 G1890 (.A1(W291), .A2(I941), .ZN(W1265));
  NOR2X1 G1891 (.A1(W114), .A2(I320), .ZN(W606));
  NOR2X1 G1892 (.A1(W6), .A2(I909), .ZN(W613));
  NOR2X1 G1893 (.A1(I342), .A2(W110), .ZN(W1267));
  NOR2X1 G1894 (.A1(W1186), .A2(I724), .ZN(W1270));
  NOR2X1 G1895 (.A1(W156), .A2(I944), .ZN(W617));
  NOR2X1 G1896 (.A1(W438), .A2(I734), .ZN(W1253));
  NOR2X1 G1897 (.A1(I508), .A2(W537), .ZN(W651));
  NOR2X1 G1898 (.A1(I504), .A2(W1084), .ZN(W1247));
  NOR2X1 G1899 (.A1(W294), .A2(I349), .ZN(W561));
  NOR2X1 G1900 (.A1(W465), .A2(W352), .ZN(W562));
  NOR2X1 G1901 (.A1(W521), .A2(W45), .ZN(W650));
  NOR2X1 G1902 (.A1(W623), .A2(I548), .ZN(W1249));
  NOR2X1 G1903 (.A1(W439), .A2(W240), .ZN(W1250));
  NOR2X1 G1904 (.A1(I970), .A2(W250), .ZN(W649));
  NOR2X1 G1905 (.A1(I509), .A2(W296), .ZN(W647));
  NOR2X1 G1906 (.A1(I861), .A2(W352), .ZN(W565));
  NOR2X1 G1907 (.A1(I457), .A2(I452), .ZN(W646));
  NOR2X1 G1908 (.A1(I486), .A2(W272), .ZN(W1324));
  NOR2X1 G1909 (.A1(W303), .A2(W264), .ZN(W644));
  NOR2X1 G1910 (.A1(I4), .A2(I996), .ZN(W567));
  NOR2X1 G1911 (.A1(W145), .A2(W393), .ZN(W1291));
  NOR2X1 G1912 (.A1(W429), .A2(I764), .ZN(W643));
  NOR2X1 G1913 (.A1(I136), .A2(I19), .ZN(W569));
  NOR2X1 G1914 (.A1(I457), .A2(I601), .ZN(W570));
  NOR2X1 G1915 (.A1(I649), .A2(I760), .ZN(W571));
  NOR2X1 G1916 (.A1(W62), .A2(W629), .ZN(W1289));
  NOR2X1 G1917 (.A1(W1104), .A2(W491), .ZN(W1288));
  NOR2X1 G1918 (.A1(W339), .A2(I297), .ZN(W573));
  NOR2X1 G1919 (.A1(W1090), .A2(W1169), .ZN(W1363));
  NOR2X1 G1920 (.A1(I862), .A2(I863), .ZN(W431));
  NOR2X1 G1921 (.A1(I870), .A2(I871), .ZN(O9));
  NOR2X1 G1922 (.A1(I244), .A2(W164), .ZN(W1369));
  NOR2X1 G1923 (.A1(I974), .A2(I422), .ZN(W1368));
  NOR2X1 G1924 (.A1(I874), .A2(I875), .ZN(W437));
  NOR2X1 G1925 (.A1(W257), .A2(I365), .ZN(W739));
  NOR2X1 G1926 (.A1(W612), .A2(I568), .ZN(O52));
  NOR2X1 G1927 (.A1(I880), .A2(I881), .ZN(W440));
  NOR2X1 G1928 (.A1(I884), .A2(I885), .ZN(W442));
  NOR2X1 G1929 (.A1(I299), .A2(I365), .ZN(W735));
  NOR2X1 G1930 (.A1(I223), .A2(I5), .ZN(W1364));
  NOR2X1 G1931 (.A1(I860), .A2(I861), .ZN(W430));
  NOR2X1 G1932 (.A1(I760), .A2(I22), .ZN(W734));
  NOR2X1 G1933 (.A1(I853), .A2(I113), .ZN(W733));
  NOR2X1 G1934 (.A1(I499), .A2(I200), .ZN(W732));
  NOR2X1 G1935 (.A1(I888), .A2(I889), .ZN(W444));
  NOR2X1 G1936 (.A1(I894), .A2(I895), .ZN(W447));
  NOR2X1 G1937 (.A1(I450), .A2(W529), .ZN(W730));
  NOR2X1 G1938 (.A1(I922), .A2(W250), .ZN(W1356));
  NOR2X1 G1939 (.A1(W496), .A2(I694), .ZN(W723));
  NOR2X1 G1940 (.A1(I908), .A2(I909), .ZN(W454));
  NOR2X1 G1941 (.A1(I910), .A2(I911), .ZN(O11));
  NOR2X1 G1942 (.A1(I912), .A2(I913), .ZN(O12));
  NOR2X1 G1943 (.A1(W346), .A2(I854), .ZN(W750));
  NOR2X1 G1944 (.A1(W473), .A2(W361), .ZN(O25));
  NOR2X1 G1945 (.A1(I814), .A2(I815), .ZN(W407));
  NOR2X1 G1946 (.A1(I816), .A2(I817), .ZN(W408));
  NOR2X1 G1947 (.A1(I818), .A2(I819), .ZN(W409));
  NOR2X1 G1948 (.A1(W1172), .A2(I145), .ZN(W1185));
  NOR2X1 G1949 (.A1(W548), .A2(W978), .ZN(W1186));
  NOR2X1 G1950 (.A1(I824), .A2(I825), .ZN(W412));
  NOR2X1 G1951 (.A1(W971), .A2(W832), .ZN(W1381));
  NOR2X1 G1952 (.A1(I830), .A2(I831), .ZN(W415));
  NOR2X1 G1953 (.A1(W231), .A2(I679), .ZN(W1379));
  NOR2X1 G1954 (.A1(W969), .A2(W617), .ZN(W1189));
  NOR2X1 G1955 (.A1(I914), .A2(I915), .ZN(W457));
  NOR2X1 G1956 (.A1(I196), .A2(I50), .ZN(W749));
  NOR2X1 G1957 (.A1(I832), .A2(I833), .ZN(W416));
  NOR2X1 G1958 (.A1(W499), .A2(W443), .ZN(W748));
  NOR2X1 G1959 (.A1(W1357), .A2(I581), .ZN(W1374));
  NOR2X1 G1960 (.A1(I838), .A2(I839), .ZN(W419));
  NOR2X1 G1961 (.A1(W865), .A2(I213), .ZN(O64));
  NOR2X1 G1962 (.A1(I687), .A2(I628), .ZN(W1192));
  NOR2X1 G1963 (.A1(I852), .A2(I853), .ZN(W426));
  NOR2X1 G1964 (.A1(I856), .A2(I857), .ZN(W428));
  NOR2X1 G1965 (.A1(I858), .A2(I859), .ZN(W429));
  NOR2X1 G1966 (.A1(I662), .A2(W149), .ZN(W505));
  NOR2X1 G1967 (.A1(I195), .A2(W252), .ZN(O22));
  NOR2X1 G1968 (.A1(W1303), .A2(W1066), .ZN(W1332));
  NOR2X1 G1969 (.A1(I988), .A2(I989), .ZN(W494));
  NOR2X1 G1970 (.A1(I990), .A2(I991), .ZN(W495));
  NOR2X1 G1971 (.A1(I998), .A2(I999), .ZN(W499));
  NOR2X1 G1972 (.A1(I794), .A2(W123), .ZN(W698));
  NOR2X1 G1973 (.A1(I446), .A2(W103), .ZN(W500));
  NOR2X1 G1974 (.A1(I829), .A2(I726), .ZN(W697));
  NOR2X1 G1975 (.A1(I687), .A2(W163), .ZN(W695));
  NOR2X1 G1976 (.A1(W549), .A2(W110), .ZN(W1329));
  NOR2X1 G1977 (.A1(I23), .A2(I563), .ZN(W504));
  NOR2X1 G1978 (.A1(W379), .A2(I388), .ZN(W1333));
  NOR2X1 G1979 (.A1(W678), .A2(I284), .ZN(W692));
  NOR2X1 G1980 (.A1(I824), .A2(I688), .ZN(W508));
  NOR2X1 G1981 (.A1(I375), .A2(I766), .ZN(W689));
  NOR2X1 G1982 (.A1(W427), .A2(W1138), .ZN(W1225));
  NOR2X1 G1983 (.A1(I862), .A2(W222), .ZN(W688));
  NOR2X1 G1984 (.A1(I259), .A2(I674), .ZN(W511));
  NOR2X1 G1985 (.A1(W139), .A2(W3), .ZN(W512));
  NOR2X1 G1986 (.A1(I42), .A2(W423), .ZN(W513));
  NOR2X1 G1987 (.A1(W342), .A2(W995), .ZN(W1226));
  NOR2X1 G1988 (.A1(I204), .A2(W566), .ZN(W1227));
  NOR2X1 G1989 (.A1(W1214), .A2(I730), .ZN(W1345));
  NOR2X1 G1990 (.A1(I390), .A2(W117), .ZN(W1206));
  NOR2X1 G1991 (.A1(I916), .A2(I917), .ZN(W458));
  NOR2X1 G1992 (.A1(I415), .A2(I396), .ZN(W1207));
  NOR2X1 G1993 (.A1(W687), .A2(I437), .ZN(O23));
  NOR2X1 G1994 (.A1(I236), .A2(W674), .ZN(W1209));
  NOR2X1 G1995 (.A1(I922), .A2(I923), .ZN(W461));
  NOR2X1 G1996 (.A1(I924), .A2(I925), .ZN(W462));
  NOR2X1 G1997 (.A1(I458), .A2(W510), .ZN(W718));
  NOR2X1 G1998 (.A1(I928), .A2(I929), .ZN(W464));
  NOR2X1 G1999 (.A1(I936), .A2(I937), .ZN(W468));
  NOR2X1 G2000 (.A1(I942), .A2(I943), .ZN(W471));
  NOR2X1 G2001 (.A1(W232), .A2(I413), .ZN(W1438));
  NOR2X1 G2002 (.A1(W51), .A2(W903), .ZN(W1213));
  NOR2X1 G2003 (.A1(W517), .A2(I784), .ZN(W1214));
  NOR2X1 G2004 (.A1(I956), .A2(I957), .ZN(W478));
  NOR2X1 G2005 (.A1(W651), .A2(W439), .ZN(W715));
  NOR2X1 G2006 (.A1(I968), .A2(I969), .ZN(W484));
  NOR2X1 G2007 (.A1(W959), .A2(I716), .ZN(W1339));
  NOR2X1 G2008 (.A1(I974), .A2(I975), .ZN(W487));
  NOR2X1 G2009 (.A1(W482), .A2(I466), .ZN(W1336));
  NOR2X1 G2010 (.A1(I590), .A2(I894), .ZN(W1335));
  NOR2X1 G2011 (.A1(I982), .A2(I983), .ZN(W491));
  NOR2X1 G2012 (.A1(I530), .A2(W87), .ZN(W1565));
  NOR2X1 G2013 (.A1(I416), .A2(I417), .ZN(W208));
  NOR2X1 G2014 (.A1(W114), .A2(I715), .ZN(W955));
  NOR2X1 G2015 (.A1(I356), .A2(W662), .ZN(W954));
  NOR2X1 G2016 (.A1(W975), .A2(W674), .ZN(W1046));
  NOR2X1 G2017 (.A1(W1082), .A2(I579), .ZN(W1570));
  NOR2X1 G2018 (.A1(I230), .A2(I231), .ZN(W115));
  NOR2X1 G2019 (.A1(I76), .A2(W573), .ZN(W1047));
  NOR2X1 G2020 (.A1(I234), .A2(I235), .ZN(W117));
  NOR2X1 G2021 (.A1(W640), .A2(I166), .ZN(W1566));
  NOR2X1 G2022 (.A1(I224), .A2(I225), .ZN(W112));
  NOR2X1 G2023 (.A1(I546), .A2(I572), .ZN(W1048));
  NOR2X1 G2024 (.A1(I240), .A2(I241), .ZN(W120));
  NOR2X1 G2025 (.A1(W287), .A2(I208), .ZN(W1049));
  NOR2X1 G2026 (.A1(W941), .A2(W568), .ZN(W948));
  NOR2X1 G2027 (.A1(I244), .A2(I245), .ZN(W122));
  NOR2X1 G2028 (.A1(W856), .A2(W1436), .ZN(W1562));
  NOR2X1 G2029 (.A1(W409), .A2(W1181), .ZN(W1561));
  NOR2X1 G2030 (.A1(I246), .A2(I247), .ZN(W123));
  NOR2X1 G2031 (.A1(I248), .A2(I249), .ZN(W124));
  NOR2X1 G2032 (.A1(W596), .A2(W217), .ZN(W961));
  NOR2X1 G2033 (.A1(I178), .A2(I179), .ZN(W89));
  NOR2X1 G2034 (.A1(I180), .A2(I181), .ZN(W90));
  NOR2X1 G2035 (.A1(I184), .A2(I185), .ZN(W92));
  NOR2X1 G2036 (.A1(I190), .A2(I191), .ZN(W95));
  NOR2X1 G2037 (.A1(I192), .A2(I193), .ZN(W96));
  NOR2X1 G2038 (.A1(I604), .A2(I788), .ZN(W965));
  NOR2X1 G2039 (.A1(I956), .A2(W135), .ZN(W963));
  NOR2X1 G2040 (.A1(W939), .A2(I175), .ZN(W1039));
  NOR2X1 G2041 (.A1(W334), .A2(W180), .ZN(W1040));
  NOR2X1 G2042 (.A1(I252), .A2(I253), .ZN(W126));
  NOR2X1 G2043 (.A1(I661), .A2(I996), .ZN(O81));
  NOR2X1 G2044 (.A1(I231), .A2(W527), .ZN(W1041));
  NOR2X1 G2045 (.A1(W31), .A2(I873), .ZN(W960));
  NOR2X1 G2046 (.A1(W505), .A2(W411), .ZN(W1042));
  NOR2X1 G2047 (.A1(W377), .A2(I418), .ZN(W959));
  NOR2X1 G2048 (.A1(I216), .A2(I217), .ZN(W108));
  NOR2X1 G2049 (.A1(I176), .A2(W1028), .ZN(W1573));
  NOR2X1 G2050 (.A1(I218), .A2(I219), .ZN(W109));
  NOR2X1 G2051 (.A1(I729), .A2(W230), .ZN(W1537));
  NOR2X1 G2052 (.A1(W46), .A2(W1084), .ZN(O80));
  NOR2X1 G2053 (.A1(W593), .A2(W197), .ZN(W937));
  NOR2X1 G2054 (.A1(W154), .A2(W605), .ZN(W935));
  NOR2X1 G2055 (.A1(W1335), .A2(I446), .ZN(W1543));
  NOR2X1 G2056 (.A1(W724), .A2(I786), .ZN(W933));
  NOR2X1 G2057 (.A1(W935), .A2(I405), .ZN(W1063));
  NOR2X1 G2058 (.A1(I514), .A2(W395), .ZN(W932));
  NOR2X1 G2059 (.A1(I316), .A2(I317), .ZN(W158));
  NOR2X1 G2060 (.A1(W359), .A2(I5), .ZN(W925));
  NOR2X1 G2061 (.A1(W533), .A2(I216), .ZN(W1549));
  NOR2X1 G2062 (.A1(W45), .A2(W74), .ZN(W1536));
  NOR2X1 G2063 (.A1(W683), .A2(I27), .ZN(W922));
  NOR2X1 G2064 (.A1(I964), .A2(W383), .ZN(W921));
  NOR2X1 G2065 (.A1(I330), .A2(I331), .ZN(W165));
  NOR2X1 G2066 (.A1(I597), .A2(W597), .ZN(W1535));
  NOR2X1 G2067 (.A1(I334), .A2(I335), .ZN(W167));
  NOR2X1 G2068 (.A1(I336), .A2(I337), .ZN(W168));
  NOR2X1 G2069 (.A1(I338), .A2(I339), .ZN(W169));
  NOR2X1 G2070 (.A1(W589), .A2(I948), .ZN(W945));
  NOR2X1 G2071 (.A1(W966), .A2(I639), .ZN(W1052));
  NOR2X1 G2072 (.A1(I256), .A2(I257), .ZN(W128));
  NOR2X1 G2073 (.A1(W1185), .A2(I670), .ZN(W1558));
  NOR2X1 G2074 (.A1(W641), .A2(W494), .ZN(W1055));
  NOR2X1 G2075 (.A1(I260), .A2(I261), .ZN(W130));
  NOR2X1 G2076 (.A1(W33), .A2(W998), .ZN(W1556));
  NOR2X1 G2077 (.A1(I85), .A2(I574), .ZN(W947));
  NOR2X1 G2078 (.A1(I262), .A2(I263), .ZN(W131));
  NOR2X1 G2079 (.A1(W1181), .A2(W1271), .ZN(W1555));
  NOR2X1 G2080 (.A1(I174), .A2(I175), .ZN(W87));
  NOR2X1 G2081 (.A1(W279), .A2(I277), .ZN(W1057));
  NOR2X1 G2082 (.A1(W661), .A2(W63), .ZN(W1058));
  NOR2X1 G2083 (.A1(W520), .A2(I864), .ZN(W943));
  NOR2X1 G2084 (.A1(I266), .A2(I267), .ZN(W133));
  NOR2X1 G2085 (.A1(W758), .A2(W1062), .ZN(W1551));
  NOR2X1 G2086 (.A1(I270), .A2(I271), .ZN(W135));
  NOR2X1 G2087 (.A1(I5), .A2(W460), .ZN(W1059));
  NOR2X1 G2088 (.A1(I282), .A2(I283), .ZN(W141));
  NOR2X1 G2089 (.A1(I64), .A2(I65), .ZN(W32));
  NOR2X1 G2090 (.A1(I881), .A2(W252), .ZN(W1000));
  NOR2X1 G2091 (.A1(W261), .A2(W565), .ZN(W998));
  NOR2X1 G2092 (.A1(I48), .A2(I49), .ZN(W24));
  NOR2X1 G2093 (.A1(I50), .A2(I51), .ZN(W25));
  NOR2X1 G2094 (.A1(W735), .A2(W678), .ZN(W991));
  NOR2X1 G2095 (.A1(I56), .A2(I57), .ZN(W28));
  NOR2X1 G2096 (.A1(I366), .A2(I208), .ZN(W1621));
  NOR2X1 G2097 (.A1(W1226), .A2(W713), .ZN(W1620));
  NOR2X1 G2098 (.A1(W764), .A2(W1589), .ZN(W1617));
  NOR2X1 G2099 (.A1(W698), .A2(W785), .ZN(W1017));
  NOR2X1 G2100 (.A1(I8), .A2(I657), .ZN(W1615));
  NOR2X1 G2101 (.A1(W619), .A2(W917), .ZN(W988));
  NOR2X1 G2102 (.A1(I70), .A2(I71), .ZN(W35));
  NOR2X1 G2103 (.A1(W192), .A2(W678), .ZN(W1021));
  NOR2X1 G2104 (.A1(I74), .A2(I75), .ZN(W37));
  NOR2X1 G2105 (.A1(W944), .A2(W116), .ZN(W1611));
  NOR2X1 G2106 (.A1(W851), .A2(I566), .ZN(W1610));
  NOR2X1 G2107 (.A1(W866), .A2(I302), .ZN(W985));
  NOR2X1 G2108 (.A1(I78), .A2(I79), .ZN(W39));
  NOR2X1 G2109 (.A1(I26), .A2(I27), .ZN(W13));
  NOR2X1 G2110 (.A1(W1202), .A2(I180), .ZN(W1638));
  NOR2X1 G2111 (.A1(I6), .A2(I7), .ZN(W3));
  NOR2X1 G2112 (.A1(I543), .A2(I681), .ZN(W1634));
  NOR2X1 G2113 (.A1(I8), .A2(I9), .ZN(W4));
  NOR2X1 G2114 (.A1(I10), .A2(I11), .ZN(W5));
  NOR2X1 G2115 (.A1(I396), .A2(W550), .ZN(O88));
  NOR2X1 G2116 (.A1(I806), .A2(W127), .ZN(W1005));
  NOR2X1 G2117 (.A1(I20), .A2(I21), .ZN(W10));
  NOR2X1 G2118 (.A1(W37), .A2(W1441), .ZN(W1630));
  NOR2X1 G2119 (.A1(I80), .A2(I81), .ZN(W40));
  NOR2X1 G2120 (.A1(W915), .A2(W474), .ZN(W1629));
  NOR2X1 G2121 (.A1(W1464), .A2(W1455), .ZN(W1628));
  NOR2X1 G2122 (.A1(I30), .A2(I31), .ZN(W15));
  NOR2X1 G2123 (.A1(I714), .A2(W804), .ZN(W1014));
  NOR2X1 G2124 (.A1(I200), .A2(I970), .ZN(W1627));
  NOR2X1 G2125 (.A1(W579), .A2(I455), .ZN(W1015));
  NOR2X1 G2126 (.A1(I42), .A2(I43), .ZN(W21));
  NOR2X1 G2127 (.A1(W51), .A2(W1190), .ZN(W1625));
  NOR2X1 G2128 (.A1(W337), .A2(I560), .ZN(W968));
  NOR2X1 G2129 (.A1(W912), .A2(I958), .ZN(W976));
  NOR2X1 G2130 (.A1(W17), .A2(I242), .ZN(W1589));
  NOR2X1 G2131 (.A1(W118), .A2(I370), .ZN(W1588));
  NOR2X1 G2132 (.A1(I146), .A2(I147), .ZN(W73));
  NOR2X1 G2133 (.A1(I474), .A2(I547), .ZN(W969));
  NOR2X1 G2134 (.A1(I844), .A2(W127), .ZN(W1586));
  NOR2X1 G2135 (.A1(W764), .A2(W1231), .ZN(W1585));
  NOR2X1 G2136 (.A1(I150), .A2(I151), .ZN(W75));
  NOR2X1 G2137 (.A1(W700), .A2(W826), .ZN(W1583));
  NOR2X1 G2138 (.A1(I157), .A2(I27), .ZN(W1592));
  NOR2X1 G2139 (.A1(I152), .A2(I153), .ZN(W76));
  NOR2X1 G2140 (.A1(I570), .A2(I304), .ZN(W967));
  NOR2X1 G2141 (.A1(I160), .A2(I161), .ZN(W80));
  NOR2X1 G2142 (.A1(I162), .A2(I163), .ZN(W81));
  NOR2X1 G2143 (.A1(I907), .A2(I581), .ZN(W1035));
  NOR2X1 G2144 (.A1(I168), .A2(I169), .ZN(W84));
  NOR2X1 G2145 (.A1(I170), .A2(I171), .ZN(O1));
  NOR2X1 G2146 (.A1(W182), .A2(W1145), .ZN(W1582));
  NOR2X1 G2147 (.A1(W681), .A2(W766), .ZN(W979));
  NOR2X1 G2148 (.A1(W1268), .A2(W149), .ZN(O85));
  NOR2X1 G2149 (.A1(W872), .A2(I981), .ZN(W1023));
  NOR2X1 G2150 (.A1(W687), .A2(W294), .ZN(W1024));
  NOR2X1 G2151 (.A1(W922), .A2(W1246), .ZN(W1607));
  NOR2X1 G2152 (.A1(I219), .A2(I111), .ZN(O84));
  NOR2X1 G2153 (.A1(I90), .A2(I91), .ZN(W45));
  NOR2X1 G2154 (.A1(I110), .A2(I111), .ZN(W55));
  NOR2X1 G2155 (.A1(I112), .A2(I113), .ZN(W56));
  NOR2X1 G2156 (.A1(I114), .A2(I115), .ZN(W57));
  NOR2X1 G2157 (.A1(W32), .A2(W1250), .ZN(W1572));
  NOR2X1 G2158 (.A1(W747), .A2(W37), .ZN(W1027));
  NOR2X1 G2159 (.A1(I612), .A2(W585), .ZN(W1028));
  NOR2X1 G2160 (.A1(I337), .A2(W375), .ZN(W1600));
  NOR2X1 G2161 (.A1(I464), .A2(I546), .ZN(W1599));
  NOR2X1 G2162 (.A1(I120), .A2(I121), .ZN(W60));
  NOR2X1 G2163 (.A1(I122), .A2(I123), .ZN(W61));
  NOR2X1 G2164 (.A1(I137), .A2(W1280), .ZN(W1596));
  NOR2X1 G2165 (.A1(I819), .A2(W917), .ZN(W977));
  NOR2X1 G2166 (.A1(W797), .A2(W734), .ZN(W1075));
  NOR2X1 G2167 (.A1(I72), .A2(W1054), .ZN(W1078));
  NOR2X1 G2168 (.A1(W182), .A2(W114), .ZN(W894));
  NOR2X1 G2169 (.A1(I400), .A2(I401), .ZN(W200));
  NOR2X1 G2170 (.A1(I102), .A2(W151), .ZN(W892));
  NOR2X1 G2171 (.A1(W597), .A2(W80), .ZN(W1091));
  NOR2X1 G2172 (.A1(I406), .A2(I407), .ZN(W203));
  NOR2X1 G2173 (.A1(I975), .A2(W539), .ZN(W1508));
  NOR2X1 G2174 (.A1(I203), .A2(I303), .ZN(W1076));
  NOR2X1 G2175 (.A1(W8), .A2(W418), .ZN(W1511));
  NOR2X1 G2176 (.A1(I332), .A2(W489), .ZN(O76));
  NOR2X1 G2177 (.A1(W599), .A2(I509), .ZN(W888));
  NOR2X1 G2178 (.A1(I218), .A2(W806), .ZN(W1531));
  NOR2X1 G2179 (.A1(I225), .A2(W864), .ZN(W918));
  NOR2X1 G2180 (.A1(I412), .A2(I413), .ZN(W206));
  NOR2X1 G2181 (.A1(I414), .A2(I415), .ZN(W207));
  NOR2X1 G2182 (.A1(I625), .A2(I674), .ZN(W1092));
  NOR2X1 G2183 (.A1(W1040), .A2(W969), .ZN(W1094));
  NOR2X1 G2184 (.A1(W358), .A2(I972), .ZN(W1525));
  NOR2X1 G2185 (.A1(W626), .A2(I240), .ZN(W1089));
  NOR2X1 G2186 (.A1(W1358), .A2(I440), .ZN(W1513));
  NOR2X1 G2187 (.A1(I364), .A2(I365), .ZN(W182));
  NOR2X1 G2188 (.A1(W554), .A2(W521), .ZN(W1514));
  NOR2X1 G2189 (.A1(I245), .A2(I354), .ZN(W896));
  NOR2X1 G2190 (.A1(I384), .A2(I385), .ZN(W192));
  NOR2X1 G2191 (.A1(I121), .A2(W325), .ZN(W906));
  NOR2X1 G2192 (.A1(W566), .A2(W451), .ZN(W1086));
  NOR2X1 G2193 (.A1(I46), .A2(W1133), .ZN(W1516));
  NOR2X1 G2194 (.A1(I374), .A2(I375), .ZN(W187));
  NOR2X1 G2195 (.A1(I96), .A2(W289), .ZN(W1084));
  NOR2X1 G2196 (.A1(I598), .A2(I284), .ZN(W1085));
  NOR2X1 G2197 (.A1(I943), .A2(W728), .ZN(W902));
  NOR2X1 G2198 (.A1(I414), .A2(I208), .ZN(W1518));
  NOR2X1 G2199 (.A1(I860), .A2(W364), .ZN(W920));
  NOR2X1 G2200 (.A1(W901), .A2(W322), .ZN(W919));
  NOR2X1 G2201 (.A1(I176), .A2(I182), .ZN(W887));
  NOR2X1 G2202 (.A1(I346), .A2(I347), .ZN(W173));
  NOR2X1 G2203 (.A1(W130), .A2(W1465), .ZN(O78));
  NOR2X1 G2204 (.A1(W875), .A2(I294), .ZN(W1072));
  NANDX1 G2205 (.A1(W1070), .A2(W2358), .ZN(O929));
  NANDX1 G2206 (.A1(I488), .A2(W366), .ZN(W693));
  NANDX1 G2207 (.A1(W1357), .A2(W1368), .ZN(W3616));
  NANDX1 G2208 (.A1(W1542), .A2(W790), .ZN(O928));
  NANDX1 G2209 (.A1(I288), .A2(W1343), .ZN(O677));
  NANDX1 G2210 (.A1(W615), .A2(I352), .ZN(W898));
  NANDX1 G2211 (.A1(I285), .A2(I640), .ZN(W694));
  NANDX1 G2212 (.A1(W2442), .A2(W395), .ZN(W3983));
  NANDX1 G2213 (.A1(W2408), .A2(W2255), .ZN(W3614));
  NANDX1 G2214 (.A1(W2562), .A2(W2533), .ZN(W4528));
  NANDX1 G2215 (.A1(W281), .A2(W1402), .ZN(O523));
  NANDX1 G2216 (.A1(W3917), .A2(I112), .ZN(O676));
  NANDX1 G2217 (.A1(I54), .A2(I974), .ZN(W978));
  NANDX1 G2218 (.A1(W1851), .A2(W1775), .ZN(W4534));
  NANDX1 G2219 (.A1(W2889), .A2(W2638), .ZN(W4502));
  NANDX1 G2220 (.A1(W2087), .A2(W3005), .ZN(W4485));
  NANDX1 G2221 (.A1(W411), .A2(W238), .ZN(W972));
  NANDX1 G2222 (.A1(I546), .A2(I374), .ZN(W702));
  NANDX1 G2223 (.A1(W1302), .A2(W1962), .ZN(W3629));
  NANDX1 G2224 (.A1(W261), .A2(I198), .ZN(W973));
  NANDX1 G2225 (.A1(W483), .A2(I120), .ZN(W3625));
  NANDX1 G2226 (.A1(W3827), .A2(W2278), .ZN(W4495));
  NANDX1 G2227 (.A1(W639), .A2(W1814), .ZN(W4498));
  NANDX1 G2228 (.A1(W4134), .A2(W2012), .ZN(O937));
  NANDX1 G2229 (.A1(W2296), .A2(I518), .ZN(W4504));
  NANDX1 G2230 (.A1(W1297), .A2(W3500), .ZN(W4508));
  NANDX1 G2231 (.A1(I79), .A2(I939), .ZN(W975));
  NANDX1 G2232 (.A1(W3946), .A2(W1800), .ZN(O924));
  NANDX1 G2233 (.A1(W545), .A2(W3306), .ZN(O626));
  NANDX1 G2234 (.A1(W1696), .A2(W3750), .ZN(O1048));
  NANDX1 G2235 (.A1(W1805), .A2(W1802), .ZN(O527));
  NANDX1 G2236 (.A1(W3385), .A2(W2713), .ZN(W3618));
  NANDX1 G2237 (.A1(I702), .A2(I623), .ZN(W683));
  NANDX1 G2238 (.A1(W242), .A2(W505), .ZN(W983));
  NANDX1 G2239 (.A1(W209), .A2(W380), .ZN(W982));
  NANDX1 G2240 (.A1(W86), .A2(W601), .ZN(O519));
  NANDX1 G2241 (.A1(W1449), .A2(W1816), .ZN(O633));
  NANDX1 G2242 (.A1(W623), .A2(W308), .ZN(W679));
  NANDX1 G2243 (.A1(W3352), .A2(W515), .ZN(W4554));
  NANDX1 G2244 (.A1(W1817), .A2(W3370), .ZN(W3601));
  NANDX1 G2245 (.A1(W4080), .A2(W349), .ZN(W4553));
  NANDX1 G2246 (.A1(W2872), .A2(W3713), .ZN(O946));
  NANDX1 G2247 (.A1(W2336), .A2(W3329), .ZN(W3603));
  NANDX1 G2248 (.A1(W3256), .A2(I777), .ZN(O520));
  NANDX1 G2249 (.A1(W120), .A2(I323), .ZN(W682));
  NANDX1 G2250 (.A1(W2294), .A2(W2564), .ZN(W4740));
  NANDX1 G2251 (.A1(W96), .A2(W4421), .ZN(W4547));
  NANDX1 G2252 (.A1(W3223), .A2(W3314), .ZN(W3608));
  NANDX1 G2253 (.A1(I272), .A2(I871), .ZN(W687));
  NANDX1 G2254 (.A1(W1144), .A2(W1398), .ZN(W3884));
  NANDX1 G2255 (.A1(I543), .A2(I587), .ZN(O941));
  NANDX1 G2256 (.A1(W3646), .A2(W812), .ZN(W3879));
  NANDX1 G2257 (.A1(W2009), .A2(W2178), .ZN(O940));
  NANDX1 G2258 (.A1(W29), .A2(I730), .ZN(W618));
  NANDX1 G2259 (.A1(I284), .A2(I713), .ZN(O630));
  NANDX1 G2260 (.A1(W432), .A2(W582), .ZN(W859));
  NANDX1 G2261 (.A1(I895), .A2(I104), .ZN(W3875));
  NANDX1 G2262 (.A1(W1283), .A2(W787), .ZN(O521));
  NANDX1 G2263 (.A1(W3121), .A2(W1341), .ZN(O675));
  NANDX1 G2264 (.A1(W3442), .A2(I350), .ZN(O938));
  NANDX1 G2265 (.A1(W4270), .A2(W772), .ZN(O908));
  NANDX1 G2266 (.A1(W157), .A2(W145), .ZN(W685));
  NANDX1 G2267 (.A1(W496), .A2(W41), .ZN(W686));
  NANDX1 G2268 (.A1(W1630), .A2(W211), .ZN(W3641));
  NANDX1 G2269 (.A1(W1168), .A2(W14), .ZN(O857));
  NANDX1 G2270 (.A1(W4584), .A2(W4012), .ZN(W4747));
  NANDX1 G2271 (.A1(W1383), .A2(W2402), .ZN(W4430));
  NANDX1 G2272 (.A1(W579), .A2(I511), .ZN(W719));
  NANDX1 G2273 (.A1(W631), .A2(W1536), .ZN(W3644));
  NANDX1 G2274 (.A1(W356), .A2(W2077), .ZN(O880));
  NANDX1 G2275 (.A1(W793), .A2(W817), .ZN(O34));
  NANDX1 G2276 (.A1(I840), .A2(I17), .ZN(W4437));
  NANDX1 G2277 (.A1(W2924), .A2(W2455), .ZN(W4009));
  NANDX1 G2278 (.A1(W1053), .A2(I550), .ZN(W1639));
  NANDX1 G2279 (.A1(W1794), .A2(W1930), .ZN(W4438));
  NANDX1 G2280 (.A1(W4190), .A2(W622), .ZN(W4439));
  NANDX1 G2281 (.A1(I929), .A2(W65), .ZN(W717));
  NANDX1 G2282 (.A1(W804), .A2(I728), .ZN(W849));
  NANDX1 G2283 (.A1(I14), .A2(W651), .ZN(W899));
  NANDX1 G2284 (.A1(W3522), .A2(W1789), .ZN(O883));
  NANDX1 G2285 (.A1(W262), .A2(W2719), .ZN(W4016));
  NANDX1 G2286 (.A1(W475), .A2(W892), .ZN(W4416));
  NANDX1 G2287 (.A1(W709), .A2(I964), .ZN(W724));
  NANDX1 G2288 (.A1(W1087), .A2(W3616), .ZN(W3652));
  NANDX1 G2289 (.A1(I240), .A2(W2448), .ZN(O870));
  NANDX1 G2290 (.A1(W1692), .A2(W2714), .ZN(W4421));
  NANDX1 G2291 (.A1(I758), .A2(W340), .ZN(W722));
  NANDX1 G2292 (.A1(W263), .A2(I537), .ZN(W903));
  NANDX1 G2293 (.A1(I198), .A2(I587), .ZN(W966));
  NANDX1 G2294 (.A1(W1594), .A2(W4010), .ZN(O884));
  NANDX1 G2295 (.A1(I81), .A2(I868), .ZN(W848));
  NANDX1 G2296 (.A1(I533), .A2(W760), .ZN(W4010));
  NANDX1 G2297 (.A1(I686), .A2(W2824), .ZN(O540));
  NANDX1 G2298 (.A1(W2081), .A2(W1814), .ZN(W3648));
  NANDX1 G2299 (.A1(W135), .A2(W3093), .ZN(O872));
  NANDX1 G2300 (.A1(W2576), .A2(I288), .ZN(O538));
  NANDX1 G2301 (.A1(W276), .A2(I179), .ZN(W4429));
  NANDX1 G2302 (.A1(W4190), .A2(W1861), .ZN(W4468));
  NANDX1 G2303 (.A1(W1966), .A2(W96), .ZN(W4743));
  NANDX1 G2304 (.A1(W3223), .A2(W1516), .ZN(O896));
  NANDX1 G2305 (.A1(W1039), .A2(W1534), .ZN(W4463));
  NANDX1 G2306 (.A1(W3419), .A2(W3942), .ZN(O897));
  NANDX1 G2307 (.A1(W57), .A2(I958), .ZN(W855));
  NANDX1 G2308 (.A1(W940), .A2(W722), .ZN(W970));
  NANDX1 G2309 (.A1(W1207), .A2(W124), .ZN(W3634));
  NANDX1 G2310 (.A1(W1977), .A2(W163), .ZN(O898));
  NANDX1 G2311 (.A1(W685), .A2(W268), .ZN(W711));
  NANDX1 G2312 (.A1(I491), .A2(I191), .ZN(W707));
  NANDX1 G2313 (.A1(W351), .A2(W1738), .ZN(O904));
  NANDX1 G2314 (.A1(I965), .A2(W539), .ZN(O906));
  NANDX1 G2315 (.A1(W3563), .A2(I755), .ZN(W3866));
  NANDX1 G2316 (.A1(I658), .A2(W1156), .ZN(W3867));
  NANDX1 G2317 (.A1(W2722), .A2(I907), .ZN(O907));
  NANDX1 G2318 (.A1(W4392), .A2(W1599), .ZN(W4564));
  NANDX1 G2319 (.A1(W3140), .A2(W3336), .ZN(O911));
  NANDX1 G2320 (.A1(W1194), .A2(W1569), .ZN(W4458));
  NANDX1 G2321 (.A1(I393), .A2(I352), .ZN(W854));
  NANDX1 G2322 (.A1(W1021), .A2(I424), .ZN(W3638));
  NANDX1 G2323 (.A1(I721), .A2(I563), .ZN(W712));
  NANDX1 G2324 (.A1(W3429), .A2(W1035), .ZN(O891));
  NANDX1 G2325 (.A1(I634), .A2(I285), .ZN(W713));
  NANDX1 G2326 (.A1(I756), .A2(W296), .ZN(W714));
  NANDX1 G2327 (.A1(W2395), .A2(W3060), .ZN(W3992));
  NANDX1 G2328 (.A1(W668), .A2(I165), .ZN(W4450));
  NANDX1 G2329 (.A1(W15), .A2(I794), .ZN(W1008));
  NANDX1 G2330 (.A1(W4236), .A2(W1990), .ZN(O886));
  NANDX1 G2331 (.A1(W4362), .A2(W2956), .ZN(W4446));
  NANDX1 G2332 (.A1(I864), .A2(I682), .ZN(W4003));
  NANDX1 G2333 (.A1(W139), .A2(W1366), .ZN(W3510));
  NANDX1 G2334 (.A1(W874), .A2(W2773), .ZN(O885));
  NANDX1 G2335 (.A1(I401), .A2(W3386), .ZN(O652));
  NANDX1 G2336 (.A1(I100), .A2(W1913), .ZN(O994));
  NANDX1 G2337 (.A1(I382), .A2(W265), .ZN(W1001));
  NANDX1 G2338 (.A1(W286), .A2(I233), .ZN(W874));
  NANDX1 G2339 (.A1(W3509), .A2(W2771), .ZN(W3541));
  NANDX1 G2340 (.A1(W4104), .A2(W3638), .ZN(O995));
  NANDX1 G2341 (.A1(W2854), .A2(W2304), .ZN(O654));
  NANDX1 G2342 (.A1(I530), .A2(W235), .ZN(W877));
  NANDX1 G2343 (.A1(W2285), .A2(W3473), .ZN(W4661));
  NANDX1 G2344 (.A1(W981), .A2(W3395), .ZN(W3905));
  NANDX1 G2345 (.A1(I960), .A2(I80), .ZN(W627));
  NANDX1 G2346 (.A1(W3757), .A2(W4640), .ZN(W4662));
  NANDX1 G2347 (.A1(W2507), .A2(I240), .ZN(W4663));
  NANDX1 G2348 (.A1(W416), .A2(I257), .ZN(W3540));
  NANDX1 G2349 (.A1(I625), .A2(W4439), .ZN(O996));
  NANDX1 G2350 (.A1(W3880), .A2(W3710), .ZN(O1030));
  NANDX1 G2351 (.A1(W3362), .A2(W1674), .ZN(O499));
  NANDX1 G2352 (.A1(W497), .A2(I274), .ZN(O998));
  NANDX1 G2353 (.A1(W855), .A2(I580), .ZN(W891));
  NANDX1 G2354 (.A1(I23), .A2(W2699), .ZN(O658));
  NANDX1 G2355 (.A1(W1584), .A2(I941), .ZN(W4651));
  NANDX1 G2356 (.A1(W3286), .A2(I829), .ZN(O659));
  NANDX1 G2357 (.A1(W1587), .A2(W930), .ZN(W3900));
  NANDX1 G2358 (.A1(W723), .A2(W2128), .ZN(W4724));
  NANDX1 G2359 (.A1(I493), .A2(I666), .ZN(W648));
  NANDX1 G2360 (.A1(W1701), .A2(W10), .ZN(W3547));
  NANDX1 G2361 (.A1(W606), .A2(I817), .ZN(W997));
  NANDX1 G2362 (.A1(I875), .A2(I134), .ZN(W3552));
  NANDX1 G2363 (.A1(I534), .A2(I499), .ZN(W995));
  NANDX1 G2364 (.A1(W3428), .A2(W3407), .ZN(O660));
  NANDX1 G2365 (.A1(I777), .A2(W537), .ZN(W873));
  NANDX1 G2366 (.A1(W668), .A2(W2193), .ZN(W4642));
  NANDX1 G2367 (.A1(W2607), .A2(W521), .ZN(O503));
  NANDX1 G2368 (.A1(W2548), .A2(W3954), .ZN(W4700));
  NANDX1 G2369 (.A1(W4249), .A2(W2338), .ZN(O1014));
  NANDX1 G2370 (.A1(W476), .A2(W3217), .ZN(W3527));
  NANDX1 G2371 (.A1(W2065), .A2(I562), .ZN(W3927));
  NANDX1 G2372 (.A1(W1063), .A2(I188), .ZN(W4694));
  NANDX1 G2373 (.A1(W1367), .A2(I902), .ZN(O1025));
  NANDX1 G2374 (.A1(W833), .A2(W722), .ZN(W1006));
  NANDX1 G2375 (.A1(W81), .A2(W773), .ZN(O1016));
  NANDX1 G2376 (.A1(W1048), .A2(W3425), .ZN(O1017));
  NANDX1 G2377 (.A1(W1764), .A2(W4499), .ZN(W4690));
  NANDX1 G2378 (.A1(W2422), .A2(I198), .ZN(W4702));
  NANDX1 G2379 (.A1(W2913), .A2(W3244), .ZN(O495));
  NANDX1 G2380 (.A1(W71), .A2(W2443), .ZN(W3518));
  NANDX1 G2381 (.A1(W1360), .A2(W3381), .ZN(W3517));
  NANDX1 G2382 (.A1(W675), .A2(I894), .ZN(O1021));
  NANDX1 G2383 (.A1(I246), .A2(I182), .ZN(O493));
  NANDX1 G2384 (.A1(W160), .A2(I457), .ZN(W629));
  NANDX1 G2385 (.A1(W454), .A2(W1206), .ZN(O505));
  NANDX1 G2386 (.A1(I909), .A2(I357), .ZN(W635));
  NANDX1 G2387 (.A1(W994), .A2(W1942), .ZN(O1008));
  NANDX1 G2388 (.A1(W2340), .A2(W504), .ZN(O1006));
  NANDX1 G2389 (.A1(I885), .A2(W2940), .ZN(W3529));
  NANDX1 G2390 (.A1(W2610), .A2(W1543), .ZN(O497));
  NANDX1 G2391 (.A1(W386), .A2(I184), .ZN(W640));
  NANDX1 G2392 (.A1(W2520), .A2(W2223), .ZN(W3909));
  NANDX1 G2393 (.A1(I633), .A2(W4007), .ZN(W4671));
  NANDX1 G2394 (.A1(I778), .A2(W1045), .ZN(O1000));
  NANDX1 G2395 (.A1(W684), .A2(W740), .ZN(W880));
  NANDX1 G2396 (.A1(W4169), .A2(W3977), .ZN(O1027));
  NANDX1 G2397 (.A1(W1526), .A2(W4480), .ZN(O999));
  NANDX1 G2398 (.A1(W1758), .A2(W651), .ZN(W4715));
  NANDX1 G2399 (.A1(W1315), .A2(W2874), .ZN(W3535));
  NANDX1 G2400 (.A1(W3653), .A2(W1663), .ZN(W4667));
  NANDX1 G2401 (.A1(I815), .A2(W531), .ZN(O966));
  NANDX1 G2402 (.A1(I138), .A2(I478), .ZN(W621));
  NANDX1 G2403 (.A1(I706), .A2(W2802), .ZN(O670));
  NANDX1 G2404 (.A1(I870), .A2(I838), .ZN(W671));
  NANDX1 G2405 (.A1(I989), .A2(W3054), .ZN(O1042));
  NANDX1 G2406 (.A1(W1837), .A2(W325), .ZN(O1040));
  NANDX1 G2407 (.A1(W1133), .A2(W3141), .ZN(W3896));
  NANDX1 G2408 (.A1(W53), .A2(W1193), .ZN(W4590));
  NANDX1 G2409 (.A1(W133), .A2(I732), .ZN(O964));
  NANDX1 G2410 (.A1(W2888), .A2(W1067), .ZN(W3590));
  NANDX1 G2411 (.A1(W1498), .A2(W2720), .ZN(W4600));
  NANDX1 G2412 (.A1(W3798), .A2(I991), .ZN(O969));
  NANDX1 G2413 (.A1(W1525), .A2(I172), .ZN(W3588));
  NANDX1 G2414 (.A1(I991), .A2(W2509), .ZN(W3587));
  NANDX1 G2415 (.A1(W1543), .A2(W210), .ZN(O511));
  NANDX1 G2416 (.A1(W1427), .A2(W45), .ZN(W3957));
  NANDX1 G2417 (.A1(W987), .A2(W2138), .ZN(O665));
  NANDX1 G2418 (.A1(I386), .A2(I108), .ZN(W989));
  NANDX1 G2419 (.A1(I534), .A2(W4084), .ZN(W4581));
  NANDX1 G2420 (.A1(W1091), .A2(W1040), .ZN(O634));
  NANDX1 G2421 (.A1(I209), .A2(W530), .ZN(W984));
  NANDX1 G2422 (.A1(W2775), .A2(W427), .ZN(W3512));
  NANDX1 G2423 (.A1(W2516), .A2(W3510), .ZN(O1044));
  NANDX1 G2424 (.A1(W87), .A2(I980), .ZN(W674));
  NANDX1 G2425 (.A1(I598), .A2(W166), .ZN(O960));
  NANDX1 G2426 (.A1(W2803), .A2(W3157), .ZN(W3970));
  NANDX1 G2427 (.A1(W3358), .A2(W3985), .ZN(W4574));
  NANDX1 G2428 (.A1(W1303), .A2(W2992), .ZN(O957));
  NANDX1 G2429 (.A1(W323), .A2(W339), .ZN(W619));
  NANDX1 G2430 (.A1(I409), .A2(I730), .ZN(W4572));
  NANDX1 G2431 (.A1(W348), .A2(I957), .ZN(O32));
  NANDX1 G2432 (.A1(I352), .A2(I982), .ZN(W628));
  NANDX1 G2433 (.A1(W845), .A2(W2886), .ZN(O951));
  NANDX1 G2434 (.A1(W124), .A2(W284), .ZN(W656));
  NANDX1 G2435 (.A1(W701), .A2(I405), .ZN(W994));
  NANDX1 G2436 (.A1(I885), .A2(W689), .ZN(W3563));
  NANDX1 G2437 (.A1(W2773), .A2(W727), .ZN(O984));
  NANDX1 G2438 (.A1(I607), .A2(W2901), .ZN(W4635));
  NANDX1 G2439 (.A1(I8), .A2(I285), .ZN(W654));
  NANDX1 G2440 (.A1(W2484), .A2(W876), .ZN(W4633));
  NANDX1 G2441 (.A1(W2063), .A2(W2386), .ZN(W3568));
  NANDX1 G2442 (.A1(W689), .A2(W242), .ZN(W3570));
  NANDX1 G2443 (.A1(W2619), .A2(W1047), .ZN(W4632));
  NANDX1 G2444 (.A1(W2272), .A2(I768), .ZN(W4631));
  NANDX1 G2445 (.A1(I635), .A2(W81), .ZN(W625));
  NANDX1 G2446 (.A1(I711), .A2(W3527), .ZN(W3571));
  NANDX1 G2447 (.A1(I176), .A2(W1840), .ZN(W3899));
  NANDX1 G2448 (.A1(W297), .A2(W3974), .ZN(W4629));
  NANDX1 G2449 (.A1(W844), .A2(W150), .ZN(W881));
  NANDX1 G2450 (.A1(W3438), .A2(W1506), .ZN(W3977));
  NANDX1 G2451 (.A1(W850), .A2(I43), .ZN(W872));
  NANDX1 G2452 (.A1(W2797), .A2(W2451), .ZN(O661));
  NANDX1 G2453 (.A1(I686), .A2(I950), .ZN(W658));
  NANDX1 G2454 (.A1(W206), .A2(I303), .ZN(W659));
  NANDX1 G2455 (.A1(W1586), .A2(W2586), .ZN(W4621));
  NANDX1 G2456 (.A1(I866), .A2(I355), .ZN(O977));
  NANDX1 G2457 (.A1(W4504), .A2(W57), .ZN(O973));
  NANDX1 G2458 (.A1(W552), .A2(W586), .ZN(O33));
  NANDX1 G2459 (.A1(W2647), .A2(W301), .ZN(W3576));
  NANDX1 G2460 (.A1(W663), .A2(I280), .ZN(W990));
  NANDX1 G2461 (.A1(W1748), .A2(W2259), .ZN(W3578));
  NANDX1 G2462 (.A1(W1636), .A2(W3267), .ZN(O509));
  NANDX1 G2463 (.A1(W3180), .A2(W3901), .ZN(O971));
  NANDX1 G2464 (.A1(W123), .A2(W3699), .ZN(W3954));
  NANDX1 G2465 (.A1(W1479), .A2(W1412), .ZN(O645));
  NANDX1 G2466 (.A1(I106), .A2(W700), .ZN(O569));
  NANDX1 G2467 (.A1(W402), .A2(W195), .ZN(W4184));
  NANDX1 G2468 (.A1(I987), .A2(I659), .ZN(O769));
  NANDX1 G2469 (.A1(I982), .A2(W781), .ZN(O570));
  NANDX1 G2470 (.A1(W416), .A2(W710), .ZN(W915));
  NANDX1 G2471 (.A1(W1982), .A2(W1613), .ZN(W4191));
  NANDX1 G2472 (.A1(W2476), .A2(W3400), .ZN(W3829));
  NANDX1 G2473 (.A1(W3447), .A2(W3288), .ZN(O771));
  NANDX1 G2474 (.A1(W654), .A2(W199), .ZN(W824));
  NANDX1 G2475 (.A1(W2017), .A2(I660), .ZN(W4183));
  NANDX1 G2476 (.A1(I486), .A2(W888), .ZN(O776));
  NANDX1 G2477 (.A1(W258), .A2(W403), .ZN(W3737));
  NANDX1 G2478 (.A1(W2619), .A2(W236), .ZN(O777));
  NANDX1 G2479 (.A1(W3606), .A2(W1789), .ZN(O778));
  NANDX1 G2480 (.A1(W3415), .A2(I100), .ZN(O779));
  NANDX1 G2481 (.A1(I117), .A2(I476), .ZN(W942));
  NANDX1 G2482 (.A1(I145), .A2(W493), .ZN(O36));
  NANDX1 G2483 (.A1(W1827), .A2(W1594), .ZN(W4080));
  NANDX1 G2484 (.A1(W627), .A2(W3379), .ZN(O573));
  NANDX1 G2485 (.A1(W1487), .A2(W1316), .ZN(W4169));
  NANDX1 G2486 (.A1(W662), .A2(W502), .ZN(W939));
  NANDX1 G2487 (.A1(I264), .A2(W564), .ZN(W940));
  NANDX1 G2488 (.A1(I786), .A2(W37), .ZN(W793));
  NANDX1 G2489 (.A1(W1121), .A2(W581), .ZN(W4172));
  NANDX1 G2490 (.A1(W2329), .A2(W3672), .ZN(W3825));
  NANDX1 G2491 (.A1(W1838), .A2(W946), .ZN(W3747));
  NANDX1 G2492 (.A1(W1307), .A2(W3503), .ZN(O766));
  NANDX1 G2493 (.A1(W173), .A2(I508), .ZN(W944));
  NANDX1 G2494 (.A1(I812), .A2(I376), .ZN(W792));
  NANDX1 G2495 (.A1(I556), .A2(I541), .ZN(W791));
  NANDX1 G2496 (.A1(W748), .A2(I990), .ZN(W822));
  NANDX1 G2497 (.A1(W2503), .A2(W2300), .ZN(W4178));
  NANDX1 G2498 (.A1(W1579), .A2(W2884), .ZN(W4182));
  NANDX1 G2499 (.A1(W1560), .A2(W2465), .ZN(W3745));
  NANDX1 G2500 (.A1(W736), .A2(W1780), .ZN(O572));
  NANDX1 G2501 (.A1(W1604), .A2(W2645), .ZN(W3742));
  NANDX1 G2502 (.A1(W84), .A2(W676), .ZN(W831));
  NANDX1 G2503 (.A1(W815), .A2(W309), .ZN(W4235));
  NANDX1 G2504 (.A1(W969), .A2(I587), .ZN(O718));
  NANDX1 G2505 (.A1(W2248), .A2(W3400), .ZN(O563));
  NANDX1 G2506 (.A1(I203), .A2(I244), .ZN(W779));
  NANDX1 G2507 (.A1(W850), .A2(W2868), .ZN(O800));
  NANDX1 G2508 (.A1(I280), .A2(W565), .ZN(W912));
  NANDX1 G2509 (.A1(W2079), .A2(W785), .ZN(W4239));
  NANDX1 G2510 (.A1(W1209), .A2(W3695), .ZN(O562));
  NANDX1 G2511 (.A1(I204), .A2(I734), .ZN(O799));
  NANDX1 G2512 (.A1(W856), .A2(W2410), .ZN(O802));
  NANDX1 G2513 (.A1(I909), .A2(I241), .ZN(W3716));
  NANDX1 G2514 (.A1(I844), .A2(W2007), .ZN(O803));
  NANDX1 G2515 (.A1(W2284), .A2(W1252), .ZN(O561));
  NANDX1 G2516 (.A1(W2796), .A2(W3819), .ZN(W4243));
  NANDX1 G2517 (.A1(I134), .A2(W500), .ZN(O607));
  NANDX1 G2518 (.A1(I444), .A2(I925), .ZN(W776));
  NANDX1 G2519 (.A1(W2388), .A2(W1738), .ZN(W3711));
  NANDX1 G2520 (.A1(W1374), .A2(W3716), .ZN(O791));
  NANDX1 G2521 (.A1(W736), .A2(I456), .ZN(W783));
  NANDX1 G2522 (.A1(I973), .A2(W631), .ZN(W826));
  NANDX1 G2523 (.A1(I530), .A2(W1448), .ZN(O786));
  NANDX1 G2524 (.A1(W1837), .A2(I780), .ZN(O787));
  NANDX1 G2525 (.A1(W1510), .A2(W1454), .ZN(W3729));
  NANDX1 G2526 (.A1(W805), .A2(I889), .ZN(W827));
  NANDX1 G2527 (.A1(W353), .A2(W532), .ZN(W946));
  NANDX1 G2528 (.A1(I272), .A2(W3517), .ZN(O790));
  NANDX1 G2529 (.A1(W519), .A2(W645), .ZN(W794));
  NANDX1 G2530 (.A1(I681), .A2(I186), .ZN(O792));
  NANDX1 G2531 (.A1(I170), .A2(I128), .ZN(W828));
  NANDX1 G2532 (.A1(W1007), .A2(I682), .ZN(O793));
  NANDX1 G2533 (.A1(W519), .A2(W531), .ZN(W780));
  NANDX1 G2534 (.A1(I402), .A2(I675), .ZN(W829));
  NANDX1 G2535 (.A1(W1268), .A2(W927), .ZN(W3721));
  NANDX1 G2536 (.A1(W3017), .A2(W3417), .ZN(O797));
  NANDX1 G2537 (.A1(W295), .A2(W892), .ZN(W924));
  NANDX1 G2538 (.A1(I600), .A2(W3765), .ZN(O744));
  NANDX1 G2539 (.A1(W3107), .A2(W888), .ZN(W3810));
  NANDX1 G2540 (.A1(W2999), .A2(W4074), .ZN(W4130));
  NANDX1 G2541 (.A1(W807), .A2(I666), .ZN(W818));
  NANDX1 G2542 (.A1(W633), .A2(W893), .ZN(W1009));
  NANDX1 G2543 (.A1(W1001), .A2(I646), .ZN(W3809));
  NANDX1 G2544 (.A1(W259), .A2(W2042), .ZN(W3806));
  NANDX1 G2545 (.A1(W799), .A2(W567), .ZN(W819));
  NANDX1 G2546 (.A1(W203), .A2(I910), .ZN(W923));
  NANDX1 G2547 (.A1(W2655), .A2(W3243), .ZN(O730));
  NANDX1 G2548 (.A1(W2098), .A2(W1429), .ZN(O597));
  NANDX1 G2549 (.A1(W643), .A2(W1217), .ZN(W4134));
  NANDX1 G2550 (.A1(W3494), .A2(W1566), .ZN(W4136));
  NANDX1 G2551 (.A1(W499), .A2(W279), .ZN(W803));
  NANDX1 G2552 (.A1(W149), .A2(W138), .ZN(O28));
  NANDX1 G2553 (.A1(I408), .A2(W88), .ZN(W802));
  NANDX1 G2554 (.A1(W256), .A2(I432), .ZN(W4141));
  NANDX1 G2555 (.A1(W2134), .A2(W1847), .ZN(O739));
  NANDX1 G2556 (.A1(W3967), .A2(W1756), .ZN(W4101));
  NANDX1 G2557 (.A1(W200), .A2(W2385), .ZN(W3815));
  NANDX1 G2558 (.A1(I693), .A2(W796), .ZN(W813));
  NANDX1 G2559 (.A1(W3813), .A2(W1649), .ZN(O734));
  NANDX1 G2560 (.A1(W678), .A2(I872), .ZN(W812));
  NANDX1 G2561 (.A1(W2159), .A2(I660), .ZN(W3814));
  NANDX1 G2562 (.A1(W3182), .A2(W280), .ZN(W4109));
  NANDX1 G2563 (.A1(W1770), .A2(W496), .ZN(W4112));
  NANDX1 G2564 (.A1(W1269), .A2(I692), .ZN(O595));
  NANDX1 G2565 (.A1(W1041), .A2(W1844), .ZN(O732));
  NANDX1 G2566 (.A1(W1744), .A2(W2979), .ZN(W4115));
  NANDX1 G2567 (.A1(W1993), .A2(W4081), .ZN(O741));
  NANDX1 G2568 (.A1(W3407), .A2(W1397), .ZN(W4118));
  NANDX1 G2569 (.A1(I121), .A2(I446), .ZN(W810));
  NANDX1 G2570 (.A1(W3525), .A2(W2217), .ZN(W4121));
  NANDX1 G2571 (.A1(W1227), .A2(W351), .ZN(O743));
  NANDX1 G2572 (.A1(I290), .A2(W294), .ZN(W934));
  NANDX1 G2573 (.A1(W1861), .A2(W3874), .ZN(W4150));
  NANDX1 G2574 (.A1(W1855), .A2(W2255), .ZN(O754));
  NANDX1 G2575 (.A1(W2316), .A2(W3079), .ZN(W3819));
  NANDX1 G2576 (.A1(W3071), .A2(W327), .ZN(O756));
  NANDX1 G2577 (.A1(I116), .A2(W1839), .ZN(W3763));
  NANDX1 G2578 (.A1(W3636), .A2(I584), .ZN(O757));
  NANDX1 G2579 (.A1(W1112), .A2(W2893), .ZN(O582));
  NANDX1 G2580 (.A1(W872), .A2(W1), .ZN(O758));
  NANDX1 G2581 (.A1(W2332), .A2(I88), .ZN(W4088));
  NANDX1 G2582 (.A1(I937), .A2(W2378), .ZN(O760));
  NANDX1 G2583 (.A1(W1784), .A2(W2783), .ZN(W4159));
  NANDX1 G2584 (.A1(I223), .A2(W2931), .ZN(W3759));
  NANDX1 G2585 (.A1(W1056), .A2(W1069), .ZN(W4161));
  NANDX1 G2586 (.A1(W1851), .A2(W2721), .ZN(O580));
  NANDX1 G2587 (.A1(I20), .A2(W664), .ZN(W795));
  NANDX1 G2588 (.A1(W1824), .A2(W2040), .ZN(O577));
  NANDX1 G2589 (.A1(I833), .A2(W1632), .ZN(O604));
  NANDX1 G2590 (.A1(W295), .A2(I224), .ZN(W930));
  NANDX1 G2591 (.A1(I982), .A2(W2291), .ZN(W3797));
  NANDX1 G2592 (.A1(W3346), .A2(W1520), .ZN(W3796));
  NANDX1 G2593 (.A1(W2235), .A2(W799), .ZN(O594));
  NANDX1 G2594 (.A1(W3543), .A2(W1355), .ZN(W4144));
  NANDX1 G2595 (.A1(W515), .A2(W2531), .ZN(W3794));
  NANDX1 G2596 (.A1(W1757), .A2(W525), .ZN(W3792));
  NANDX1 G2597 (.A1(W48), .A2(W1151), .ZN(O591));
  NANDX1 G2598 (.A1(I848), .A2(W688), .ZN(W928));
  NANDX1 G2599 (.A1(W3186), .A2(W87), .ZN(O608));
  NANDX1 G2600 (.A1(W2093), .A2(W3013), .ZN(W3778));
  NANDX1 G2601 (.A1(W2645), .A2(W2438), .ZN(W3773));
  NANDX1 G2602 (.A1(W2393), .A2(W1932), .ZN(W4148));
  NANDX1 G2603 (.A1(W1653), .A2(W382), .ZN(W3768));
  NANDX1 G2604 (.A1(W3123), .A2(W1460), .ZN(W4149));
  NANDX1 G2605 (.A1(I262), .A2(W2977), .ZN(O584));
  NANDX1 G2606 (.A1(W368), .A2(W3771), .ZN(W3818));
  NANDX1 G2607 (.A1(W1338), .A2(W3665), .ZN(O615));
  NANDX1 G2608 (.A1(W372), .A2(I944), .ZN(W745));
  NANDX1 G2609 (.A1(I206), .A2(W3119), .ZN(W4348));
  NANDX1 G2610 (.A1(W86), .A2(I821), .ZN(W744));
  NANDX1 G2611 (.A1(W1325), .A2(I966), .ZN(W4029));
  NANDX1 G2612 (.A1(W59), .A2(W3914), .ZN(W4354));
  NANDX1 G2613 (.A1(W2454), .A2(W1655), .ZN(W4028));
  NANDX1 G2614 (.A1(W2618), .A2(W3361), .ZN(O549));
  NANDX1 G2615 (.A1(W3134), .A2(W3374), .ZN(W3673));
  NANDX1 G2616 (.A1(W476), .A2(W1722), .ZN(O551));
  NANDX1 G2617 (.A1(W43), .A2(I636), .ZN(W743));
  NANDX1 G2618 (.A1(W8), .A2(I132), .ZN(W741));
  NANDX1 G2619 (.A1(W1336), .A2(W1438), .ZN(W4361));
  NANDX1 G2620 (.A1(I136), .A2(W924), .ZN(W962));
  NANDX1 G2621 (.A1(W3564), .A2(W4162), .ZN(W4362));
  NANDX1 G2622 (.A1(W400), .A2(W644), .ZN(W844));
  NANDX1 G2623 (.A1(W2181), .A2(W1566), .ZN(O546));
  NANDX1 G2624 (.A1(W2359), .A2(W928), .ZN(O545));
  NANDX1 G2625 (.A1(W1823), .A2(W1844), .ZN(W4035));
  NANDX1 G2626 (.A1(W2836), .A2(W3183), .ZN(W4329));
  NANDX1 G2627 (.A1(W1245), .A2(W1345), .ZN(W4335));
  NANDX1 G2628 (.A1(W676), .A2(I132), .ZN(W957));
  NANDX1 G2629 (.A1(W2715), .A2(W3084), .ZN(W3688));
  NANDX1 G2630 (.A1(W441), .A2(W2380), .ZN(W3849));
  NANDX1 G2631 (.A1(W256), .A2(W672), .ZN(W841));
  NANDX1 G2632 (.A1(W3078), .A2(W1867), .ZN(O554));
  NANDX1 G2633 (.A1(W2423), .A2(W3548), .ZN(O833));
  NANDX1 G2634 (.A1(W2155), .A2(W3385), .ZN(W4363));
  NANDX1 G2635 (.A1(W2798), .A2(W3283), .ZN(O834));
  NANDX1 G2636 (.A1(I36), .A2(W2339), .ZN(O699));
  NANDX1 G2637 (.A1(W1347), .A2(W1985), .ZN(W3682));
  NANDX1 G2638 (.A1(W2924), .A2(W3128), .ZN(O836));
  NANDX1 G2639 (.A1(W1384), .A2(W88), .ZN(W4342));
  NANDX1 G2640 (.A1(W2006), .A2(I342), .ZN(O698));
  NANDX1 G2641 (.A1(W3888), .A2(I439), .ZN(O837));
  NANDX1 G2642 (.A1(W132), .A2(W84), .ZN(W746));
  NANDX1 G2643 (.A1(I91), .A2(I831), .ZN(O856));
  NANDX1 G2644 (.A1(W509), .A2(W1262), .ZN(O853));
  NANDX1 G2645 (.A1(W1315), .A2(I862), .ZN(O854));
  NANDX1 G2646 (.A1(I923), .A2(I120), .ZN(W731));
  NANDX1 G2647 (.A1(I160), .A2(W2179), .ZN(O693));
  NANDX1 G2648 (.A1(W1500), .A2(W2144), .ZN(W3653));
  NANDX1 G2649 (.A1(W118), .A2(W284), .ZN(W729));
  NANDX1 G2650 (.A1(W101), .A2(I888), .ZN(W4394));
  NANDX1 G2651 (.A1(W3841), .A2(W3673), .ZN(W4399));
  NANDX1 G2652 (.A1(W3270), .A2(I705), .ZN(O543));
  NANDX1 G2653 (.A1(I683), .A2(W9), .ZN(W816));
  NANDX1 G2654 (.A1(W3742), .A2(W847), .ZN(O860));
  NANDX1 G2655 (.A1(W2449), .A2(W2282), .ZN(O861));
  NANDX1 G2656 (.A1(I721), .A2(I203), .ZN(O862));
  NANDX1 G2657 (.A1(W1069), .A2(I353), .ZN(O863));
  NANDX1 G2658 (.A1(I210), .A2(W3957), .ZN(O864));
  NANDX1 G2659 (.A1(W2106), .A2(W3624), .ZN(O692));
  NANDX1 G2660 (.A1(W110), .A2(W437), .ZN(W726));
  NANDX1 G2661 (.A1(I170), .A2(W1636), .ZN(W4378));
  NANDX1 G2662 (.A1(I288), .A2(W1564), .ZN(O619));
  NANDX1 G2663 (.A1(W2330), .A2(W4130), .ZN(W4368));
  NANDX1 G2664 (.A1(W993), .A2(W536), .ZN(O847));
  NANDX1 G2665 (.A1(I665), .A2(W275), .ZN(W738));
  NANDX1 G2666 (.A1(W3458), .A2(W204), .ZN(O848));
  NANDX1 G2667 (.A1(W3062), .A2(I904), .ZN(W3665));
  NANDX1 G2668 (.A1(W965), .A2(W2309), .ZN(W4373));
  NANDX1 G2669 (.A1(I655), .A2(W699), .ZN(W737));
  NANDX1 G2670 (.A1(W695), .A2(W3169), .ZN(O830));
  NANDX1 G2671 (.A1(W396), .A2(W15), .ZN(W964));
  NANDX1 G2672 (.A1(I788), .A2(I437), .ZN(W736));
  NANDX1 G2673 (.A1(W3308), .A2(I414), .ZN(O695));
  NANDX1 G2674 (.A1(W2274), .A2(W2420), .ZN(W3657));
  NANDX1 G2675 (.A1(W650), .A2(W1341), .ZN(W3656));
  NANDX1 G2676 (.A1(I481), .A2(I557), .ZN(W4021));
  NANDX1 G2677 (.A1(W3610), .A2(W943), .ZN(O851));
  NANDX1 G2678 (.A1(I633), .A2(W2467), .ZN(W4283));
  NANDX1 G2679 (.A1(I23), .A2(W1581), .ZN(W4268));
  NANDX1 G2680 (.A1(W1154), .A2(W1640), .ZN(O811));
  NANDX1 G2681 (.A1(I174), .A2(W509), .ZN(O812));
  NANDX1 G2682 (.A1(W584), .A2(W1645), .ZN(W4274));
  NANDX1 G2683 (.A1(W2183), .A2(W3639), .ZN(W3706));
  NANDX1 G2684 (.A1(W2665), .A2(W873), .ZN(W4276));
  NANDX1 G2685 (.A1(W106), .A2(I224), .ZN(W765));
  NANDX1 G2686 (.A1(W3110), .A2(W1911), .ZN(W4282));
  NANDX1 G2687 (.A1(W1442), .A2(W1222), .ZN(O712));
  NANDX1 G2688 (.A1(W3338), .A2(W2307), .ZN(W3840));
  NANDX1 G2689 (.A1(W1133), .A2(W3601), .ZN(W4053));
  NANDX1 G2690 (.A1(W601), .A2(W3709), .ZN(W4284));
  NANDX1 G2691 (.A1(W1685), .A2(W3771), .ZN(W4052));
  NANDX1 G2692 (.A1(W805), .A2(W662), .ZN(W950));
  NANDX1 G2693 (.A1(W622), .A2(W2018), .ZN(W3704));
  NANDX1 G2694 (.A1(W500), .A2(W68), .ZN(W764));
  NANDX1 G2695 (.A1(W3979), .A2(W2703), .ZN(O815));
  NANDX1 G2696 (.A1(W326), .A2(I58), .ZN(W832));
  NANDX1 G2697 (.A1(W2058), .A2(W2), .ZN(W4247));
  NANDX1 G2698 (.A1(W735), .A2(I544), .ZN(W775));
  NANDX1 G2699 (.A1(W3377), .A2(I820), .ZN(W3710));
  NANDX1 G2700 (.A1(W1264), .A2(I338), .ZN(W4065));
  NANDX1 G2701 (.A1(W212), .A2(W798), .ZN(W911));
  NANDX1 G2702 (.A1(W2974), .A2(W2977), .ZN(W3837));
  NANDX1 G2703 (.A1(W412), .A2(W154), .ZN(W4254));
  NANDX1 G2704 (.A1(W1709), .A2(W1827), .ZN(W4260));
  NANDX1 G2705 (.A1(W645), .A2(W3999), .ZN(O709));
  NANDX1 G2706 (.A1(W361), .A2(W2149), .ZN(W4061));
  NANDX1 G2707 (.A1(W860), .A2(I887), .ZN(W949));
  NANDX1 G2708 (.A1(W4250), .A2(W580), .ZN(O809));
  NANDX1 G2709 (.A1(W2478), .A2(W65), .ZN(W3707));
  NANDX1 G2710 (.A1(I809), .A2(W652), .ZN(W769));
  NANDX1 G2711 (.A1(I13), .A2(W3130), .ZN(O715));
  NANDX1 G2712 (.A1(W3122), .A2(W2062), .ZN(O810));
  NANDX1 G2713 (.A1(W1041), .A2(W3652), .ZN(W4317));
  NANDX1 G2714 (.A1(I469), .A2(I290), .ZN(O613));
  NANDX1 G2715 (.A1(W324), .A2(W78), .ZN(W752));
  NANDX1 G2716 (.A1(W796), .A2(I647), .ZN(W4046));
  NANDX1 G2717 (.A1(I983), .A2(I175), .ZN(W953));
  NANDX1 G2718 (.A1(I402), .A2(W2779), .ZN(O706));
  NANDX1 G2719 (.A1(W1253), .A2(I817), .ZN(W4041));
  NANDX1 G2720 (.A1(W1035), .A2(W3259), .ZN(O826));
  NANDX1 G2721 (.A1(W206), .A2(W540), .ZN(W840));
  NANDX1 G2722 (.A1(W2490), .A2(W3408), .ZN(O822));
  NANDX1 G2723 (.A1(W81), .A2(W2261), .ZN(O827));
  NANDX1 G2724 (.A1(W2616), .A2(W2117), .ZN(W4320));
  NANDX1 G2725 (.A1(W1673), .A2(W15), .ZN(W3847));
  NANDX1 G2726 (.A1(W3144), .A2(I368), .ZN(W4321));
  NANDX1 G2727 (.A1(W4300), .A2(W559), .ZN(W4322));
  NANDX1 G2728 (.A1(W899), .A2(W4305), .ZN(W4323));
  NANDX1 G2729 (.A1(W508), .A2(I636), .ZN(W956));
  NANDX1 G2730 (.A1(W3656), .A2(I163), .ZN(O828));
  NANDX1 G2731 (.A1(W3884), .A2(W1155), .ZN(W4298));
  NANDX1 G2732 (.A1(I488), .A2(I636), .ZN(O816));
  NANDX1 G2733 (.A1(I357), .A2(W504), .ZN(O26));
  NANDX1 G2734 (.A1(W275), .A2(I659), .ZN(W3701));
  NANDX1 G2735 (.A1(W205), .A2(W138), .ZN(W761));
  NANDX1 G2736 (.A1(W1263), .A2(W1597), .ZN(W4295));
  NANDX1 G2737 (.A1(W2399), .A2(W2211), .ZN(O559));
  NANDX1 G2738 (.A1(I253), .A2(W1879), .ZN(W3699));
  NANDX1 G2739 (.A1(W2139), .A2(W140), .ZN(W3841));
  NANDX1 G2740 (.A1(W3661), .A2(W4037), .ZN(O865));
  NANDX1 G2741 (.A1(W2996), .A2(I181), .ZN(W4300));
  NANDX1 G2742 (.A1(W897), .A2(W333), .ZN(W907));
  NANDX1 G2743 (.A1(I786), .A2(W363), .ZN(W756));
  NANDX1 G2744 (.A1(W493), .A2(I475), .ZN(W4305));
  NANDX1 G2745 (.A1(I402), .A2(W331), .ZN(W755));
  NANDX1 G2746 (.A1(I530), .A2(W228), .ZN(W754));
  NANDX1 G2747 (.A1(W215), .A2(I567), .ZN(W952));
  NANDX1 G2748 (.A1(W4251), .A2(W4198), .ZN(O1911));
  NANDX1 G2749 (.A1(I422), .A2(I423), .ZN(W211));
  NANDX1 G2750 (.A1(W1376), .A2(W4758), .ZN(O1889));
  NANDX1 G2751 (.A1(W5767), .A2(W632), .ZN(O1891));
  NANDX1 G2752 (.A1(W873), .A2(W2398), .ZN(W5910));
  NANDX1 G2753 (.A1(W670), .A2(W5301), .ZN(O1895));
  NANDX1 G2754 (.A1(W4386), .A2(W2488), .ZN(O1897));
  NANDX1 G2755 (.A1(W5564), .A2(W5674), .ZN(O1901));
  NANDX1 G2756 (.A1(W4895), .A2(W325), .ZN(O1903));
  NANDX1 G2757 (.A1(W2419), .A2(W152), .ZN(O1904));
  NANDX1 G2758 (.A1(W2356), .A2(W852), .ZN(O1906));
  NANDX1 G2759 (.A1(W1986), .A2(W2218), .ZN(O1909));
  NANDX1 G2760 (.A1(W627), .A2(W3187), .ZN(O1885));
  NANDX1 G2761 (.A1(W3719), .A2(W2993), .ZN(O1913));
  NANDX1 G2762 (.A1(I408), .A2(I409), .ZN(W204));
  NANDX1 G2763 (.A1(W4553), .A2(W153), .ZN(O1915));
  NANDX1 G2764 (.A1(I404), .A2(I405), .ZN(W202));
  NANDX1 G2765 (.A1(W1945), .A2(W2709), .ZN(O1917));
  NANDX1 G2766 (.A1(I970), .A2(W3801), .ZN(O1918));
  NANDX1 G2767 (.A1(W3980), .A2(W975), .ZN(O1923));
  NANDX1 G2768 (.A1(W5218), .A2(W3171), .ZN(O1925));
  NANDX1 G2769 (.A1(W3691), .A2(W1843), .ZN(O1927));
  NANDX1 G2770 (.A1(W218), .A2(W3622), .ZN(O1930));
  NANDX1 G2771 (.A1(W5144), .A2(W2355), .ZN(O1931));
  NANDX1 G2772 (.A1(W1462), .A2(W1636), .ZN(O1859));
  NANDX1 G2773 (.A1(W385), .A2(W4627), .ZN(O1843));
  NANDX1 G2774 (.A1(W337), .A2(W4024), .ZN(O1844));
  NANDX1 G2775 (.A1(W672), .A2(W601), .ZN(W5855));
  NANDX1 G2776 (.A1(W3248), .A2(W1579), .ZN(O1846));
  NANDX1 G2777 (.A1(W5399), .A2(W3865), .ZN(O1847));
  NANDX1 G2778 (.A1(I456), .A2(I457), .ZN(W228));
  NANDX1 G2779 (.A1(W840), .A2(W3166), .ZN(W5863));
  NANDX1 G2780 (.A1(W1240), .A2(W5496), .ZN(O1852));
  NANDX1 G2781 (.A1(I450), .A2(I451), .ZN(W225));
  NANDX1 G2782 (.A1(W3813), .A2(W4120), .ZN(O1854));
  NANDX1 G2783 (.A1(W1045), .A2(W4694), .ZN(O1857));
  NANDX1 G2784 (.A1(I910), .A2(W3520), .ZN(O1934));
  NANDX1 G2785 (.A1(W3288), .A2(W597), .ZN(O1863));
  NANDX1 G2786 (.A1(W3796), .A2(W5233), .ZN(O1864));
  NANDX1 G2787 (.A1(W1666), .A2(W50), .ZN(O1867));
  NANDX1 G2788 (.A1(W5121), .A2(W2420), .ZN(O1868));
  NANDX1 G2789 (.A1(I438), .A2(I439), .ZN(W219));
  NANDX1 G2790 (.A1(I436), .A2(I437), .ZN(W218));
  NANDX1 G2791 (.A1(W1630), .A2(I471), .ZN(W5891));
  NANDX1 G2792 (.A1(W4003), .A2(W4320), .ZN(O1876));
  NANDX1 G2793 (.A1(I432), .A2(I433), .ZN(W216));
  NANDX1 G2794 (.A1(W4128), .A2(I707), .ZN(O1878));
  NANDX1 G2795 (.A1(I428), .A2(I429), .ZN(W214));
  NANDX1 G2796 (.A1(W4092), .A2(W3563), .ZN(O1993));
  NANDX1 G2797 (.A1(W6006), .A2(W2471), .ZN(O1981));
  NANDX1 G2798 (.A1(W5506), .A2(I8), .ZN(O1982));
  NANDX1 G2799 (.A1(W410), .A2(W3929), .ZN(O1983));
  NANDX1 G2800 (.A1(W5547), .A2(W1660), .ZN(O1984));
  NANDX1 G2801 (.A1(W2148), .A2(W5298), .ZN(O1985));
  NANDX1 G2802 (.A1(W965), .A2(W2443), .ZN(O1986));
  NANDX1 G2803 (.A1(I360), .A2(I361), .ZN(W180));
  NANDX1 G2804 (.A1(W5763), .A2(W1028), .ZN(O1987));
  NANDX1 G2805 (.A1(W4897), .A2(W2733), .ZN(O1989));
  NANDX1 G2806 (.A1(I356), .A2(I357), .ZN(W178));
  NANDX1 G2807 (.A1(I354), .A2(I355), .ZN(W177));
  NANDX1 G2808 (.A1(W5066), .A2(W1458), .ZN(W6006));
  NANDX1 G2809 (.A1(I352), .A2(I353), .ZN(W176));
  NANDX1 G2810 (.A1(W4859), .A2(W4268), .ZN(O1995));
  NANDX1 G2811 (.A1(I350), .A2(I351), .ZN(W175));
  NANDX1 G2812 (.A1(W3991), .A2(W3535), .ZN(O1997));
  NANDX1 G2813 (.A1(I348), .A2(I349), .ZN(W174));
  NANDX1 G2814 (.A1(W2515), .A2(W1361), .ZN(O2002));
  NANDX1 G2815 (.A1(W4909), .A2(W1929), .ZN(O2004));
  NANDX1 G2816 (.A1(W3123), .A2(W4405), .ZN(O2013));
  NANDX1 G2817 (.A1(W2252), .A2(W3306), .ZN(O2015));
  NANDX1 G2818 (.A1(W4259), .A2(W3848), .ZN(O2016));
  NANDX1 G2819 (.A1(W4267), .A2(W4036), .ZN(O2017));
  NANDX1 G2820 (.A1(W378), .A2(W4521), .ZN(O1954));
  NANDX1 G2821 (.A1(I392), .A2(I393), .ZN(W196));
  NANDX1 G2822 (.A1(I390), .A2(I391), .ZN(W195));
  NANDX1 G2823 (.A1(I388), .A2(I389), .ZN(W194));
  NANDX1 G2824 (.A1(I386), .A2(I387), .ZN(W193));
  NANDX1 G2825 (.A1(W2696), .A2(W375), .ZN(O1943));
  NANDX1 G2826 (.A1(W4827), .A2(I166), .ZN(W5968));
  NANDX1 G2827 (.A1(W1777), .A2(I13), .ZN(O1947));
  NANDX1 G2828 (.A1(W978), .A2(W3337), .ZN(O1948));
  NANDX1 G2829 (.A1(W1457), .A2(W1201), .ZN(O1949));
  NANDX1 G2830 (.A1(W3162), .A2(I939), .ZN(O1951));
  NANDX1 G2831 (.A1(W1596), .A2(W732), .ZN(O1953));
  NANDX1 G2832 (.A1(W3431), .A2(I493), .ZN(O1842));
  NANDX1 G2833 (.A1(W1433), .A2(W2660), .ZN(O1957));
  NANDX1 G2834 (.A1(W4366), .A2(W4430), .ZN(O1958));
  NANDX1 G2835 (.A1(W1368), .A2(W4015), .ZN(W5987));
  NANDX1 G2836 (.A1(I502), .A2(W825), .ZN(O1962));
  NANDX1 G2837 (.A1(W1566), .A2(W4904), .ZN(O1963));
  NANDX1 G2838 (.A1(I370), .A2(I371), .ZN(W185));
  NANDX1 G2839 (.A1(W1255), .A2(W800), .ZN(O1969));
  NANDX1 G2840 (.A1(I792), .A2(W3708), .ZN(O1970));
  NANDX1 G2841 (.A1(W3294), .A2(W3964), .ZN(O1972));
  NANDX1 G2842 (.A1(W1492), .A2(W3420), .ZN(O1976));
  NANDX1 G2843 (.A1(W4656), .A2(W3890), .ZN(O1977));
  NANDX1 G2844 (.A1(W5710), .A2(W5225), .ZN(W5725));
  NANDX1 G2845 (.A1(W1825), .A2(W2012), .ZN(W5686));
  NANDX1 G2846 (.A1(W1813), .A2(W4170), .ZN(O1700));
  NANDX1 G2847 (.A1(W2987), .A2(W962), .ZN(O1707));
  NANDX1 G2848 (.A1(I564), .A2(I565), .ZN(W282));
  NANDX1 G2849 (.A1(I21), .A2(W174), .ZN(W5698));
  NANDX1 G2850 (.A1(W1542), .A2(W4927), .ZN(O1710));
  NANDX1 G2851 (.A1(W3383), .A2(W1179), .ZN(O1713));
  NANDX1 G2852 (.A1(W2290), .A2(W919), .ZN(O1714));
  NANDX1 G2853 (.A1(W5404), .A2(W982), .ZN(O1724));
  NANDX1 G2854 (.A1(I542), .A2(I543), .ZN(W271));
  NANDX1 G2855 (.A1(I536), .A2(I537), .ZN(W268));
  NANDX1 G2856 (.A1(I574), .A2(I575), .ZN(W287));
  NANDX1 G2857 (.A1(I534), .A2(I535), .ZN(W267));
  NANDX1 G2858 (.A1(I532), .A2(I533), .ZN(W266));
  NANDX1 G2859 (.A1(W1220), .A2(I872), .ZN(O1740));
  NANDX1 G2860 (.A1(W876), .A2(W3447), .ZN(O1742));
  NANDX1 G2861 (.A1(W2894), .A2(W2766), .ZN(O1745));
  NANDX1 G2862 (.A1(W2030), .A2(W1359), .ZN(W5748));
  NANDX1 G2863 (.A1(W2564), .A2(W834), .ZN(O1757));
  NANDX1 G2864 (.A1(I304), .A2(W3100), .ZN(O1758));
  NANDX1 G2865 (.A1(W5454), .A2(W3826), .ZN(O1759));
  NANDX1 G2866 (.A1(W3247), .A2(W1826), .ZN(O1761));
  NANDX1 G2867 (.A1(W3005), .A2(W986), .ZN(O1763));
  NANDX1 G2868 (.A1(I596), .A2(I597), .ZN(W298));
  NANDX1 G2869 (.A1(I608), .A2(I609), .ZN(W304));
  NANDX1 G2870 (.A1(I508), .A2(W4317), .ZN(O1663));
  NANDX1 G2871 (.A1(W4121), .A2(W5484), .ZN(O1666));
  NANDX1 G2872 (.A1(I738), .A2(W3223), .ZN(O1667));
  NANDX1 G2873 (.A1(I604), .A2(I605), .ZN(O3));
  NANDX1 G2874 (.A1(W5208), .A2(W3441), .ZN(O1669));
  NANDX1 G2875 (.A1(W3497), .A2(W2951), .ZN(O1671));
  NANDX1 G2876 (.A1(I602), .A2(I603), .ZN(W301));
  NANDX1 G2877 (.A1(W1036), .A2(W3293), .ZN(O1673));
  NANDX1 G2878 (.A1(W4172), .A2(W512), .ZN(O1674));
  NANDX1 G2879 (.A1(I600), .A2(I601), .ZN(W300));
  NANDX1 G2880 (.A1(W2908), .A2(W373), .ZN(O1768));
  NANDX1 G2881 (.A1(I594), .A2(I595), .ZN(W297));
  NANDX1 G2882 (.A1(W2376), .A2(W3985), .ZN(O1679));
  NANDX1 G2883 (.A1(W2443), .A2(W895), .ZN(O1680));
  NANDX1 G2884 (.A1(W2058), .A2(W4559), .ZN(W5662));
  NANDX1 G2885 (.A1(W450), .A2(W2068), .ZN(W5665));
  NANDX1 G2886 (.A1(W4079), .A2(W5351), .ZN(W5666));
  NANDX1 G2887 (.A1(W886), .A2(I164), .ZN(O1687));
  NANDX1 G2888 (.A1(I586), .A2(I587), .ZN(W293));
  NANDX1 G2889 (.A1(W413), .A2(W3844), .ZN(O1692));
  NANDX1 G2890 (.A1(I580), .A2(I581), .ZN(W290));
  NANDX1 G2891 (.A1(W4700), .A2(W5529), .ZN(O1695));
  NANDX1 G2892 (.A1(I474), .A2(I475), .ZN(W237));
  NANDX1 G2893 (.A1(W5084), .A2(I817), .ZN(O1804));
  NANDX1 G2894 (.A1(W5627), .A2(W4747), .ZN(O1808));
  NANDX1 G2895 (.A1(W3309), .A2(W608), .ZN(O1810));
  NANDX1 G2896 (.A1(W639), .A2(W2197), .ZN(O1812));
  NANDX1 G2897 (.A1(W916), .A2(W1362), .ZN(W5815));
  NANDX1 G2898 (.A1(I482), .A2(I483), .ZN(W241));
  NANDX1 G2899 (.A1(W4622), .A2(I874), .ZN(O1815));
  NANDX1 G2900 (.A1(W3674), .A2(W772), .ZN(O1816));
  NANDX1 G2901 (.A1(W301), .A2(W4554), .ZN(W5820));
  NANDX1 G2902 (.A1(I478), .A2(I479), .ZN(W239));
  NANDX1 G2903 (.A1(I476), .A2(I477), .ZN(W238));
  NANDX1 G2904 (.A1(I488), .A2(I489), .ZN(W244));
  NANDX1 G2905 (.A1(I470), .A2(I471), .ZN(W235));
  NANDX1 G2906 (.A1(W1613), .A2(W5766), .ZN(O1821));
  NANDX1 G2907 (.A1(W1702), .A2(W1261), .ZN(O1827));
  NANDX1 G2908 (.A1(W1925), .A2(W1507), .ZN(O1829));
  NANDX1 G2909 (.A1(W743), .A2(W1170), .ZN(O1830));
  NANDX1 G2910 (.A1(W1947), .A2(W4363), .ZN(O1831));
  NANDX1 G2911 (.A1(I842), .A2(W1569), .ZN(O1833));
  NANDX1 G2912 (.A1(W3150), .A2(W1447), .ZN(W5841));
  NANDX1 G2913 (.A1(W1854), .A2(W4584), .ZN(O1836));
  NANDX1 G2914 (.A1(W3319), .A2(W3907), .ZN(O1838));
  NANDX1 G2915 (.A1(W2563), .A2(W5408), .ZN(O1839));
  NANDX1 G2916 (.A1(W560), .A2(W1016), .ZN(O1785));
  NANDX1 G2917 (.A1(W1919), .A2(W1924), .ZN(O1769));
  NANDX1 G2918 (.A1(W1775), .A2(W4934), .ZN(W5766));
  NANDX1 G2919 (.A1(I103), .A2(W3883), .ZN(W5767));
  NANDX1 G2920 (.A1(W5437), .A2(W626), .ZN(O1770));
  NANDX1 G2921 (.A1(W5087), .A2(W4713), .ZN(O1772));
  NANDX1 G2922 (.A1(W2717), .A2(W5381), .ZN(O1774));
  NANDX1 G2923 (.A1(I508), .A2(I509), .ZN(W254));
  NANDX1 G2924 (.A1(I506), .A2(I507), .ZN(W253));
  NANDX1 G2925 (.A1(I504), .A2(I505), .ZN(W252));
  NANDX1 G2926 (.A1(W4856), .A2(W2754), .ZN(O1779));
  NANDX1 G2927 (.A1(W2436), .A2(W1918), .ZN(O1781));
  NANDX1 G2928 (.A1(W1944), .A2(W4789), .ZN(O2020));
  NANDX1 G2929 (.A1(W5076), .A2(W4560), .ZN(O1787));
  NANDX1 G2930 (.A1(I502), .A2(I503), .ZN(W251));
  NANDX1 G2931 (.A1(I500), .A2(I501), .ZN(W250));
  NANDX1 G2932 (.A1(I498), .A2(I499), .ZN(W249));
  NANDX1 G2933 (.A1(W277), .A2(W5253), .ZN(O1792));
  NANDX1 G2934 (.A1(W3297), .A2(W2651), .ZN(O1795));
  NANDX1 G2935 (.A1(W5576), .A2(W2108), .ZN(O1796));
  NANDX1 G2936 (.A1(I490), .A2(I491), .ZN(W245));
  NANDX1 G2937 (.A1(W3529), .A2(W2965), .ZN(O1798));
  NANDX1 G2938 (.A1(W5090), .A2(W2817), .ZN(O1800));
  NANDX1 G2939 (.A1(I116), .A2(I117), .ZN(W58));
  NANDX1 G2940 (.A1(I134), .A2(I135), .ZN(W67));
  NANDX1 G2941 (.A1(W5442), .A2(W5348), .ZN(O2271));
  NANDX1 G2942 (.A1(W3409), .A2(W4258), .ZN(O2272));
  NANDX1 G2943 (.A1(W3349), .A2(I349), .ZN(O2274));
  NANDX1 G2944 (.A1(W3), .A2(W994), .ZN(O2275));
  NANDX1 G2945 (.A1(W3480), .A2(W6226), .ZN(O2276));
  NANDX1 G2946 (.A1(W4508), .A2(I495), .ZN(O2283));
  NANDX1 G2947 (.A1(W5874), .A2(W3486), .ZN(O2284));
  NANDX1 G2948 (.A1(W2724), .A2(W1816), .ZN(O2290));
  NANDX1 G2949 (.A1(W104), .A2(W486), .ZN(O2292));
  NANDX1 G2950 (.A1(W3711), .A2(W3527), .ZN(O2295));
  NANDX1 G2951 (.A1(I136), .A2(I137), .ZN(W68));
  NANDX1 G2952 (.A1(I686), .A2(W5686), .ZN(O2299));
  NANDX1 G2953 (.A1(W2776), .A2(W6055), .ZN(O2306));
  NANDX1 G2954 (.A1(I108), .A2(I109), .ZN(W54));
  NANDX1 G2955 (.A1(I102), .A2(I103), .ZN(W51));
  NANDX1 G2956 (.A1(I94), .A2(I95), .ZN(O0));
  NANDX1 G2957 (.A1(W154), .A2(W3496), .ZN(O2321));
  NANDX1 G2958 (.A1(W5072), .A2(W2132), .ZN(O2322));
  NANDX1 G2959 (.A1(W501), .A2(W4478), .ZN(O2324));
  NANDX1 G2960 (.A1(W6009), .A2(W3396), .ZN(O2328));
  NANDX1 G2961 (.A1(I84), .A2(I85), .ZN(W42));
  NANDX1 G2962 (.A1(W313), .A2(W5482), .ZN(O2331));
  NANDX1 G2963 (.A1(I164), .A2(I165), .ZN(W82));
  NANDX1 G2964 (.A1(I194), .A2(I195), .ZN(W97));
  NANDX1 G2965 (.A1(W3838), .A2(W4851), .ZN(O2204));
  NANDX1 G2966 (.A1(I212), .A2(W4431), .ZN(O2206));
  NANDX1 G2967 (.A1(W3167), .A2(W363), .ZN(O2207));
  NANDX1 G2968 (.A1(W3828), .A2(W3177), .ZN(O2216));
  NANDX1 G2969 (.A1(W4655), .A2(W2624), .ZN(O2219));
  NANDX1 G2970 (.A1(W1102), .A2(W3317), .ZN(O2221));
  NANDX1 G2971 (.A1(W4514), .A2(I416), .ZN(O2226));
  NANDX1 G2972 (.A1(W4766), .A2(W822), .ZN(O2230));
  NANDX1 G2973 (.A1(W1751), .A2(W875), .ZN(W6283));
  NANDX1 G2974 (.A1(W432), .A2(W3793), .ZN(O2236));
  NANDX1 G2975 (.A1(W4212), .A2(I998), .ZN(O2336));
  NANDX1 G2976 (.A1(W6283), .A2(I734), .ZN(O2241));
  NANDX1 G2977 (.A1(I156), .A2(I157), .ZN(W78));
  NANDX1 G2978 (.A1(W5737), .A2(W3215), .ZN(O2246));
  NANDX1 G2979 (.A1(W2454), .A2(I922), .ZN(O2248));
  NANDX1 G2980 (.A1(W2639), .A2(W4877), .ZN(O2251));
  NANDX1 G2981 (.A1(W1408), .A2(W2167), .ZN(O2252));
  NANDX1 G2982 (.A1(W133), .A2(W29), .ZN(O2255));
  NANDX1 G2983 (.A1(W4260), .A2(I11), .ZN(O2256));
  NANDX1 G2984 (.A1(I144), .A2(I145), .ZN(W72));
  NANDX1 G2985 (.A1(W386), .A2(W4164), .ZN(O2258));
  NANDX1 G2986 (.A1(W3044), .A2(W939), .ZN(O2259));
  NANDX1 G2987 (.A1(I22), .A2(I23), .ZN(W11));
  NANDX1 G2988 (.A1(I44), .A2(I45), .ZN(W22));
  NANDX1 G2989 (.A1(W4467), .A2(I28), .ZN(O2387));
  NANDX1 G2990 (.A1(W2709), .A2(W3307), .ZN(O2388));
  NANDX1 G2991 (.A1(W1974), .A2(W4935), .ZN(O2392));
  NANDX1 G2992 (.A1(I38), .A2(I39), .ZN(W19));
  NANDX1 G2993 (.A1(W1040), .A2(W1372), .ZN(O2402));
  NANDX1 G2994 (.A1(W1112), .A2(W2887), .ZN(O2403));
  NANDX1 G2995 (.A1(W4578), .A2(W5637), .ZN(O2412));
  NANDX1 G2996 (.A1(I28), .A2(I29), .ZN(W14));
  NANDX1 G2997 (.A1(W1510), .A2(I476), .ZN(O2415));
  NANDX1 G2998 (.A1(W211), .A2(W4569), .ZN(O2420));
  NANDX1 G2999 (.A1(W1375), .A2(W183), .ZN(O2384));
  NANDX1 G3000 (.A1(W5004), .A2(W516), .ZN(O2423));
  NANDX1 G3001 (.A1(I18), .A2(I19), .ZN(W9));
  NANDX1 G3002 (.A1(I16), .A2(I17), .ZN(W8));
  NANDX1 G3003 (.A1(W2270), .A2(W5282), .ZN(O2434));
  NANDX1 G3004 (.A1(W1509), .A2(W324), .ZN(O2435));
  NANDX1 G3005 (.A1(I12), .A2(I13), .ZN(W6));
  NANDX1 G3006 (.A1(W3515), .A2(I827), .ZN(O2439));
  NANDX1 G3007 (.A1(W980), .A2(I514), .ZN(O2443));
  NANDX1 G3008 (.A1(I4), .A2(I5), .ZN(W2));
  NANDX1 G3009 (.A1(W2025), .A2(W3280), .ZN(O2447));
  NANDX1 G3010 (.A1(I2), .A2(I3), .ZN(W1));
  NANDX1 G3011 (.A1(I191), .A2(W4115), .ZN(O2363));
  NANDX1 G3012 (.A1(I592), .A2(W1873), .ZN(O2338));
  NANDX1 G3013 (.A1(W3291), .A2(W2053), .ZN(O2341));
  NANDX1 G3014 (.A1(W2458), .A2(W4520), .ZN(O2345));
  NANDX1 G3015 (.A1(W3483), .A2(W5185), .ZN(O2347));
  NANDX1 G3016 (.A1(I357), .A2(W3310), .ZN(O2348));
  NANDX1 G3017 (.A1(W5093), .A2(W3547), .ZN(O2349));
  NANDX1 G3018 (.A1(W5615), .A2(W3172), .ZN(O2351));
  NANDX1 G3019 (.A1(W1806), .A2(W1995), .ZN(O2354));
  NANDX1 G3020 (.A1(I687), .A2(W101), .ZN(O2355));
  NANDX1 G3021 (.A1(I60), .A2(I61), .ZN(W30));
  NANDX1 G3022 (.A1(W5121), .A2(W4604), .ZN(O2358));
  NANDX1 G3023 (.A1(I196), .A2(I197), .ZN(W98));
  NANDX1 G3024 (.A1(W3450), .A2(W2984), .ZN(O2364));
  NANDX1 G3025 (.A1(W2805), .A2(I484), .ZN(O2365));
  NANDX1 G3026 (.A1(I184), .A2(I776), .ZN(O2367));
  NANDX1 G3027 (.A1(I947), .A2(W2351), .ZN(O2368));
  NANDX1 G3028 (.A1(I54), .A2(I55), .ZN(W27));
  NANDX1 G3029 (.A1(W6223), .A2(W1255), .ZN(O2371));
  NANDX1 G3030 (.A1(I538), .A2(I387), .ZN(O2374));
  NANDX1 G3031 (.A1(W3409), .A2(W3154), .ZN(O2380));
  NANDX1 G3032 (.A1(W1525), .A2(W4800), .ZN(O2382));
  NANDX1 G3033 (.A1(W3789), .A2(W4179), .ZN(O2383));
  NANDX1 G3034 (.A1(I276), .A2(I277), .ZN(W138));
  NANDX1 G3035 (.A1(W940), .A2(W1038), .ZN(O2063));
  NANDX1 G3036 (.A1(W2113), .A2(W2314), .ZN(O2065));
  NANDX1 G3037 (.A1(W5283), .A2(W1568), .ZN(O2066));
  NANDX1 G3038 (.A1(W4389), .A2(W5454), .ZN(O2071));
  NANDX1 G3039 (.A1(I290), .A2(I291), .ZN(W145));
  NANDX1 G3040 (.A1(W2709), .A2(W4016), .ZN(O2073));
  NANDX1 G3041 (.A1(W5910), .A2(W1153), .ZN(O2074));
  NANDX1 G3042 (.A1(I288), .A2(I289), .ZN(W144));
  NANDX1 G3043 (.A1(I284), .A2(I285), .ZN(W142));
  NANDX1 G3044 (.A1(W58), .A2(I798), .ZN(O2083));
  NANDX1 G3045 (.A1(W4830), .A2(I817), .ZN(O2084));
  NANDX1 G3046 (.A1(I296), .A2(I297), .ZN(W148));
  NANDX1 G3047 (.A1(W758), .A2(W1174), .ZN(O2090));
  NANDX1 G3048 (.A1(W3046), .A2(W4174), .ZN(W6129));
  NANDX1 G3049 (.A1(I268), .A2(I269), .ZN(W134));
  NANDX1 G3050 (.A1(W2397), .A2(W791), .ZN(O2098));
  NANDX1 G3051 (.A1(W5438), .A2(W1184), .ZN(O2103));
  NANDX1 G3052 (.A1(W4922), .A2(I641), .ZN(O2104));
  NANDX1 G3053 (.A1(W3774), .A2(W3113), .ZN(O2105));
  NANDX1 G3054 (.A1(W1081), .A2(W2916), .ZN(O2106));
  NANDX1 G3055 (.A1(W5815), .A2(W116), .ZN(O2107));
  NANDX1 G3056 (.A1(W413), .A2(W5302), .ZN(O2108));
  NANDX1 G3057 (.A1(W3320), .A2(W536), .ZN(O2109));
  NANDX1 G3058 (.A1(W4383), .A2(W1761), .ZN(O2046));
  NANDX1 G3059 (.A1(I328), .A2(I329), .ZN(W164));
  NANDX1 G3060 (.A1(W1370), .A2(W4183), .ZN(W6058));
  NANDX1 G3061 (.A1(I322), .A2(I323), .ZN(W161));
  NANDX1 G3062 (.A1(I318), .A2(I319), .ZN(W159));
  NANDX1 G3063 (.A1(W2122), .A2(W1675), .ZN(O2032));
  NANDX1 G3064 (.A1(I866), .A2(W2471), .ZN(O2034));
  NANDX1 G3065 (.A1(I314), .A2(I315), .ZN(W157));
  NANDX1 G3066 (.A1(W2324), .A2(W4502), .ZN(O2036));
  NANDX1 G3067 (.A1(W5280), .A2(W2238), .ZN(O2037));
  NANDX1 G3068 (.A1(I312), .A2(I313), .ZN(W156));
  NANDX1 G3069 (.A1(I308), .A2(I309), .ZN(W154));
  NANDX1 G3070 (.A1(W2951), .A2(W156), .ZN(O2110));
  NANDX1 G3071 (.A1(W4321), .A2(W5938), .ZN(O2047));
  NANDX1 G3072 (.A1(I304), .A2(I305), .ZN(W152));
  NANDX1 G3073 (.A1(W2426), .A2(W3757), .ZN(O2049));
  NANDX1 G3074 (.A1(W3362), .A2(W193), .ZN(O2050));
  NANDX1 G3075 (.A1(I302), .A2(I303), .ZN(W151));
  NANDX1 G3076 (.A1(I357), .A2(W5253), .ZN(O2053));
  NANDX1 G3077 (.A1(I300), .A2(I301), .ZN(W150));
  NANDX1 G3078 (.A1(W4485), .A2(I965), .ZN(O2056));
  NANDX1 G3079 (.A1(W1655), .A2(W5286), .ZN(O2057));
  NANDX1 G3080 (.A1(W246), .A2(W4021), .ZN(O2059));
  NANDX1 G3081 (.A1(I298), .A2(I299), .ZN(W149));
  NANDX1 G3082 (.A1(W5007), .A2(W1837), .ZN(O2184));
  NANDX1 G3083 (.A1(I683), .A2(W1760), .ZN(O2166));
  NANDX1 G3084 (.A1(I226), .A2(I227), .ZN(W113));
  NANDX1 G3085 (.A1(W3870), .A2(W2171), .ZN(O2168));
  NANDX1 G3086 (.A1(W2512), .A2(W2566), .ZN(O2169));
  NANDX1 G3087 (.A1(W3020), .A2(W2561), .ZN(O2171));
  NANDX1 G3088 (.A1(I222), .A2(I223), .ZN(W111));
  NANDX1 G3089 (.A1(I220), .A2(I221), .ZN(W110));
  NANDX1 G3090 (.A1(W3768), .A2(W3102), .ZN(O2175));
  NANDX1 G3091 (.A1(I214), .A2(I215), .ZN(W107));
  NANDX1 G3092 (.A1(W4303), .A2(W4791), .ZN(O2181));
  NANDX1 G3093 (.A1(W3452), .A2(W4014), .ZN(W6226));
  NANDX1 G3094 (.A1(I228), .A2(I229), .ZN(W114));
  NANDX1 G3095 (.A1(I212), .A2(I213), .ZN(W106));
  NANDX1 G3096 (.A1(W4079), .A2(W4684), .ZN(O2186));
  NANDX1 G3097 (.A1(I51), .A2(W4908), .ZN(O2187));
  NANDX1 G3098 (.A1(W2034), .A2(W4277), .ZN(O2188));
  NANDX1 G3099 (.A1(W3927), .A2(W1623), .ZN(O2189));
  NANDX1 G3100 (.A1(I208), .A2(I209), .ZN(W104));
  NANDX1 G3101 (.A1(W1332), .A2(W3008), .ZN(O2192));
  NANDX1 G3102 (.A1(I206), .A2(I207), .ZN(W103));
  NANDX1 G3103 (.A1(W3546), .A2(I621), .ZN(O2196));
  NANDX1 G3104 (.A1(I202), .A2(I203), .ZN(W101));
  NANDX1 G3105 (.A1(W2434), .A2(I780), .ZN(O2200));
  NANDX1 G3106 (.A1(I732), .A2(I533), .ZN(O2143));
  NANDX1 G3107 (.A1(W1803), .A2(W4740), .ZN(O2113));
  NANDX1 G3108 (.A1(W413), .A2(W1168), .ZN(W6154));
  NANDX1 G3109 (.A1(W1804), .A2(W5122), .ZN(O2114));
  NANDX1 G3110 (.A1(I258), .A2(I259), .ZN(W129));
  NANDX1 G3111 (.A1(I441), .A2(W5511), .ZN(O2118));
  NANDX1 G3112 (.A1(W3811), .A2(W5968), .ZN(O2122));
  NANDX1 G3113 (.A1(W5836), .A2(W5860), .ZN(O2124));
  NANDX1 G3114 (.A1(I254), .A2(I255), .ZN(W127));
  NANDX1 G3115 (.A1(I756), .A2(W1133), .ZN(O2129));
  NANDX1 G3116 (.A1(W5487), .A2(W6087), .ZN(O2134));
  NANDX1 G3117 (.A1(W114), .A2(W4667), .ZN(O2139));
  NANDX1 G3118 (.A1(W2522), .A2(W153), .ZN(W5629));
  NANDX1 G3119 (.A1(I242), .A2(I243), .ZN(W121));
  NANDX1 G3120 (.A1(W3307), .A2(I32), .ZN(O2146));
  NANDX1 G3121 (.A1(I238), .A2(I239), .ZN(W119));
  NANDX1 G3122 (.A1(W6006), .A2(W4732), .ZN(O2149));
  NANDX1 G3123 (.A1(I236), .A2(I237), .ZN(W118));
  NANDX1 G3124 (.A1(W2988), .A2(W798), .ZN(O2151));
  NANDX1 G3125 (.A1(W1455), .A2(I618), .ZN(W6197));
  NANDX1 G3126 (.A1(W5156), .A2(W775), .ZN(O2155));
  NANDX1 G3127 (.A1(W3057), .A2(W1179), .ZN(O2156));
  NANDX1 G3128 (.A1(I232), .A2(I233), .ZN(W116));
  NANDX1 G3129 (.A1(W3462), .A2(W4498), .ZN(W5047));
  NANDX1 G3130 (.A1(W280), .A2(W258), .ZN(W522));
  NANDX1 G3131 (.A1(I55), .A2(W4762), .ZN(O1217));
  NANDX1 G3132 (.A1(I391), .A2(W3213), .ZN(O1219));
  NANDX1 G3133 (.A1(W3968), .A2(W3841), .ZN(W5025));
  NANDX1 G3134 (.A1(W199), .A2(I78), .ZN(W519));
  NANDX1 G3135 (.A1(W2170), .A2(W4293), .ZN(W5028));
  NANDX1 G3136 (.A1(W371), .A2(I150), .ZN(W517));
  NANDX1 G3137 (.A1(W1895), .A2(W1951), .ZN(O1223));
  NANDX1 G3138 (.A1(W1616), .A2(W2080), .ZN(O1227));
  NANDX1 G3139 (.A1(I207), .A2(W4140), .ZN(W5037));
  NANDX1 G3140 (.A1(I814), .A2(W107), .ZN(O1230));
  NANDX1 G3141 (.A1(W4564), .A2(W2284), .ZN(O1214));
  NANDX1 G3142 (.A1(I135), .A2(W2312), .ZN(O1236));
  NANDX1 G3143 (.A1(W2049), .A2(W1822), .ZN(O1237));
  NANDX1 G3144 (.A1(W3703), .A2(I948), .ZN(O1239));
  NANDX1 G3145 (.A1(I489), .A2(I422), .ZN(W5056));
  NANDX1 G3146 (.A1(W390), .A2(W4549), .ZN(O1242));
  NANDX1 G3147 (.A1(I563), .A2(I830), .ZN(O1243));
  NANDX1 G3148 (.A1(W3964), .A2(W3794), .ZN(O1245));
  NANDX1 G3149 (.A1(I587), .A2(I249), .ZN(W509));
  NANDX1 G3150 (.A1(W3913), .A2(W2464), .ZN(O1246));
  NANDX1 G3151 (.A1(W2669), .A2(W562), .ZN(O1248));
  NANDX1 G3152 (.A1(W414), .A2(I921), .ZN(W507));
  NANDX1 G3153 (.A1(I510), .A2(W4659), .ZN(W4996));
  NANDX1 G3154 (.A1(W281), .A2(I966), .ZN(W544));
  NANDX1 G3155 (.A1(I28), .A2(W26), .ZN(W543));
  NANDX1 G3156 (.A1(I283), .A2(W3877), .ZN(W4972));
  NANDX1 G3157 (.A1(W4047), .A2(W3028), .ZN(O1187));
  NANDX1 G3158 (.A1(W2932), .A2(W4135), .ZN(W4978));
  NANDX1 G3159 (.A1(W2659), .A2(W1144), .ZN(O1190));
  NANDX1 G3160 (.A1(W2127), .A2(W4965), .ZN(O1194));
  NANDX1 G3161 (.A1(I410), .A2(I770), .ZN(W4984));
  NANDX1 G3162 (.A1(I488), .A2(W161), .ZN(W536));
  NANDX1 G3163 (.A1(W1669), .A2(W3570), .ZN(O1197));
  NANDX1 G3164 (.A1(W1), .A2(W387), .ZN(W533));
  NANDX1 G3165 (.A1(W4695), .A2(W4682), .ZN(W5074));
  NANDX1 G3166 (.A1(W2775), .A2(W3056), .ZN(W4997));
  NANDX1 G3167 (.A1(I44), .A2(I983), .ZN(W532));
  NANDX1 G3168 (.A1(W1652), .A2(W3262), .ZN(W5000));
  NANDX1 G3169 (.A1(W440), .A2(W184), .ZN(W531));
  NANDX1 G3170 (.A1(W4559), .A2(W1335), .ZN(W5004));
  NANDX1 G3171 (.A1(I693), .A2(I258), .ZN(W530));
  NANDX1 G3172 (.A1(I735), .A2(W443), .ZN(W529));
  NANDX1 G3173 (.A1(W3590), .A2(W169), .ZN(O1207));
  NANDX1 G3174 (.A1(W2057), .A2(I499), .ZN(O1208));
  NANDX1 G3175 (.A1(I535), .A2(W392), .ZN(W526));
  NANDX1 G3176 (.A1(W4915), .A2(W3019), .ZN(O1213));
  NANDX1 G3177 (.A1(W932), .A2(W556), .ZN(O1306));
  NANDX1 G3178 (.A1(W4441), .A2(W451), .ZN(W5121));
  NANDX1 G3179 (.A1(W2222), .A2(W5047), .ZN(W5124));
  NANDX1 G3180 (.A1(I972), .A2(I973), .ZN(W486));
  NANDX1 G3181 (.A1(I797), .A2(W3164), .ZN(O1289));
  NANDX1 G3182 (.A1(I748), .A2(W35), .ZN(O1294));
  NANDX1 G3183 (.A1(I966), .A2(I967), .ZN(W483));
  NANDX1 G3184 (.A1(I964), .A2(I965), .ZN(W482));
  NANDX1 G3185 (.A1(W2058), .A2(W3271), .ZN(W5140));
  NANDX1 G3186 (.A1(I962), .A2(I963), .ZN(W481));
  NANDX1 G3187 (.A1(W392), .A2(I990), .ZN(O1298));
  NANDX1 G3188 (.A1(W1192), .A2(W2562), .ZN(O1301));
  NANDX1 G3189 (.A1(I115), .A2(W3898), .ZN(O1285));
  NANDX1 G3190 (.A1(I952), .A2(I953), .ZN(W476));
  NANDX1 G3191 (.A1(I946), .A2(I947), .ZN(W473));
  NANDX1 G3192 (.A1(W3233), .A2(W529), .ZN(O1312));
  NANDX1 G3193 (.A1(I944), .A2(I945), .ZN(W472));
  NANDX1 G3194 (.A1(W2385), .A2(W3653), .ZN(W5164));
  NANDX1 G3195 (.A1(W98), .A2(W4482), .ZN(O1316));
  NANDX1 G3196 (.A1(I940), .A2(I941), .ZN(W470));
  NANDX1 G3197 (.A1(I938), .A2(I939), .ZN(W469));
  NANDX1 G3198 (.A1(I932), .A2(I933), .ZN(W466));
  NANDX1 G3199 (.A1(W4355), .A2(W201), .ZN(O1326));
  NANDX1 G3200 (.A1(W4491), .A2(I485), .ZN(W5185));
  NANDX1 G3201 (.A1(W4646), .A2(W4195), .ZN(O1272));
  NANDX1 G3202 (.A1(I85), .A2(I204), .ZN(W503));
  NANDX1 G3203 (.A1(I956), .A2(W255), .ZN(W502));
  NANDX1 G3204 (.A1(W597), .A2(W3569), .ZN(O1254));
  NANDX1 G3205 (.A1(W3061), .A2(W4235), .ZN(O1257));
  NANDX1 G3206 (.A1(W2542), .A2(W4558), .ZN(W5087));
  NANDX1 G3207 (.A1(W2396), .A2(W3263), .ZN(W5088));
  NANDX1 G3208 (.A1(W389), .A2(W3442), .ZN(W5093));
  NANDX1 G3209 (.A1(I994), .A2(I995), .ZN(W497));
  NANDX1 G3210 (.A1(W2034), .A2(I797), .ZN(O1266));
  NANDX1 G3211 (.A1(I992), .A2(I993), .ZN(W496));
  NANDX1 G3212 (.A1(I206), .A2(W775), .ZN(O1268));
  NANDX1 G3213 (.A1(W527), .A2(W117), .ZN(W545));
  NANDX1 G3214 (.A1(I986), .A2(I987), .ZN(W493));
  NANDX1 G3215 (.A1(W2113), .A2(W1872), .ZN(O1275));
  NANDX1 G3216 (.A1(W4067), .A2(W3068), .ZN(O1276));
  NANDX1 G3217 (.A1(I464), .A2(W4744), .ZN(O1277));
  NANDX1 G3218 (.A1(W5088), .A2(W1265), .ZN(W5111));
  NANDX1 G3219 (.A1(W2029), .A2(W1476), .ZN(W5113));
  NANDX1 G3220 (.A1(I980), .A2(I981), .ZN(W490));
  NANDX1 G3221 (.A1(W3242), .A2(W1153), .ZN(O1281));
  NANDX1 G3222 (.A1(W4396), .A2(W3318), .ZN(O1282));
  NANDX1 G3223 (.A1(I976), .A2(I977), .ZN(W488));
  NANDX1 G3224 (.A1(W2782), .A2(W2507), .ZN(W4828));
  NANDX1 G3225 (.A1(W1892), .A2(I340), .ZN(W4811));
  NANDX1 G3226 (.A1(W245), .A2(W2755), .ZN(O1089));
  NANDX1 G3227 (.A1(I774), .A2(W218), .ZN(W589));
  NANDX1 G3228 (.A1(W1240), .A2(W1411), .ZN(O1091));
  NANDX1 G3229 (.A1(I206), .A2(W3947), .ZN(W4816));
  NANDX1 G3230 (.A1(W3816), .A2(W4191), .ZN(O1093));
  NANDX1 G3231 (.A1(W4630), .A2(W3273), .ZN(O1094));
  NANDX1 G3232 (.A1(W328), .A2(W115), .ZN(W588));
  NANDX1 G3233 (.A1(I11), .A2(W4298), .ZN(O1097));
  NANDX1 G3234 (.A1(W39), .A2(W360), .ZN(W587));
  NANDX1 G3235 (.A1(I393), .A2(W2591), .ZN(W4826));
  NANDX1 G3236 (.A1(W872), .A2(W4582), .ZN(O1088));
  NANDX1 G3237 (.A1(W418), .A2(W2528), .ZN(O1101));
  NANDX1 G3238 (.A1(W136), .A2(I932), .ZN(W584));
  NANDX1 G3239 (.A1(W2716), .A2(W473), .ZN(O1103));
  NANDX1 G3240 (.A1(W2003), .A2(W3320), .ZN(W4839));
  NANDX1 G3241 (.A1(W1992), .A2(W4009), .ZN(O1111));
  NANDX1 G3242 (.A1(W1210), .A2(I7), .ZN(O1112));
  NANDX1 G3243 (.A1(W4648), .A2(W1858), .ZN(W4849));
  NANDX1 G3244 (.A1(I175), .A2(I536), .ZN(W579));
  NANDX1 G3245 (.A1(I608), .A2(I179), .ZN(W4855));
  NANDX1 G3246 (.A1(I72), .A2(I384), .ZN(W576));
  NANDX1 G3247 (.A1(W4754), .A2(W2952), .ZN(W4864));
  NANDX1 G3248 (.A1(W1453), .A2(W2178), .ZN(O1074));
  NANDX1 G3249 (.A1(W2220), .A2(W3232), .ZN(W4754));
  NANDX1 G3250 (.A1(I962), .A2(I249), .ZN(O19));
  NANDX1 G3251 (.A1(I447), .A2(W4227), .ZN(O1053));
  NANDX1 G3252 (.A1(I798), .A2(W406), .ZN(W611));
  NANDX1 G3253 (.A1(I180), .A2(W4084), .ZN(O1058));
  NANDX1 G3254 (.A1(W347), .A2(I365), .ZN(W608));
  NANDX1 G3255 (.A1(W627), .A2(W2983), .ZN(O1060));
  NANDX1 G3256 (.A1(W457), .A2(W348), .ZN(W603));
  NANDX1 G3257 (.A1(W102), .A2(W4671), .ZN(O1064));
  NANDX1 G3258 (.A1(W195), .A2(W307), .ZN(W598));
  NANDX1 G3259 (.A1(W1968), .A2(W3979), .ZN(O1073));
  NANDX1 G3260 (.A1(W371), .A2(W2464), .ZN(O1123));
  NANDX1 G3261 (.A1(I731), .A2(W3796), .ZN(O1075));
  NANDX1 G3262 (.A1(W1468), .A2(W3039), .ZN(O1076));
  NANDX1 G3263 (.A1(W2447), .A2(W689), .ZN(O1077));
  NANDX1 G3264 (.A1(I323), .A2(I234), .ZN(W595));
  NANDX1 G3265 (.A1(W2454), .A2(W3976), .ZN(O1079));
  NANDX1 G3266 (.A1(W850), .A2(W1007), .ZN(O1081));
  NANDX1 G3267 (.A1(W2965), .A2(W1249), .ZN(W4797));
  NANDX1 G3268 (.A1(W714), .A2(W3529), .ZN(W4798));
  NANDX1 G3269 (.A1(W272), .A2(I790), .ZN(W594));
  NANDX1 G3270 (.A1(W105), .A2(W494), .ZN(W592));
  NANDX1 G3271 (.A1(W4176), .A2(I58), .ZN(O1087));
  NANDX1 G3272 (.A1(W1897), .A2(I829), .ZN(W4937));
  NANDX1 G3273 (.A1(I416), .A2(W1577), .ZN(W4922));
  NANDX1 G3274 (.A1(W84), .A2(W484), .ZN(W556));
  NANDX1 G3275 (.A1(W1394), .A2(W1887), .ZN(W4924));
  NANDX1 G3276 (.A1(W4824), .A2(I7), .ZN(O1157));
  NANDX1 G3277 (.A1(W57), .A2(W1235), .ZN(O1158));
  NANDX1 G3278 (.A1(W3509), .A2(W2227), .ZN(W4927));
  NANDX1 G3279 (.A1(W2614), .A2(W1421), .ZN(W4928));
  NANDX1 G3280 (.A1(I56), .A2(I70), .ZN(W555));
  NANDX1 G3281 (.A1(W186), .A2(I256), .ZN(W554));
  NANDX1 G3282 (.A1(I26), .A2(I197), .ZN(W553));
  NANDX1 G3283 (.A1(W3875), .A2(W3574), .ZN(O1164));
  NANDX1 G3284 (.A1(I598), .A2(W3526), .ZN(O1155));
  NANDX1 G3285 (.A1(W474), .A2(W510), .ZN(W551));
  NANDX1 G3286 (.A1(W4142), .A2(W77), .ZN(W4940));
  NANDX1 G3287 (.A1(W4497), .A2(W2842), .ZN(O1167));
  NANDX1 G3288 (.A1(I364), .A2(I431), .ZN(O1171));
  NANDX1 G3289 (.A1(W4099), .A2(W3035), .ZN(W4949));
  NANDX1 G3290 (.A1(W1386), .A2(W4014), .ZN(O1174));
  NANDX1 G3291 (.A1(I521), .A2(W1430), .ZN(O1178));
  NANDX1 G3292 (.A1(W4001), .A2(W3578), .ZN(O1179));
  NANDX1 G3293 (.A1(W4826), .A2(W115), .ZN(O1182));
  NANDX1 G3294 (.A1(I198), .A2(W988), .ZN(W4965));
  NANDX1 G3295 (.A1(W3420), .A2(W3471), .ZN(O1183));
  NANDX1 G3296 (.A1(W4397), .A2(W2439), .ZN(O1139));
  NANDX1 G3297 (.A1(W1714), .A2(W4535), .ZN(W4871));
  NANDX1 G3298 (.A1(W3390), .A2(W2133), .ZN(W4872));
  NANDX1 G3299 (.A1(W3216), .A2(W2233), .ZN(O1126));
  NANDX1 G3300 (.A1(I263), .A2(W2541), .ZN(W4878));
  NANDX1 G3301 (.A1(I296), .A2(W2875), .ZN(O1130));
  NANDX1 G3302 (.A1(W445), .A2(W25), .ZN(W568));
  NANDX1 G3303 (.A1(I392), .A2(I677), .ZN(O1134));
  NANDX1 G3304 (.A1(W2267), .A2(W2941), .ZN(O1136));
  NANDX1 G3305 (.A1(I188), .A2(W1279), .ZN(W4891));
  NANDX1 G3306 (.A1(W680), .A2(W2972), .ZN(O1137));
  NANDX1 G3307 (.A1(W1865), .A2(W3263), .ZN(W4893));
  NANDX1 G3308 (.A1(I926), .A2(I927), .ZN(W463));
  NANDX1 G3309 (.A1(W1960), .A2(W1407), .ZN(O1140));
  NANDX1 G3310 (.A1(W216), .A2(W693), .ZN(O1143));
  NANDX1 G3311 (.A1(W196), .A2(I349), .ZN(W564));
  NANDX1 G3312 (.A1(W465), .A2(W2772), .ZN(O1145));
  NANDX1 G3313 (.A1(W4855), .A2(W321), .ZN(W4906));
  NANDX1 G3314 (.A1(I233), .A2(I10), .ZN(W560));
  NANDX1 G3315 (.A1(I858), .A2(W206), .ZN(W559));
  NANDX1 G3316 (.A1(I344), .A2(W185), .ZN(W557));
  NANDX1 G3317 (.A1(I743), .A2(W1313), .ZN(O1153));
  NANDX1 G3318 (.A1(W301), .A2(W2551), .ZN(O1154));
  NANDX1 G3319 (.A1(W515), .A2(W4353), .ZN(O1548));
  NANDX1 G3320 (.A1(W5011), .A2(W954), .ZN(O1532));
  NANDX1 G3321 (.A1(W3927), .A2(W3245), .ZN(O1533));
  NANDX1 G3322 (.A1(I170), .A2(W563), .ZN(O1536));
  NANDX1 G3323 (.A1(W2062), .A2(W3425), .ZN(W5471));
  NANDX1 G3324 (.A1(I614), .A2(W845), .ZN(O1539));
  NANDX1 G3325 (.A1(W1410), .A2(W1973), .ZN(O1542));
  NANDX1 G3326 (.A1(W258), .A2(I992), .ZN(O1543));
  NANDX1 G3327 (.A1(W3839), .A2(I626), .ZN(O1544));
  NANDX1 G3328 (.A1(W2712), .A2(W2730), .ZN(O1545));
  NANDX1 G3329 (.A1(W4359), .A2(W90), .ZN(W5484));
  NANDX1 G3330 (.A1(I720), .A2(I721), .ZN(W360));
  NANDX1 G3331 (.A1(W2674), .A2(W1091), .ZN(O1531));
  NANDX1 G3332 (.A1(W3371), .A2(I164), .ZN(W5487));
  NANDX1 G3333 (.A1(W1073), .A2(W4336), .ZN(O1551));
  NANDX1 G3334 (.A1(I718), .A2(I719), .ZN(W359));
  NANDX1 G3335 (.A1(W3318), .A2(I782), .ZN(W5492));
  NANDX1 G3336 (.A1(W3820), .A2(W79), .ZN(W5493));
  NANDX1 G3337 (.A1(W733), .A2(W1063), .ZN(O1553));
  NANDX1 G3338 (.A1(I714), .A2(I715), .ZN(W357));
  NANDX1 G3339 (.A1(I503), .A2(W5118), .ZN(O1559));
  NANDX1 G3340 (.A1(W3231), .A2(W1179), .ZN(O1561));
  NANDX1 G3341 (.A1(W4297), .A2(W747), .ZN(W5506));
  NANDX1 G3342 (.A1(I704), .A2(I705), .ZN(W352));
  NANDX1 G3343 (.A1(W2925), .A2(W747), .ZN(O1513));
  NANDX1 G3344 (.A1(W4535), .A2(W2821), .ZN(O1490));
  NANDX1 G3345 (.A1(W4604), .A2(I317), .ZN(O1493));
  NANDX1 G3346 (.A1(I772), .A2(I773), .ZN(W386));
  NANDX1 G3347 (.A1(I770), .A2(I771), .ZN(W385));
  NANDX1 G3348 (.A1(W1242), .A2(W3867), .ZN(O1501));
  NANDX1 G3349 (.A1(W449), .A2(W3481), .ZN(O1504));
  NANDX1 G3350 (.A1(W3639), .A2(W1294), .ZN(W5424));
  NANDX1 G3351 (.A1(W2408), .A2(I169), .ZN(W5425));
  NANDX1 G3352 (.A1(I479), .A2(W4865), .ZN(O1505));
  NANDX1 G3353 (.A1(W370), .A2(I426), .ZN(O1507));
  NANDX1 G3354 (.A1(W3090), .A2(W273), .ZN(O1510));
  NANDX1 G3355 (.A1(W4713), .A2(W2129), .ZN(O1566));
  NANDX1 G3356 (.A1(W693), .A2(I660), .ZN(W5438));
  NANDX1 G3357 (.A1(I758), .A2(I759), .ZN(W379));
  NANDX1 G3358 (.A1(I754), .A2(I755), .ZN(W377));
  NANDX1 G3359 (.A1(W2168), .A2(W2926), .ZN(O1517));
  NANDX1 G3360 (.A1(W745), .A2(W817), .ZN(W5448));
  NANDX1 G3361 (.A1(W5435), .A2(W4723), .ZN(O1523));
  NANDX1 G3362 (.A1(I746), .A2(I747), .ZN(W373));
  NANDX1 G3363 (.A1(W4330), .A2(W722), .ZN(O1525));
  NANDX1 G3364 (.A1(I742), .A2(I743), .ZN(W371));
  NANDX1 G3365 (.A1(I740), .A2(I741), .ZN(W370));
  NANDX1 G3366 (.A1(I734), .A2(I735), .ZN(O6));
  NANDX1 G3367 (.A1(W1323), .A2(W4221), .ZN(W5595));
  NANDX1 G3368 (.A1(W2704), .A2(W4171), .ZN(O1612));
  NANDX1 G3369 (.A1(I656), .A2(I657), .ZN(W328));
  NANDX1 G3370 (.A1(W321), .A2(W2992), .ZN(W5576));
  NANDX1 G3371 (.A1(W1915), .A2(W2843), .ZN(W5577));
  NANDX1 G3372 (.A1(W1284), .A2(W1926), .ZN(O1617));
  NANDX1 G3373 (.A1(I654), .A2(I655), .ZN(W327));
  NANDX1 G3374 (.A1(W3980), .A2(W5005), .ZN(O1619));
  NANDX1 G3375 (.A1(W3716), .A2(I267), .ZN(W5587));
  NANDX1 G3376 (.A1(I642), .A2(I643), .ZN(W321));
  NANDX1 G3377 (.A1(I430), .A2(W5436), .ZN(W5591));
  NANDX1 G3378 (.A1(W4798), .A2(W3388), .ZN(O1628));
  NANDX1 G3379 (.A1(I660), .A2(I661), .ZN(W330));
  NANDX1 G3380 (.A1(W4333), .A2(W48), .ZN(O1631));
  NANDX1 G3381 (.A1(W879), .A2(W2412), .ZN(O1632));
  NANDX1 G3382 (.A1(W196), .A2(W2544), .ZN(O1633));
  NANDX1 G3383 (.A1(W663), .A2(W736), .ZN(O1636));
  NANDX1 G3384 (.A1(W952), .A2(W5148), .ZN(O1637));
  NANDX1 G3385 (.A1(W522), .A2(W1288), .ZN(O1644));
  NANDX1 G3386 (.A1(W4940), .A2(W1041), .ZN(W5613));
  NANDX1 G3387 (.A1(W148), .A2(W3510), .ZN(O1649));
  NANDX1 G3388 (.A1(I622), .A2(I623), .ZN(W311));
  NANDX1 G3389 (.A1(W3225), .A2(W725), .ZN(O1652));
  NANDX1 G3390 (.A1(W2465), .A2(W2959), .ZN(O1654));
  NANDX1 G3391 (.A1(W3229), .A2(W3533), .ZN(O1582));
  NANDX1 G3392 (.A1(I696), .A2(I697), .ZN(W348));
  NANDX1 G3393 (.A1(I692), .A2(I693), .ZN(W346));
  NANDX1 G3394 (.A1(I690), .A2(I691), .ZN(W345));
  NANDX1 G3395 (.A1(W463), .A2(W2872), .ZN(O1575));
  NANDX1 G3396 (.A1(W3554), .A2(I817), .ZN(W5525));
  NANDX1 G3397 (.A1(W2284), .A2(W985), .ZN(O1577));
  NANDX1 G3398 (.A1(I854), .A2(W2169), .ZN(W5527));
  NANDX1 G3399 (.A1(I686), .A2(I687), .ZN(W343));
  NANDX1 G3400 (.A1(I351), .A2(W1472), .ZN(O1579));
  NANDX1 G3401 (.A1(I684), .A2(I685), .ZN(W342));
  NANDX1 G3402 (.A1(W1906), .A2(W1104), .ZN(O1581));
  NANDX1 G3403 (.A1(W4879), .A2(I758), .ZN(O1485));
  NANDX1 G3404 (.A1(W4024), .A2(I552), .ZN(O1590));
  NANDX1 G3405 (.A1(W1412), .A2(W1210), .ZN(W5546));
  NANDX1 G3406 (.A1(W2387), .A2(W3691), .ZN(O1594));
  NANDX1 G3407 (.A1(I320), .A2(W1239), .ZN(O1595));
  NANDX1 G3408 (.A1(W4743), .A2(W5221), .ZN(O1596));
  NANDX1 G3409 (.A1(W5), .A2(W3351), .ZN(O1598));
  NANDX1 G3410 (.A1(W1053), .A2(W1113), .ZN(W5558));
  NANDX1 G3411 (.A1(W4839), .A2(W2238), .ZN(O1604));
  NANDX1 G3412 (.A1(W5067), .A2(W2931), .ZN(O1608));
  NANDX1 G3413 (.A1(I664), .A2(I665), .ZN(W332));
  NANDX1 G3414 (.A1(W4986), .A2(W3255), .ZN(O1376));
  NANDX1 G3415 (.A1(W3844), .A2(W5164), .ZN(W5233));
  NANDX1 G3416 (.A1(W1398), .A2(W4651), .ZN(O1358));
  NANDX1 G3417 (.A1(I892), .A2(I893), .ZN(O10));
  NANDX1 G3418 (.A1(W1933), .A2(W2697), .ZN(W5239));
  NANDX1 G3419 (.A1(W833), .A2(W4098), .ZN(O1366));
  NANDX1 G3420 (.A1(W498), .A2(W822), .ZN(O1369));
  NANDX1 G3421 (.A1(W4653), .A2(W4690), .ZN(O1370));
  NANDX1 G3422 (.A1(W566), .A2(W447), .ZN(O1371));
  NANDX1 G3423 (.A1(I886), .A2(I887), .ZN(W443));
  NANDX1 G3424 (.A1(W1699), .A2(W63), .ZN(O1372));
  NANDX1 G3425 (.A1(W9), .A2(W5025), .ZN(W5253));
  NANDX1 G3426 (.A1(W488), .A2(W2159), .ZN(W5232));
  NANDX1 G3427 (.A1(W4787), .A2(W2090), .ZN(O1377));
  NANDX1 G3428 (.A1(W2887), .A2(W3020), .ZN(O1378));
  NANDX1 G3429 (.A1(W3551), .A2(W471), .ZN(O1379));
  NANDX1 G3430 (.A1(I878), .A2(I879), .ZN(W439));
  NANDX1 G3431 (.A1(I135), .A2(W2611), .ZN(O1381));
  NANDX1 G3432 (.A1(W112), .A2(W2937), .ZN(O1382));
  NANDX1 G3433 (.A1(I876), .A2(I877), .ZN(W438));
  NANDX1 G3434 (.A1(W624), .A2(W1977), .ZN(O1385));
  NANDX1 G3435 (.A1(I798), .A2(W4486), .ZN(W5267));
  NANDX1 G3436 (.A1(I872), .A2(I873), .ZN(W436));
  NANDX1 G3437 (.A1(W388), .A2(W4111), .ZN(W5273));
  NANDX1 G3438 (.A1(W1992), .A2(W3320), .ZN(W5213));
  NANDX1 G3439 (.A1(I810), .A2(W4732), .ZN(O1328));
  NANDX1 G3440 (.A1(W2829), .A2(W4293), .ZN(W5191));
  NANDX1 G3441 (.A1(I920), .A2(I921), .ZN(W460));
  NANDX1 G3442 (.A1(I264), .A2(W404), .ZN(O1332));
  NANDX1 G3443 (.A1(I918), .A2(I919), .ZN(O13));
  NANDX1 G3444 (.A1(W2942), .A2(W4684), .ZN(O1334));
  NANDX1 G3445 (.A1(W1624), .A2(W2940), .ZN(W5199));
  NANDX1 G3446 (.A1(I906), .A2(I907), .ZN(W453));
  NANDX1 G3447 (.A1(I904), .A2(I905), .ZN(W452));
  NANDX1 G3448 (.A1(I755), .A2(I113), .ZN(W5210));
  NANDX1 G3449 (.A1(W1544), .A2(I147), .ZN(W5211));
  NANDX1 G3450 (.A1(W2367), .A2(W4371), .ZN(O1393));
  NANDX1 G3451 (.A1(W3898), .A2(W1369), .ZN(O1346));
  NANDX1 G3452 (.A1(I902), .A2(I903), .ZN(W451));
  NANDX1 G3453 (.A1(I900), .A2(I901), .ZN(W450));
  NANDX1 G3454 (.A1(W2251), .A2(W2003), .ZN(W5221));
  NANDX1 G3455 (.A1(W115), .A2(I606), .ZN(W5222));
  NANDX1 G3456 (.A1(W2210), .A2(W3224), .ZN(O1351));
  NANDX1 G3457 (.A1(I730), .A2(W415), .ZN(W5225));
  NANDX1 G3458 (.A1(W4827), .A2(W4501), .ZN(O1352));
  NANDX1 G3459 (.A1(W1642), .A2(W3098), .ZN(O1353));
  NANDX1 G3460 (.A1(W2955), .A2(W1153), .ZN(W5228));
  NANDX1 G3461 (.A1(W4856), .A2(W1740), .ZN(O1356));
  NANDX1 G3462 (.A1(W5183), .A2(W2909), .ZN(O1460));
  NANDX1 G3463 (.A1(I820), .A2(I821), .ZN(W410));
  NANDX1 G3464 (.A1(W4343), .A2(W5228), .ZN(W5338));
  NANDX1 G3465 (.A1(W3722), .A2(W1390), .ZN(O1437));
  NANDX1 G3466 (.A1(I428), .A2(W4893), .ZN(O1438));
  NANDX1 G3467 (.A1(W3218), .A2(W3526), .ZN(O1443));
  NANDX1 G3468 (.A1(W5168), .A2(W4880), .ZN(O1444));
  NANDX1 G3469 (.A1(I812), .A2(I813), .ZN(W406));
  NANDX1 G3470 (.A1(I810), .A2(I811), .ZN(W405));
  NANDX1 G3471 (.A1(W5215), .A2(W675), .ZN(O1450));
  NANDX1 G3472 (.A1(W4505), .A2(W223), .ZN(O1452));
  NANDX1 G3473 (.A1(W3391), .A2(W5101), .ZN(W5362));
  NANDX1 G3474 (.A1(I826), .A2(I827), .ZN(W413));
  NANDX1 G3475 (.A1(I798), .A2(I799), .ZN(W399));
  NANDX1 G3476 (.A1(W584), .A2(W4331), .ZN(O1462));
  NANDX1 G3477 (.A1(I796), .A2(I797), .ZN(W398));
  NANDX1 G3478 (.A1(W202), .A2(W897), .ZN(O1467));
  NANDX1 G3479 (.A1(W4282), .A2(I158), .ZN(W5381));
  NANDX1 G3480 (.A1(W4689), .A2(W3479), .ZN(O1471));
  NANDX1 G3481 (.A1(W4748), .A2(W4938), .ZN(O1474));
  NANDX1 G3482 (.A1(W2635), .A2(W342), .ZN(O1479));
  NANDX1 G3483 (.A1(W4707), .A2(W1093), .ZN(O1480));
  NANDX1 G3484 (.A1(W4302), .A2(W2559), .ZN(O1482));
  NANDX1 G3485 (.A1(W791), .A2(W4633), .ZN(W5396));
  NANDX1 G3486 (.A1(W123), .A2(W1190), .ZN(O1414));
  NANDX1 G3487 (.A1(W879), .A2(W5030), .ZN(O1395));
  NANDX1 G3488 (.A1(I152), .A2(W378), .ZN(W5288));
  NANDX1 G3489 (.A1(W3201), .A2(W4094), .ZN(O1403));
  NANDX1 G3490 (.A1(I848), .A2(I849), .ZN(W424));
  NANDX1 G3491 (.A1(W121), .A2(W4035), .ZN(O1405));
  NANDX1 G3492 (.A1(I661), .A2(W1789), .ZN(W5298));
  NANDX1 G3493 (.A1(W918), .A2(I843), .ZN(W5300));
  NANDX1 G3494 (.A1(I842), .A2(I843), .ZN(W421));
  NANDX1 G3495 (.A1(I409), .A2(I728), .ZN(W5307));
  NANDX1 G3496 (.A1(W3798), .A2(W2747), .ZN(O1411));
  NANDX1 G3497 (.A1(W2017), .A2(W3957), .ZN(O1413));
  NANDX1 G3498 (.A1(W351), .A2(I245), .ZN(W616));
  NANDX1 G3499 (.A1(I85), .A2(W3279), .ZN(O1417));
  NANDX1 G3500 (.A1(W5028), .A2(W784), .ZN(O1418));
  NANDX1 G3501 (.A1(W2417), .A2(W3738), .ZN(O1419));
  NANDX1 G3502 (.A1(W2178), .A2(I956), .ZN(O1420));
  NANDX1 G3503 (.A1(W4247), .A2(I17), .ZN(O1425));
  NANDX1 G3504 (.A1(W3038), .A2(W2039), .ZN(W5325));
  NANDX1 G3505 (.A1(I828), .A2(I829), .ZN(W414));
  NANDX1 G3506 (.A1(W1016), .A2(W2556), .ZN(O1429));
  NANDX1 G3507 (.A1(W1295), .A2(W2588), .ZN(O1430));
  NANDX1 G3508 (.A1(I750), .A2(W668), .ZN(W5331));
  NANDX1 G3509 (.A1(W1072), .A2(W157), .ZN(W2611));
  NANDX1 G3510 (.A1(I355), .A2(I646), .ZN(O240));
  NANDX1 G3511 (.A1(I148), .A2(I454), .ZN(W1317));
  NANDX1 G3512 (.A1(W408), .A2(W801), .ZN(W1315));
  NANDX1 G3513 (.A1(W1882), .A2(W2911), .ZN(W3508));
  NANDX1 G3514 (.A1(W1566), .A2(W436), .ZN(W2597));
  NANDX1 G3515 (.A1(W2192), .A2(W2112), .ZN(O243));
  NANDX1 G3516 (.A1(W299), .A2(W2361), .ZN(W2602));
  NANDX1 G3517 (.A1(W2112), .A2(I217), .ZN(W2603));
  NANDX1 G3518 (.A1(W1776), .A2(W386), .ZN(W2606));
  NANDX1 G3519 (.A1(W180), .A2(W1623), .ZN(W2607));
  NANDX1 G3520 (.A1(I975), .A2(W2140), .ZN(W2586));
  NANDX1 G3521 (.A1(W2379), .A2(W2456), .ZN(W2612));
  NANDX1 G3522 (.A1(I52), .A2(I122), .ZN(W2613));
  NANDX1 G3523 (.A1(I781), .A2(W2396), .ZN(W2614));
  NANDX1 G3524 (.A1(W1898), .A2(W1832), .ZN(W2616));
  NANDX1 G3525 (.A1(W420), .A2(W265), .ZN(W2619));
  NANDX1 G3526 (.A1(W1291), .A2(W740), .ZN(W2623));
  NANDX1 G3527 (.A1(W863), .A2(W288), .ZN(W1310));
  NANDX1 G3528 (.A1(I793), .A2(W735), .ZN(W2631));
  NANDX1 G3529 (.A1(W1256), .A2(W895), .ZN(W2634));
  NANDX1 G3530 (.A1(W1277), .A2(I259), .ZN(W2563));
  NANDX1 G3531 (.A1(W2462), .A2(W662), .ZN(W2545));
  NANDX1 G3532 (.A1(I296), .A2(W1044), .ZN(W2549));
  NANDX1 G3533 (.A1(W1267), .A2(W2530), .ZN(W2552));
  NANDX1 G3534 (.A1(I437), .A2(W1446), .ZN(O234));
  NANDX1 G3535 (.A1(W2074), .A2(W1804), .ZN(O235));
  NANDX1 G3536 (.A1(W1456), .A2(I664), .ZN(W2557));
  NANDX1 G3537 (.A1(W875), .A2(W1540), .ZN(W2559));
  NANDX1 G3538 (.A1(W2489), .A2(W887), .ZN(O236));
  NANDX1 G3539 (.A1(I818), .A2(I284), .ZN(W2561));
  NANDX1 G3540 (.A1(W687), .A2(I405), .ZN(W1327));
  NANDX1 G3541 (.A1(I944), .A2(W1695), .ZN(W2637));
  NANDX1 G3542 (.A1(W1814), .A2(I222), .ZN(W2565));
  NANDX1 G3543 (.A1(W1211), .A2(W653), .ZN(W1326));
  NANDX1 G3544 (.A1(W1341), .A2(W1493), .ZN(O237));
  NANDX1 G3545 (.A1(W410), .A2(W1097), .ZN(W1323));
  NANDX1 G3546 (.A1(I57), .A2(W921), .ZN(W1322));
  NANDX1 G3547 (.A1(I90), .A2(I49), .ZN(W1321));
  NANDX1 G3548 (.A1(W1814), .A2(W948), .ZN(W2576));
  NANDX1 G3549 (.A1(W1544), .A2(W1810), .ZN(W2580));
  NANDX1 G3550 (.A1(W532), .A2(W2412), .ZN(O238));
  NANDX1 G3551 (.A1(I688), .A2(I391), .ZN(O269));
  NANDX1 G3552 (.A1(W1756), .A2(I948), .ZN(O262));
  NANDX1 G3553 (.A1(W573), .A2(W1271), .ZN(W2683));
  NANDX1 G3554 (.A1(W1198), .A2(W41), .ZN(W1287));
  NANDX1 G3555 (.A1(I704), .A2(W1456), .ZN(W2688));
  NANDX1 G3556 (.A1(W211), .A2(W1115), .ZN(W2690));
  NANDX1 G3557 (.A1(I719), .A2(W2441), .ZN(W2695));
  NANDX1 G3558 (.A1(I668), .A2(W1276), .ZN(W2699));
  NANDX1 G3559 (.A1(W841), .A2(W450), .ZN(W2700));
  NANDX1 G3560 (.A1(W1005), .A2(W2069), .ZN(W2701));
  NANDX1 G3561 (.A1(W83), .A2(W1659), .ZN(W2706));
  NANDX1 G3562 (.A1(I594), .A2(W2442), .ZN(O261));
  NANDX1 G3563 (.A1(W531), .A2(W1797), .ZN(W2709));
  NANDX1 G3564 (.A1(I455), .A2(W590), .ZN(W1282));
  NANDX1 G3565 (.A1(I958), .A2(W1714), .ZN(O270));
  NANDX1 G3566 (.A1(W2298), .A2(W1211), .ZN(W2717));
  NANDX1 G3567 (.A1(W707), .A2(W2139), .ZN(W2719));
  NANDX1 G3568 (.A1(W292), .A2(W775), .ZN(W1278));
  NANDX1 G3569 (.A1(I794), .A2(W691), .ZN(W2722));
  NANDX1 G3570 (.A1(W803), .A2(W899), .ZN(W2726));
  NANDX1 G3571 (.A1(I920), .A2(W597), .ZN(W1277));
  NANDX1 G3572 (.A1(I223), .A2(I442), .ZN(W1294));
  NANDX1 G3573 (.A1(W2611), .A2(W1353), .ZN(W2638));
  NANDX1 G3574 (.A1(W1258), .A2(W2442), .ZN(W2639));
  NANDX1 G3575 (.A1(W2117), .A2(I317), .ZN(W2643));
  NANDX1 G3576 (.A1(W2284), .A2(W1912), .ZN(W2648));
  NANDX1 G3577 (.A1(W1271), .A2(W1693), .ZN(W2651));
  NANDX1 G3578 (.A1(W298), .A2(W1686), .ZN(O254));
  NANDX1 G3579 (.A1(W1221), .A2(I702), .ZN(W1297));
  NANDX1 G3580 (.A1(I170), .A2(I890), .ZN(W1295));
  NANDX1 G3581 (.A1(W1134), .A2(I798), .ZN(O256));
  NANDX1 G3582 (.A1(W2037), .A2(I894), .ZN(W2544));
  NANDX1 G3583 (.A1(I337), .A2(W560), .ZN(W2664));
  NANDX1 G3584 (.A1(W143), .A2(I388), .ZN(W2666));
  NANDX1 G3585 (.A1(W2396), .A2(W1681), .ZN(W2668));
  NANDX1 G3586 (.A1(W308), .A2(W2635), .ZN(W2669));
  NANDX1 G3587 (.A1(I154), .A2(I152), .ZN(W2671));
  NANDX1 G3588 (.A1(W991), .A2(W888), .ZN(W1293));
  NANDX1 G3589 (.A1(I174), .A2(I170), .ZN(W2676));
  NANDX1 G3590 (.A1(W479), .A2(W2565), .ZN(W2677));
  NANDX1 G3591 (.A1(W997), .A2(W2243), .ZN(O260));
  NANDX1 G3592 (.A1(W868), .A2(W682), .ZN(W2453));
  NANDX1 G3593 (.A1(W2223), .A2(W2122), .ZN(W2426));
  NANDX1 G3594 (.A1(W1497), .A2(W29), .ZN(O210));
  NANDX1 G3595 (.A1(W2162), .A2(W1424), .ZN(O211));
  NANDX1 G3596 (.A1(W1820), .A2(W1075), .ZN(O213));
  NANDX1 G3597 (.A1(W604), .A2(W2210), .ZN(W2443));
  NANDX1 G3598 (.A1(W1097), .A2(W984), .ZN(W1362));
  NANDX1 G3599 (.A1(I896), .A2(I887), .ZN(W1360));
  NANDX1 G3600 (.A1(W1565), .A2(W1554), .ZN(W2449));
  NANDX1 G3601 (.A1(W90), .A2(W87), .ZN(W2451));
  NANDX1 G3602 (.A1(W403), .A2(W433), .ZN(W1358));
  NANDX1 G3603 (.A1(W716), .A2(W230), .ZN(W2423));
  NANDX1 G3604 (.A1(W1513), .A2(W1456), .ZN(W2454));
  NANDX1 G3605 (.A1(W628), .A2(W630), .ZN(W1357));
  NANDX1 G3606 (.A1(W519), .A2(W2083), .ZN(W2457));
  NANDX1 G3607 (.A1(W2341), .A2(W2380), .ZN(W2458));
  NANDX1 G3608 (.A1(I269), .A2(W1036), .ZN(W2459));
  NANDX1 G3609 (.A1(W685), .A2(W930), .ZN(W2460));
  NANDX1 G3610 (.A1(I822), .A2(W704), .ZN(W2461));
  NANDX1 G3611 (.A1(W799), .A2(W2282), .ZN(W2462));
  NANDX1 G3612 (.A1(W968), .A2(W342), .ZN(W1355));
  NANDX1 G3613 (.A1(W1009), .A2(W1401), .ZN(W2397));
  NANDX1 G3614 (.A1(W2261), .A2(W1502), .ZN(O203));
  NANDX1 G3615 (.A1(W276), .A2(W497), .ZN(W2386));
  NANDX1 G3616 (.A1(W2282), .A2(I375), .ZN(W2387));
  NANDX1 G3617 (.A1(I56), .A2(W1964), .ZN(W2389));
  NANDX1 G3618 (.A1(W310), .A2(W336), .ZN(W2391));
  NANDX1 G3619 (.A1(W492), .A2(I637), .ZN(W2392));
  NANDX1 G3620 (.A1(W776), .A2(I301), .ZN(W1380));
  NANDX1 G3621 (.A1(W564), .A2(I495), .ZN(W1378));
  NANDX1 G3622 (.A1(W438), .A2(I696), .ZN(W1377));
  NANDX1 G3623 (.A1(W1353), .A2(I192), .ZN(W1354));
  NANDX1 G3624 (.A1(W1639), .A2(I213), .ZN(W2398));
  NANDX1 G3625 (.A1(W29), .A2(W924), .ZN(W1376));
  NANDX1 G3626 (.A1(W1048), .A2(W738), .ZN(W2401));
  NANDX1 G3627 (.A1(I92), .A2(W537), .ZN(W1373));
  NANDX1 G3628 (.A1(W272), .A2(W2255), .ZN(O205));
  NANDX1 G3629 (.A1(W1667), .A2(I80), .ZN(W2412));
  NANDX1 G3630 (.A1(W400), .A2(W762), .ZN(W1370));
  NANDX1 G3631 (.A1(W2340), .A2(W1918), .ZN(W2421));
  NANDX1 G3632 (.A1(W783), .A2(W341), .ZN(W2422));
  NANDX1 G3633 (.A1(W1046), .A2(W2436), .ZN(W2526));
  NANDX1 G3634 (.A1(W2249), .A2(I480), .ZN(W2505));
  NANDX1 G3635 (.A1(I618), .A2(I975), .ZN(W1341));
  NANDX1 G3636 (.A1(W1994), .A2(W2411), .ZN(W2507));
  NANDX1 G3637 (.A1(W495), .A2(W767), .ZN(W1340));
  NANDX1 G3638 (.A1(I787), .A2(W1524), .ZN(W2509));
  NANDX1 G3639 (.A1(W2407), .A2(I542), .ZN(W2511));
  NANDX1 G3640 (.A1(W1125), .A2(I518), .ZN(W2516));
  NANDX1 G3641 (.A1(W2113), .A2(W1762), .ZN(W2522));
  NANDX1 G3642 (.A1(W770), .A2(W2400), .ZN(W2523));
  NANDX1 G3643 (.A1(W1404), .A2(W1462), .ZN(O226));
  NANDX1 G3644 (.A1(W1258), .A2(W950), .ZN(W2504));
  NANDX1 G3645 (.A1(I888), .A2(W2127), .ZN(W2528));
  NANDX1 G3646 (.A1(I86), .A2(W664), .ZN(W2531));
  NANDX1 G3647 (.A1(W1835), .A2(W1812), .ZN(O228));
  NANDX1 G3648 (.A1(W917), .A2(W1048), .ZN(O63));
  NANDX1 G3649 (.A1(I668), .A2(W134), .ZN(W2537));
  NANDX1 G3650 (.A1(W1344), .A2(W228), .ZN(W2539));
  NANDX1 G3651 (.A1(I50), .A2(W2124), .ZN(W2540));
  NANDX1 G3652 (.A1(I50), .A2(W2308), .ZN(W2542));
  NANDX1 G3653 (.A1(W1824), .A2(W1682), .ZN(O229));
  NANDX1 G3654 (.A1(I752), .A2(W1288), .ZN(W2488));
  NANDX1 G3655 (.A1(W663), .A2(I552), .ZN(W1353));
  NANDX1 G3656 (.A1(W1348), .A2(I538), .ZN(W2471));
  NANDX1 G3657 (.A1(I746), .A2(W716), .ZN(W2472));
  NANDX1 G3658 (.A1(W829), .A2(W1913), .ZN(W2473));
  NANDX1 G3659 (.A1(W2350), .A2(W1526), .ZN(W2477));
  NANDX1 G3660 (.A1(W209), .A2(W1201), .ZN(W1351));
  NANDX1 G3661 (.A1(W546), .A2(W845), .ZN(W2482));
  NANDX1 G3662 (.A1(I154), .A2(I302), .ZN(W1349));
  NANDX1 G3663 (.A1(W1274), .A2(I9), .ZN(W2487));
  NANDX1 G3664 (.A1(I132), .A2(I225), .ZN(W1276));
  NANDX1 G3665 (.A1(I386), .A2(W629), .ZN(W2489));
  NANDX1 G3666 (.A1(I43), .A2(W1196), .ZN(W1348));
  NANDX1 G3667 (.A1(W745), .A2(W428), .ZN(W1347));
  NANDX1 G3668 (.A1(W2365), .A2(W1416), .ZN(O219));
  NANDX1 G3669 (.A1(W370), .A2(W764), .ZN(W1346));
  NANDX1 G3670 (.A1(W817), .A2(I946), .ZN(W2497));
  NANDX1 G3671 (.A1(W439), .A2(W279), .ZN(W1344));
  NANDX1 G3672 (.A1(W275), .A2(W794), .ZN(W1343));
  NANDX1 G3673 (.A1(I62), .A2(I284), .ZN(W2503));
  NANDX1 G3674 (.A1(W2362), .A2(W183), .ZN(W2997));
  NANDX1 G3675 (.A1(W2050), .A2(W1572), .ZN(W2971));
  NANDX1 G3676 (.A1(W2452), .A2(W2150), .ZN(O337));
  NANDX1 G3677 (.A1(W423), .A2(I696), .ZN(W1196));
  NANDX1 G3678 (.A1(W2874), .A2(W353), .ZN(W2976));
  NANDX1 G3679 (.A1(W56), .A2(W679), .ZN(W2980));
  NANDX1 G3680 (.A1(W2308), .A2(W281), .ZN(W2983));
  NANDX1 G3681 (.A1(I375), .A2(W72), .ZN(W2984));
  NANDX1 G3682 (.A1(W644), .A2(I962), .ZN(O340));
  NANDX1 G3683 (.A1(I804), .A2(W1748), .ZN(W2993));
  NANDX1 G3684 (.A1(W1959), .A2(W2481), .ZN(W2994));
  NANDX1 G3685 (.A1(W272), .A2(W91), .ZN(O53));
  NANDX1 G3686 (.A1(W1718), .A2(W406), .ZN(W2999));
  NANDX1 G3687 (.A1(W334), .A2(W975), .ZN(W3001));
  NANDX1 G3688 (.A1(W1105), .A2(W118), .ZN(O51));
  NANDX1 G3689 (.A1(I100), .A2(I113), .ZN(W3005));
  NANDX1 G3690 (.A1(W24), .A2(W2731), .ZN(O343));
  NANDX1 G3691 (.A1(W619), .A2(W132), .ZN(W1187));
  NANDX1 G3692 (.A1(W619), .A2(W497), .ZN(W3009));
  NANDX1 G3693 (.A1(I314), .A2(W2057), .ZN(W3011));
  NANDX1 G3694 (.A1(W59), .A2(I753), .ZN(O345));
  NANDX1 G3695 (.A1(W770), .A2(W2110), .ZN(W2951));
  NANDX1 G3696 (.A1(W1614), .A2(W207), .ZN(W2926));
  NANDX1 G3697 (.A1(W2866), .A2(W2641), .ZN(O328));
  NANDX1 G3698 (.A1(I572), .A2(I767), .ZN(W2931));
  NANDX1 G3699 (.A1(I964), .A2(I766), .ZN(W2932));
  NANDX1 G3700 (.A1(W1318), .A2(W371), .ZN(W2941));
  NANDX1 G3701 (.A1(W979), .A2(W708), .ZN(W1208));
  NANDX1 G3702 (.A1(I560), .A2(I64), .ZN(O332));
  NANDX1 G3703 (.A1(W1058), .A2(W709), .ZN(W1205));
  NANDX1 G3704 (.A1(W498), .A2(I356), .ZN(W1203));
  NANDX1 G3705 (.A1(I600), .A2(I297), .ZN(W3016));
  NANDX1 G3706 (.A1(I212), .A2(W502), .ZN(W1201));
  NANDX1 G3707 (.A1(W585), .A2(W2172), .ZN(W2958));
  NANDX1 G3708 (.A1(W2389), .A2(W1476), .ZN(W2959));
  NANDX1 G3709 (.A1(I564), .A2(I974), .ZN(W1200));
  NANDX1 G3710 (.A1(I588), .A2(W468), .ZN(W1199));
  NANDX1 G3711 (.A1(W1276), .A2(I684), .ZN(W2964));
  NANDX1 G3712 (.A1(W2082), .A2(W2884), .ZN(W2965));
  NANDX1 G3713 (.A1(W418), .A2(I346), .ZN(W2968));
  NANDX1 G3714 (.A1(I227), .A2(W427), .ZN(W1198));
  NANDX1 G3715 (.A1(W2149), .A2(W150), .ZN(O360));
  NANDX1 G3716 (.A1(W151), .A2(W2793), .ZN(O356));
  NANDX1 G3717 (.A1(I271), .A2(I843), .ZN(W1161));
  NANDX1 G3718 (.A1(W1010), .A2(W125), .ZN(W3069));
  NANDX1 G3719 (.A1(I196), .A2(W2668), .ZN(O357));
  NANDX1 G3720 (.A1(I431), .A2(W2127), .ZN(O358));
  NANDX1 G3721 (.A1(W867), .A2(W2800), .ZN(W3074));
  NANDX1 G3722 (.A1(I978), .A2(W540), .ZN(W3076));
  NANDX1 G3723 (.A1(I264), .A2(W821), .ZN(W1158));
  NANDX1 G3724 (.A1(I312), .A2(W2801), .ZN(W3080));
  NANDX1 G3725 (.A1(I5), .A2(I2), .ZN(W1157));
  NANDX1 G3726 (.A1(I555), .A2(I676), .ZN(W1164));
  NANDX1 G3727 (.A1(W386), .A2(I482), .ZN(W1156));
  NANDX1 G3728 (.A1(W1018), .A2(W1464), .ZN(W3087));
  NANDX1 G3729 (.A1(I800), .A2(I191), .ZN(W1155));
  NANDX1 G3730 (.A1(W437), .A2(W779), .ZN(O362));
  NANDX1 G3731 (.A1(W1749), .A2(W1440), .ZN(W3092));
  NANDX1 G3732 (.A1(W2268), .A2(W482), .ZN(O364));
  NANDX1 G3733 (.A1(W658), .A2(W266), .ZN(W1152));
  NANDX1 G3734 (.A1(W1048), .A2(I253), .ZN(W1150));
  NANDX1 G3735 (.A1(W2791), .A2(I61), .ZN(O368));
  NANDX1 G3736 (.A1(W2196), .A2(W2786), .ZN(O350));
  NANDX1 G3737 (.A1(I735), .A2(I446), .ZN(W1183));
  NANDX1 G3738 (.A1(I581), .A2(I776), .ZN(W1179));
  NANDX1 G3739 (.A1(I58), .A2(W627), .ZN(W3023));
  NANDX1 G3740 (.A1(W2916), .A2(W2819), .ZN(W3025));
  NANDX1 G3741 (.A1(W1320), .A2(W2747), .ZN(W3028));
  NANDX1 G3742 (.A1(I929), .A2(I148), .ZN(W1175));
  NANDX1 G3743 (.A1(I81), .A2(W2646), .ZN(W3031));
  NANDX1 G3744 (.A1(I598), .A2(W52), .ZN(W1174));
  NANDX1 G3745 (.A1(W1754), .A2(W1975), .ZN(W3039));
  NANDX1 G3746 (.A1(W1597), .A2(I924), .ZN(W2923));
  NANDX1 G3747 (.A1(W2629), .A2(W449), .ZN(W3042));
  NANDX1 G3748 (.A1(W597), .A2(W2189), .ZN(W3045));
  NANDX1 G3749 (.A1(W386), .A2(W436), .ZN(W1169));
  NANDX1 G3750 (.A1(I820), .A2(W2085), .ZN(W3049));
  NANDX1 G3751 (.A1(W1702), .A2(W974), .ZN(W3050));
  NANDX1 G3752 (.A1(W1134), .A2(W741), .ZN(W1167));
  NANDX1 G3753 (.A1(W2457), .A2(W878), .ZN(W3055));
  NANDX1 G3754 (.A1(W807), .A2(W1146), .ZN(W3060));
  NANDX1 G3755 (.A1(I543), .A2(W1004), .ZN(W1165));
  NANDX1 G3756 (.A1(W1177), .A2(W201), .ZN(W2806));
  NANDX1 G3757 (.A1(W693), .A2(W638), .ZN(W1258));
  NANDX1 G3758 (.A1(I457), .A2(I2), .ZN(W2791));
  NANDX1 G3759 (.A1(W345), .A2(I237), .ZN(W2792));
  NANDX1 G3760 (.A1(W1573), .A2(W379), .ZN(W2794));
  NANDX1 G3761 (.A1(I862), .A2(W547), .ZN(W2796));
  NANDX1 G3762 (.A1(I480), .A2(W1966), .ZN(W2797));
  NANDX1 G3763 (.A1(W1918), .A2(I538), .ZN(W2800));
  NANDX1 G3764 (.A1(I510), .A2(W1076), .ZN(W2802));
  NANDX1 G3765 (.A1(W2393), .A2(I582), .ZN(W2803));
  NANDX1 G3766 (.A1(I683), .A2(W338), .ZN(W1254));
  NANDX1 G3767 (.A1(W1564), .A2(I55), .ZN(O288));
  NANDX1 G3768 (.A1(I332), .A2(W60), .ZN(W1252));
  NANDX1 G3769 (.A1(W996), .A2(I126), .ZN(W2808));
  NANDX1 G3770 (.A1(W907), .A2(W1225), .ZN(W1248));
  NANDX1 G3771 (.A1(I511), .A2(W2374), .ZN(W2814));
  NANDX1 G3772 (.A1(I12), .A2(I336), .ZN(W1245));
  NANDX1 G3773 (.A1(W1632), .A2(I121), .ZN(W2819));
  NANDX1 G3774 (.A1(W600), .A2(I967), .ZN(W1244));
  NANDX1 G3775 (.A1(W771), .A2(W1080), .ZN(O296));
  NANDX1 G3776 (.A1(I993), .A2(W1975), .ZN(W2823));
  NANDX1 G3777 (.A1(W254), .A2(W829), .ZN(W1266));
  NANDX1 G3778 (.A1(W1736), .A2(I722), .ZN(W2733));
  NANDX1 G3779 (.A1(W1190), .A2(W2059), .ZN(W2735));
  NANDX1 G3780 (.A1(I656), .A2(W1088), .ZN(W1272));
  NANDX1 G3781 (.A1(W405), .A2(I945), .ZN(W2740));
  NANDX1 G3782 (.A1(W1053), .A2(I137), .ZN(O276));
  NANDX1 G3783 (.A1(W1274), .A2(W2160), .ZN(W2747));
  NANDX1 G3784 (.A1(W256), .A2(I65), .ZN(W1268));
  NANDX1 G3785 (.A1(W1717), .A2(W2200), .ZN(W2752));
  NANDX1 G3786 (.A1(W234), .A2(W895), .ZN(W2753));
  NANDX1 G3787 (.A1(I539), .A2(W1454), .ZN(W2825));
  NANDX1 G3788 (.A1(W778), .A2(I531), .ZN(W1264));
  NANDX1 G3789 (.A1(I166), .A2(W1934), .ZN(O282));
  NANDX1 G3790 (.A1(W2349), .A2(I560), .ZN(W2764));
  NANDX1 G3791 (.A1(W970), .A2(I439), .ZN(W1263));
  NANDX1 G3792 (.A1(W760), .A2(W415), .ZN(W1262));
  NANDX1 G3793 (.A1(W1143), .A2(I310), .ZN(W2770));
  NANDX1 G3794 (.A1(I831), .A2(W704), .ZN(W1260));
  NANDX1 G3795 (.A1(W2279), .A2(W2321), .ZN(O285));
  NANDX1 G3796 (.A1(I718), .A2(W1518), .ZN(W2786));
  NANDX1 G3797 (.A1(W1997), .A2(W2320), .ZN(O320));
  NANDX1 G3798 (.A1(I19), .A2(I987), .ZN(O55));
  NANDX1 G3799 (.A1(W875), .A2(W1800), .ZN(O312));
  NANDX1 G3800 (.A1(W2024), .A2(W405), .ZN(O313));
  NANDX1 G3801 (.A1(W1993), .A2(W1242), .ZN(O314));
  NANDX1 G3802 (.A1(W2000), .A2(I94), .ZN(W2884));
  NANDX1 G3803 (.A1(I226), .A2(W656), .ZN(O317));
  NANDX1 G3804 (.A1(W578), .A2(I511), .ZN(W2887));
  NANDX1 G3805 (.A1(W2530), .A2(W1902), .ZN(W2892));
  NANDX1 G3806 (.A1(W1038), .A2(W1565), .ZN(W2893));
  NANDX1 G3807 (.A1(I74), .A2(I463), .ZN(W2894));
  NANDX1 G3808 (.A1(W1054), .A2(W741), .ZN(W1231));
  NANDX1 G3809 (.A1(I374), .A2(I21), .ZN(W1221));
  NANDX1 G3810 (.A1(W156), .A2(W571), .ZN(W1220));
  NANDX1 G3811 (.A1(W405), .A2(W1605), .ZN(W2901));
  NANDX1 G3812 (.A1(W1910), .A2(I20), .ZN(W2902));
  NANDX1 G3813 (.A1(I50), .A2(I598), .ZN(W1216));
  NANDX1 G3814 (.A1(W2862), .A2(W629), .ZN(W2913));
  NANDX1 G3815 (.A1(W2726), .A2(W1827), .ZN(O323));
  NANDX1 G3816 (.A1(I832), .A2(W18), .ZN(W2921));
  NANDX1 G3817 (.A1(I490), .A2(I738), .ZN(O326));
  NANDX1 G3818 (.A1(W590), .A2(W6), .ZN(O306));
  NANDX1 G3819 (.A1(W1027), .A2(I452), .ZN(O299));
  NANDX1 G3820 (.A1(W887), .A2(W1387), .ZN(O300));
  NANDX1 G3821 (.A1(W2116), .A2(W1393), .ZN(W2831));
  NANDX1 G3822 (.A1(W1406), .A2(W365), .ZN(W2833));
  NANDX1 G3823 (.A1(I554), .A2(I401), .ZN(W1241));
  NANDX1 G3824 (.A1(I302), .A2(W1408), .ZN(W2841));
  NANDX1 G3825 (.A1(W2251), .A2(W86), .ZN(W2842));
  NANDX1 G3826 (.A1(I4), .A2(I498), .ZN(W2844));
  NANDX1 G3827 (.A1(W2249), .A2(W2062), .ZN(O303));
  NANDX1 G3828 (.A1(I551), .A2(W1124), .ZN(W2383));
  NANDX1 G3829 (.A1(I531), .A2(W1077), .ZN(O307));
  NANDX1 G3830 (.A1(W2746), .A2(W2591), .ZN(W2860));
  NANDX1 G3831 (.A1(W334), .A2(W3), .ZN(O310));
  NANDX1 G3832 (.A1(W770), .A2(I203), .ZN(W1232));
  NANDX1 G3833 (.A1(W2216), .A2(W666), .ZN(W2865));
  NANDX1 G3834 (.A1(W70), .A2(W1307), .ZN(W2866));
  NANDX1 G3835 (.A1(W2028), .A2(W1607), .ZN(W2867));
  NANDX1 G3836 (.A1(W800), .A2(I305), .ZN(W2869));
  NANDX1 G3837 (.A1(W128), .A2(W910), .ZN(O311));
  NANDX1 G3838 (.A1(I726), .A2(W837), .ZN(W1540));
  NANDX1 G3839 (.A1(I998), .A2(W1398), .ZN(O119));
  NANDX1 G3840 (.A1(W1855), .A2(W1861), .ZN(W1879));
  NANDX1 G3841 (.A1(W1295), .A2(W869), .ZN(W1880));
  NANDX1 G3842 (.A1(W388), .A2(W783), .ZN(W1550));
  NANDX1 G3843 (.A1(W1505), .A2(I147), .ZN(W1885));
  NANDX1 G3844 (.A1(I842), .A2(W224), .ZN(W1548));
  NANDX1 G3845 (.A1(W436), .A2(W1171), .ZN(W1891));
  NANDX1 G3846 (.A1(I798), .A2(W314), .ZN(W1541));
  NANDX1 G3847 (.A1(W1390), .A2(W553), .ZN(W1904));
  NANDX1 G3848 (.A1(W122), .A2(W1483), .ZN(W1905));
  NANDX1 G3849 (.A1(W1062), .A2(W1064), .ZN(W1875));
  NANDX1 G3850 (.A1(W111), .A2(W1027), .ZN(O124));
  NANDX1 G3851 (.A1(W1651), .A2(W854), .ZN(W1911));
  NANDX1 G3852 (.A1(W1711), .A2(W1203), .ZN(W1913));
  NANDX1 G3853 (.A1(W1856), .A2(W1520), .ZN(W1914));
  NANDX1 G3854 (.A1(I794), .A2(W348), .ZN(W1917));
  NANDX1 G3855 (.A1(W1299), .A2(I834), .ZN(W1918));
  NANDX1 G3856 (.A1(W1037), .A2(W1023), .ZN(O127));
  NANDX1 G3857 (.A1(W80), .A2(I268), .ZN(W1924));
  NANDX1 G3858 (.A1(W412), .A2(W983), .ZN(W1926));
  NANDX1 G3859 (.A1(I192), .A2(I408), .ZN(W1557));
  NANDX1 G3860 (.A1(W532), .A2(W1801), .ZN(O115));
  NANDX1 G3861 (.A1(W695), .A2(W1408), .ZN(W1833));
  NANDX1 G3862 (.A1(I195), .A2(W1647), .ZN(W1836));
  NANDX1 G3863 (.A1(W1190), .A2(W1056), .ZN(W1837));
  NANDX1 G3864 (.A1(I75), .A2(I330), .ZN(W1839));
  NANDX1 G3865 (.A1(W1605), .A2(I66), .ZN(W1840));
  NANDX1 G3866 (.A1(I202), .A2(W148), .ZN(W1564));
  NANDX1 G3867 (.A1(W203), .A2(W1142), .ZN(W1560));
  NANDX1 G3868 (.A1(W468), .A2(I613), .ZN(W1847));
  NANDX1 G3869 (.A1(W42), .A2(I620), .ZN(W1559));
  NANDX1 G3870 (.A1(W1585), .A2(I412), .ZN(W1929));
  NANDX1 G3871 (.A1(W898), .A2(W172), .ZN(W1855));
  NANDX1 G3872 (.A1(I52), .A2(W828), .ZN(W1857));
  NANDX1 G3873 (.A1(W1067), .A2(W860), .ZN(W1858));
  NANDX1 G3874 (.A1(W1821), .A2(W266), .ZN(W1861));
  NANDX1 G3875 (.A1(I526), .A2(I878), .ZN(W1863));
  NANDX1 G3876 (.A1(I974), .A2(W580), .ZN(W1553));
  NANDX1 G3877 (.A1(W1804), .A2(I297), .ZN(W1870));
  NANDX1 G3878 (.A1(W1344), .A2(W1361), .ZN(W1872));
  NANDX1 G3879 (.A1(W403), .A2(W398), .ZN(W1552));
  NANDX1 G3880 (.A1(W281), .A2(W321), .ZN(W1982));
  NANDX1 G3881 (.A1(W827), .A2(W926), .ZN(O75));
  NANDX1 G3882 (.A1(I537), .A2(W278), .ZN(O131));
  NANDX1 G3883 (.A1(I285), .A2(I940), .ZN(O74));
  NANDX1 G3884 (.A1(W1902), .A2(W1040), .ZN(O132));
  NANDX1 G3885 (.A1(W34), .A2(W1416), .ZN(W1520));
  NANDX1 G3886 (.A1(W1352), .A2(W462), .ZN(W1971));
  NANDX1 G3887 (.A1(I827), .A2(I3), .ZN(W1973));
  NANDX1 G3888 (.A1(W1326), .A2(W1355), .ZN(W1977));
  NANDX1 G3889 (.A1(W400), .A2(I702), .ZN(W1978));
  NANDX1 G3890 (.A1(W1482), .A2(W1341), .ZN(W1981));
  NANDX1 G3891 (.A1(W277), .A2(W1573), .ZN(W1962));
  NANDX1 G3892 (.A1(W1237), .A2(W849), .ZN(W1985));
  NANDX1 G3893 (.A1(I180), .A2(W665), .ZN(W1986));
  NANDX1 G3894 (.A1(W1681), .A2(W247), .ZN(W1994));
  NANDX1 G3895 (.A1(I312), .A2(W1915), .ZN(W1995));
  NANDX1 G3896 (.A1(W213), .A2(I457), .ZN(W1997));
  NANDX1 G3897 (.A1(W268), .A2(I542), .ZN(W1998));
  NANDX1 G3898 (.A1(W346), .A2(W1277), .ZN(W2001));
  NANDX1 G3899 (.A1(W1700), .A2(W344), .ZN(W2005));
  NANDX1 G3900 (.A1(W470), .A2(I215), .ZN(W1506));
  NANDX1 G3901 (.A1(W122), .A2(I791), .ZN(W1528));
  NANDX1 G3902 (.A1(I214), .A2(I440), .ZN(W1930));
  NANDX1 G3903 (.A1(I12), .A2(I350), .ZN(O79));
  NANDX1 G3904 (.A1(I348), .A2(I192), .ZN(W1934));
  NANDX1 G3905 (.A1(W816), .A2(I315), .ZN(W1935));
  NANDX1 G3906 (.A1(W538), .A2(W1919), .ZN(W1936));
  NANDX1 G3907 (.A1(W147), .A2(I94), .ZN(W1937));
  NANDX1 G3908 (.A1(I541), .A2(W337), .ZN(W1940));
  NANDX1 G3909 (.A1(I306), .A2(W1398), .ZN(O77));
  NANDX1 G3910 (.A1(W521), .A2(W1150), .ZN(W1946));
  NANDX1 G3911 (.A1(W1807), .A2(W996), .ZN(W1830));
  NANDX1 G3912 (.A1(I348), .A2(I347), .ZN(W1948));
  NANDX1 G3913 (.A1(W380), .A2(I601), .ZN(W1527));
  NANDX1 G3914 (.A1(W642), .A2(W358), .ZN(W1526));
  NANDX1 G3915 (.A1(I737), .A2(W393), .ZN(W1952));
  NANDX1 G3916 (.A1(I436), .A2(W314), .ZN(W1524));
  NANDX1 G3917 (.A1(I687), .A2(I128), .ZN(W1957));
  NANDX1 G3918 (.A1(I786), .A2(I255), .ZN(O129));
  NANDX1 G3919 (.A1(W1320), .A2(W1644), .ZN(W1960));
  NANDX1 G3920 (.A1(I207), .A2(W327), .ZN(O130));
  NANDX1 G3921 (.A1(W40), .A2(W1314), .ZN(W1700));
  NANDX1 G3922 (.A1(W845), .A2(I695), .ZN(W1681));
  NANDX1 G3923 (.A1(I306), .A2(I162), .ZN(W1683));
  NANDX1 G3924 (.A1(W1085), .A2(W408), .ZN(O93));
  NANDX1 G3925 (.A1(W1209), .A2(W1143), .ZN(W1686));
  NANDX1 G3926 (.A1(W38), .A2(W319), .ZN(O94));
  NANDX1 G3927 (.A1(W238), .A2(W409), .ZN(W1688));
  NANDX1 G3928 (.A1(I910), .A2(I317), .ZN(W1690));
  NANDX1 G3929 (.A1(W207), .A2(W770), .ZN(W1694));
  NANDX1 G3930 (.A1(W1406), .A2(W987), .ZN(W1696));
  NANDX1 G3931 (.A1(W9), .A2(W312), .ZN(W1616));
  NANDX1 G3932 (.A1(W1409), .A2(I673), .ZN(W1624));
  NANDX1 G3933 (.A1(W27), .A2(W203), .ZN(W1704));
  NANDX1 G3934 (.A1(W652), .A2(W1171), .ZN(O86));
  NANDX1 G3935 (.A1(W1191), .A2(I692), .ZN(W1713));
  NANDX1 G3936 (.A1(W1575), .A2(W642), .ZN(W1718));
  NANDX1 G3937 (.A1(I621), .A2(I941), .ZN(W1605));
  NANDX1 G3938 (.A1(I656), .A2(W1689), .ZN(W1723));
  NANDX1 G3939 (.A1(W906), .A2(W185), .ZN(W1730));
  NANDX1 G3940 (.A1(W570), .A2(W540), .ZN(W1732));
  NANDX1 G3941 (.A1(W1373), .A2(W711), .ZN(W1733));
  NANDX1 G3942 (.A1(W98), .A2(I832), .ZN(W1663));
  NANDX1 G3943 (.A1(I679), .A2(W689), .ZN(W1637));
  NANDX1 G3944 (.A1(W1405), .A2(W1218), .ZN(O89));
  NANDX1 G3945 (.A1(W795), .A2(W734), .ZN(W1644));
  NANDX1 G3946 (.A1(W595), .A2(I142), .ZN(W1649));
  NANDX1 G3947 (.A1(W87), .A2(W1086), .ZN(W1631));
  NANDX1 G3948 (.A1(W950), .A2(I357), .ZN(W1654));
  NANDX1 G3949 (.A1(W1230), .A2(W621), .ZN(O92));
  NANDX1 G3950 (.A1(W1536), .A2(W1132), .ZN(W1657));
  NANDX1 G3951 (.A1(I890), .A2(I530), .ZN(W1660));
  NANDX1 G3952 (.A1(W1356), .A2(W1675), .ZN(W1736));
  NANDX1 G3953 (.A1(W1629), .A2(W810), .ZN(W1664));
  NANDX1 G3954 (.A1(W377), .A2(W1114), .ZN(W1666));
  NANDX1 G3955 (.A1(W318), .A2(I594), .ZN(W1671));
  NANDX1 G3956 (.A1(I120), .A2(W711), .ZN(W1626));
  NANDX1 G3957 (.A1(W1090), .A2(W929), .ZN(W1675));
  NANDX1 G3958 (.A1(W937), .A2(W1379), .ZN(W1676));
  NANDX1 G3959 (.A1(W1075), .A2(I644), .ZN(W1677));
  NANDX1 G3960 (.A1(W799), .A2(W1388), .ZN(W1678));
  NANDX1 G3961 (.A1(W1441), .A2(W683), .ZN(W1679));
  NANDX1 G3962 (.A1(I259), .A2(W1308), .ZN(W1574));
  NANDX1 G3963 (.A1(W798), .A2(W851), .ZN(W1794));
  NANDX1 G3964 (.A1(I525), .A2(I286), .ZN(W1799));
  NANDX1 G3965 (.A1(W130), .A2(W952), .ZN(W1800));
  NANDX1 G3966 (.A1(W619), .A2(W1120), .ZN(W1577));
  NANDX1 G3967 (.A1(W673), .A2(W1725), .ZN(W1802));
  NANDX1 G3968 (.A1(I394), .A2(W187), .ZN(W1805));
  NANDX1 G3969 (.A1(W1277), .A2(W1070), .ZN(W1807));
  NANDX1 G3970 (.A1(W1474), .A2(W481), .ZN(O110));
  NANDX1 G3971 (.A1(W604), .A2(I885), .ZN(W1575));
  NANDX1 G3972 (.A1(W1277), .A2(I909), .ZN(W1810));
  NANDX1 G3973 (.A1(W180), .A2(W1076), .ZN(W1790));
  NANDX1 G3974 (.A1(I661), .A2(W929), .ZN(W1812));
  NANDX1 G3975 (.A1(W651), .A2(I440), .ZN(W1815));
  NANDX1 G3976 (.A1(I558), .A2(W1368), .ZN(W1816));
  NANDX1 G3977 (.A1(I238), .A2(W116), .ZN(W1817));
  NANDX1 G3978 (.A1(W124), .A2(W1418), .ZN(O112));
  NANDX1 G3979 (.A1(W1651), .A2(I752), .ZN(W1822));
  NANDX1 G3980 (.A1(W1041), .A2(I782), .ZN(W1823));
  NANDX1 G3981 (.A1(I747), .A2(W661), .ZN(W1569));
  NANDX1 G3982 (.A1(W1053), .A2(W288), .ZN(W1568));
  NANDX1 G3983 (.A1(W735), .A2(W516), .ZN(W1584));
  NANDX1 G3984 (.A1(W1734), .A2(W1078), .ZN(W1738));
  NANDX1 G3985 (.A1(I298), .A2(W343), .ZN(O102));
  NANDX1 G3986 (.A1(I437), .A2(I109), .ZN(O83));
  NANDX1 G3987 (.A1(W856), .A2(W1288), .ZN(W1747));
  NANDX1 G3988 (.A1(I368), .A2(W1668), .ZN(W1750));
  NANDX1 G3989 (.A1(W823), .A2(W1298), .ZN(W1751));
  NANDX1 G3990 (.A1(W355), .A2(W1511), .ZN(W1754));
  NANDX1 G3991 (.A1(W159), .A2(I36), .ZN(W1758));
  NANDX1 G3992 (.A1(I880), .A2(I440), .ZN(W1759));
  NANDX1 G3993 (.A1(W1476), .A2(W1185), .ZN(W2008));
  NANDX1 G3994 (.A1(I875), .A2(I528), .ZN(W1768));
  NANDX1 G3995 (.A1(I541), .A2(W168), .ZN(O106));
  NANDX1 G3996 (.A1(W1421), .A2(W785), .ZN(W1772));
  NANDX1 G3997 (.A1(I524), .A2(W110), .ZN(W1773));
  NANDX1 G3998 (.A1(W1216), .A2(I117), .ZN(W1774));
  NANDX1 G3999 (.A1(I636), .A2(I29), .ZN(W1775));
  NANDX1 G4000 (.A1(W498), .A2(I472), .ZN(W1776));
  NANDX1 G4001 (.A1(W406), .A2(W90), .ZN(W1777));
  NANDX1 G4002 (.A1(W188), .A2(I592), .ZN(W1579));
  NANDX1 G4003 (.A1(W442), .A2(W308), .ZN(W2272));
  NANDX1 G4004 (.A1(W1759), .A2(W770), .ZN(O182));
  NANDX1 G4005 (.A1(I631), .A2(W66), .ZN(W2253));
  NANDX1 G4006 (.A1(W259), .A2(I583), .ZN(W1421));
  NANDX1 G4007 (.A1(W431), .A2(W448), .ZN(O184));
  NANDX1 G4008 (.A1(W737), .A2(W1051), .ZN(W1419));
  NANDX1 G4009 (.A1(W1497), .A2(I885), .ZN(W2263));
  NANDX1 G4010 (.A1(W1355), .A2(W541), .ZN(W1417));
  NANDX1 G4011 (.A1(W270), .A2(W264), .ZN(W2267));
  NANDX1 G4012 (.A1(W219), .A2(I197), .ZN(W1415));
  NANDX1 G4013 (.A1(I509), .A2(I413), .ZN(O185));
  NANDX1 G4014 (.A1(W96), .A2(W443), .ZN(W2249));
  NANDX1 G4015 (.A1(I368), .A2(I843), .ZN(W1413));
  NANDX1 G4016 (.A1(W1216), .A2(W55), .ZN(W1412));
  NANDX1 G4017 (.A1(I967), .A2(I463), .ZN(W2280));
  NANDX1 G4018 (.A1(W682), .A2(W231), .ZN(W2284));
  NANDX1 G4019 (.A1(W1769), .A2(W524), .ZN(W2286));
  NANDX1 G4020 (.A1(I934), .A2(W1590), .ZN(O187));
  NANDX1 G4021 (.A1(W1384), .A2(I114), .ZN(W1408));
  NANDX1 G4022 (.A1(I257), .A2(W895), .ZN(W1407));
  NANDX1 G4023 (.A1(I960), .A2(W1624), .ZN(W2294));
  NANDX1 G4024 (.A1(W2135), .A2(I906), .ZN(W2219));
  NANDX1 G4025 (.A1(W891), .A2(W710), .ZN(W1440));
  NANDX1 G4026 (.A1(W391), .A2(W2031), .ZN(W2197));
  NANDX1 G4027 (.A1(W1624), .A2(W961), .ZN(O172));
  NANDX1 G4028 (.A1(W255), .A2(W1430), .ZN(W1435));
  NANDX1 G4029 (.A1(W461), .A2(I785), .ZN(O174));
  NANDX1 G4030 (.A1(W1836), .A2(W1623), .ZN(O176));
  NANDX1 G4031 (.A1(W2172), .A2(W1953), .ZN(W2210));
  NANDX1 G4032 (.A1(W313), .A2(W1548), .ZN(W2211));
  NANDX1 G4033 (.A1(W1766), .A2(I323), .ZN(W2212));
  NANDX1 G4034 (.A1(W1647), .A2(W79), .ZN(W2295));
  NANDX1 G4035 (.A1(W754), .A2(I745), .ZN(W1431));
  NANDX1 G4036 (.A1(W82), .A2(I207), .ZN(O177));
  NANDX1 G4037 (.A1(W1257), .A2(W811), .ZN(W2226));
  NANDX1 G4038 (.A1(W1126), .A2(I742), .ZN(W2230));
  NANDX1 G4039 (.A1(I202), .A2(I216), .ZN(W2240));
  NANDX1 G4040 (.A1(W279), .A2(I643), .ZN(W1425));
  NANDX1 G4041 (.A1(I347), .A2(W887), .ZN(W1423));
  NANDX1 G4042 (.A1(W1812), .A2(I648), .ZN(W2246));
  NANDX1 G4043 (.A1(I168), .A2(W289), .ZN(W2247));
  NANDX1 G4044 (.A1(W432), .A2(W1021), .ZN(W2352));
  NANDX1 G4045 (.A1(W712), .A2(W80), .ZN(W1395));
  NANDX1 G4046 (.A1(W1810), .A2(W154), .ZN(W2336));
  NANDX1 G4047 (.A1(W166), .A2(W257), .ZN(W1393));
  NANDX1 G4048 (.A1(W2151), .A2(W1105), .ZN(W2339));
  NANDX1 G4049 (.A1(W1942), .A2(W1794), .ZN(W2341));
  NANDX1 G4050 (.A1(W896), .A2(W18), .ZN(W2343));
  NANDX1 G4051 (.A1(I821), .A2(W745), .ZN(O197));
  NANDX1 G4052 (.A1(W662), .A2(I123), .ZN(O198));
  NANDX1 G4053 (.A1(W966), .A2(W53), .ZN(W2349));
  NANDX1 G4054 (.A1(W743), .A2(W478), .ZN(W1390));
  NANDX1 G4055 (.A1(W692), .A2(W178), .ZN(W2332));
  NANDX1 G4056 (.A1(W780), .A2(W1990), .ZN(W2356));
  NANDX1 G4057 (.A1(W1075), .A2(W238), .ZN(W1387));
  NANDX1 G4058 (.A1(W4), .A2(W2099), .ZN(W2361));
  NANDX1 G4059 (.A1(I264), .A2(I92), .ZN(W2364));
  NANDX1 G4060 (.A1(I734), .A2(W1227), .ZN(W2369));
  NANDX1 G4061 (.A1(W1465), .A2(I888), .ZN(W2370));
  NANDX1 G4062 (.A1(W2192), .A2(I84), .ZN(O202));
  NANDX1 G4063 (.A1(W2240), .A2(I352), .ZN(W2376));
  NANDX1 G4064 (.A1(W1422), .A2(I169), .ZN(W2382));
  NANDX1 G4065 (.A1(I352), .A2(W1020), .ZN(W2311));
  NANDX1 G4066 (.A1(W115), .A2(W923), .ZN(W2297));
  NANDX1 G4067 (.A1(W1051), .A2(W451), .ZN(W2298));
  NANDX1 G4068 (.A1(W472), .A2(I315), .ZN(W1402));
  NANDX1 G4069 (.A1(W1956), .A2(W1322), .ZN(W2300));
  NANDX1 G4070 (.A1(W1390), .A2(I19), .ZN(W2302));
  NANDX1 G4071 (.A1(W1307), .A2(W1185), .ZN(W2305));
  NANDX1 G4072 (.A1(W1513), .A2(W2030), .ZN(W2306));
  NANDX1 G4073 (.A1(W1201), .A2(W865), .ZN(W2309));
  NANDX1 G4074 (.A1(W1015), .A2(W1017), .ZN(W1399));
  NANDX1 G4075 (.A1(W1008), .A2(W1784), .ZN(W2187));
  NANDX1 G4076 (.A1(W239), .A2(W1931), .ZN(W2312));
  NANDX1 G4077 (.A1(W2181), .A2(I336), .ZN(W2313));
  NANDX1 G4078 (.A1(I274), .A2(W918), .ZN(W2316));
  NANDX1 G4079 (.A1(W2225), .A2(W1456), .ZN(W2318));
  NANDX1 G4080 (.A1(I838), .A2(I5), .ZN(W2320));
  NANDX1 G4081 (.A1(W2060), .A2(W969), .ZN(W2321));
  NANDX1 G4082 (.A1(I691), .A2(W408), .ZN(W2322));
  NANDX1 G4083 (.A1(W281), .A2(W1041), .ZN(W2323));
  NANDX1 G4084 (.A1(I521), .A2(I71), .ZN(O194));
  NANDX1 G4085 (.A1(W347), .A2(W850), .ZN(W2079));
  NANDX1 G4086 (.A1(W104), .A2(W492), .ZN(W1493));
  NANDX1 G4087 (.A1(W965), .A2(W1369), .ZN(W2059));
  NANDX1 G4088 (.A1(W880), .A2(W1163), .ZN(O142));
  NANDX1 G4089 (.A1(W163), .A2(I732), .ZN(W1490));
  NANDX1 G4090 (.A1(W1490), .A2(I877), .ZN(W2065));
  NANDX1 G4091 (.A1(W748), .A2(W528), .ZN(W2066));
  NANDX1 G4092 (.A1(W1959), .A2(I64), .ZN(W2069));
  NANDX1 G4093 (.A1(W671), .A2(I650), .ZN(W2072));
  NANDX1 G4094 (.A1(W1475), .A2(W278), .ZN(W1484));
  NANDX1 G4095 (.A1(I179), .A2(W34), .ZN(W1483));
  NANDX1 G4096 (.A1(I960), .A2(W1865), .ZN(W2053));
  NANDX1 G4097 (.A1(W752), .A2(I300), .ZN(W2081));
  NANDX1 G4098 (.A1(I556), .A2(W1264), .ZN(W2083));
  NANDX1 G4099 (.A1(I925), .A2(W624), .ZN(W1478));
  NANDX1 G4100 (.A1(W1155), .A2(I424), .ZN(W2090));
  NANDX1 G4101 (.A1(W118), .A2(W710), .ZN(O147));
  NANDX1 G4102 (.A1(W1042), .A2(I797), .ZN(W1476));
  NANDX1 G4103 (.A1(W125), .A2(W1659), .ZN(O149));
  NANDX1 G4104 (.A1(W1208), .A2(W110), .ZN(W1475));
  NANDX1 G4105 (.A1(I526), .A2(W570), .ZN(W2098));
  NANDX1 G4106 (.A1(W1460), .A2(W1928), .ZN(W2026));
  NANDX1 G4107 (.A1(W719), .A2(W1431), .ZN(W2011));
  NANDX1 G4108 (.A1(W1118), .A2(W901), .ZN(W2013));
  NANDX1 G4109 (.A1(I346), .A2(W1339), .ZN(O136));
  NANDX1 G4110 (.A1(W432), .A2(W313), .ZN(W2017));
  NANDX1 G4111 (.A1(W482), .A2(W857), .ZN(W2018));
  NANDX1 G4112 (.A1(W1502), .A2(W1674), .ZN(W2019));
  NANDX1 G4113 (.A1(W590), .A2(I941), .ZN(O138));
  NANDX1 G4114 (.A1(W563), .A2(I163), .ZN(W2023));
  NANDX1 G4115 (.A1(I522), .A2(I506), .ZN(W2025));
  NANDX1 G4116 (.A1(W1044), .A2(I657), .ZN(W1473));
  NANDX1 G4117 (.A1(W117), .A2(W612), .ZN(W2030));
  NANDX1 G4118 (.A1(W1249), .A2(W14), .ZN(W2033));
  NANDX1 G4119 (.A1(W1325), .A2(W935), .ZN(W2034));
  NANDX1 G4120 (.A1(I271), .A2(W1240), .ZN(W1502));
  NANDX1 G4121 (.A1(W663), .A2(W765), .ZN(W2042));
  NANDX1 G4122 (.A1(W344), .A2(I536), .ZN(W1500));
  NANDX1 G4123 (.A1(W856), .A2(W584), .ZN(O73));
  NANDX1 G4124 (.A1(W1159), .A2(W1037), .ZN(W2050));
  NANDX1 G4125 (.A1(I231), .A2(I646), .ZN(O141));
  NANDX1 G4126 (.A1(W1880), .A2(W651), .ZN(O165));
  NANDX1 G4127 (.A1(W77), .A2(W1407), .ZN(W2149));
  NANDX1 G4128 (.A1(W374), .A2(W1200), .ZN(W1456));
  NANDX1 G4129 (.A1(W125), .A2(W1763), .ZN(O162));
  NANDX1 G4130 (.A1(I469), .A2(W1080), .ZN(W2153));
  NANDX1 G4131 (.A1(W1797), .A2(I241), .ZN(W2154));
  NANDX1 G4132 (.A1(W580), .A2(W50), .ZN(W1455));
  NANDX1 G4133 (.A1(I318), .A2(I248), .ZN(W1454));
  NANDX1 G4134 (.A1(I152), .A2(W452), .ZN(W1453));
  NANDX1 G4135 (.A1(W994), .A2(W1042), .ZN(W1451));
  NANDX1 G4136 (.A1(W724), .A2(W2035), .ZN(W2163));
  NANDX1 G4137 (.A1(I468), .A2(I980), .ZN(W1457));
  NANDX1 G4138 (.A1(I491), .A2(I916), .ZN(W2167));
  NANDX1 G4139 (.A1(I844), .A2(W249), .ZN(W2170));
  NANDX1 G4140 (.A1(W487), .A2(W304), .ZN(W2171));
  NANDX1 G4141 (.A1(W970), .A2(I550), .ZN(W1446));
  NANDX1 G4142 (.A1(W694), .A2(W310), .ZN(W2174));
  NANDX1 G4143 (.A1(W77), .A2(W1313), .ZN(W2175));
  NANDX1 G4144 (.A1(W1927), .A2(W174), .ZN(W2177));
  NANDX1 G4145 (.A1(W950), .A2(I765), .ZN(W2179));
  NANDX1 G4146 (.A1(W2098), .A2(I857), .ZN(W2181));
  NANDX1 G4147 (.A1(W306), .A2(W1973), .ZN(W2124));
  NANDX1 G4148 (.A1(I3), .A2(W1012), .ZN(W2100));
  NANDX1 G4149 (.A1(W1628), .A2(W1185), .ZN(O154));
  NANDX1 G4150 (.A1(W428), .A2(I65), .ZN(W1472));
  NANDX1 G4151 (.A1(W1174), .A2(I398), .ZN(W1471));
  NANDX1 G4152 (.A1(W49), .A2(W167), .ZN(W1470));
  NANDX1 G4153 (.A1(W545), .A2(W1168), .ZN(W2113));
  NANDX1 G4154 (.A1(I355), .A2(W1463), .ZN(O156));
  NANDX1 G4155 (.A1(W57), .A2(W1634), .ZN(O157));
  NANDX1 G4156 (.A1(I30), .A2(W1213), .ZN(W2119));
  NANDX1 G4157 (.A1(W2394), .A2(I412), .ZN(O242));
  NANDX1 G4158 (.A1(W52), .A2(I266), .ZN(W2129));
  NANDX1 G4159 (.A1(W461), .A2(W245), .ZN(W1466));
  NANDX1 G4160 (.A1(I967), .A2(W216), .ZN(W1465));
  NANDX1 G4161 (.A1(W1054), .A2(W1743), .ZN(W2132));
  NANDX1 G4162 (.A1(I499), .A2(W2026), .ZN(W2134));
  NANDX1 G4163 (.A1(I838), .A2(I788), .ZN(W1463));
  NANDX1 G4164 (.A1(W521), .A2(W396), .ZN(W1461));
  NANDX1 G4165 (.A1(W681), .A2(I457), .ZN(W2142));
  NANDX1 G4166 (.A1(W1020), .A2(W378), .ZN(W2146));
  NANDX1 G4167 (.A1(W2470), .A2(W2556), .ZN(W3333));
  NANDX1 G4168 (.A1(W811), .A2(W1021), .ZN(W3140));
  NANDX1 G4169 (.A1(W2701), .A2(W211), .ZN(W3429));
  NANDX1 G4170 (.A1(W1866), .A2(W889), .ZN(O420));
  NANDX1 G4171 (.A1(W806), .A2(W747), .ZN(W1133));
  NANDX1 G4172 (.A1(W2675), .A2(I782), .ZN(O406));
  NANDX1 G4173 (.A1(W1468), .A2(W2584), .ZN(O398));
  NANDX1 G4174 (.A1(W492), .A2(W143), .ZN(W1054));
  NANDX1 G4175 (.A1(W1595), .A2(W239), .ZN(W3271));
  NANDX1 G4176 (.A1(W2637), .A2(W1788), .ZN(W3230));
  NANDX1 G4177 (.A1(W3159), .A2(W858), .ZN(W3371));
  NANDX1 G4178 (.A1(W559), .A2(W1519), .ZN(W3196));
  NANDX1 G4179 (.A1(W1747), .A2(I734), .ZN(W3370));
  NANDX1 G4180 (.A1(I756), .A2(W58), .ZN(O396));
  NANDX1 G4181 (.A1(W980), .A2(W633), .ZN(O395));
  NANDX1 G4182 (.A1(W1041), .A2(W3293), .ZN(O446));
  NANDX1 G4183 (.A1(I609), .A2(W123), .ZN(W1033));
  NANDX1 G4184 (.A1(I876), .A2(I977), .ZN(W1018));
  NANDX1 G4185 (.A1(W1464), .A2(W1210), .ZN(O380));
  NANDX1 G4186 (.A1(W1219), .A2(W1558), .ZN(W3334));
  NANDX1 G4187 (.A1(W2949), .A2(I673), .ZN(W3148));
  NANDX1 G4188 (.A1(W1175), .A2(W3102), .ZN(W3189));
  NANDX1 G4189 (.A1(W186), .A2(I715), .ZN(W1090));
  NANDX1 G4190 (.A1(W2607), .A2(W1291), .ZN(O462));
  NANDX1 G4191 (.A1(W1978), .A2(W747), .ZN(O482));
  NANDX1 G4192 (.A1(W1094), .A2(I766), .ZN(W1121));
  NANDX1 G4193 (.A1(I872), .A2(W879), .ZN(W1067));
  NANDX1 G4194 (.A1(W259), .A2(I549), .ZN(W1032));
  NANDX1 G4195 (.A1(W148), .A2(I71), .ZN(O442));
  NANDX1 G4196 (.A1(W487), .A2(W657), .ZN(W1051));
  NANDX1 G4197 (.A1(W1863), .A2(W2048), .ZN(W3202));
  NANDX1 G4198 (.A1(W2582), .A2(W1801), .ZN(W3321));
  NANDX1 G4199 (.A1(W2807), .A2(W2793), .ZN(O429));
  NANDX1 G4200 (.A1(I346), .A2(W868), .ZN(W1016));
  NANDX1 G4201 (.A1(W2148), .A2(W2436), .ZN(O484));
  NANDX1 G4202 (.A1(I357), .A2(W1971), .ZN(W3385));
  NANDX1 G4203 (.A1(W2068), .A2(W2189), .ZN(O431));
  NANDX1 G4204 (.A1(W1288), .A2(I460), .ZN(W3384));
  NANDX1 G4205 (.A1(W1835), .A2(W3142), .ZN(O422));
  NANDX1 G4206 (.A1(W2196), .A2(I827), .ZN(O448));
  NANDX1 G4207 (.A1(I656), .A2(W265), .ZN(W1138));
  NANDX1 G4208 (.A1(W63), .A2(W3301), .ZN(W3420));
  NANDX1 G4209 (.A1(W860), .A2(W646), .ZN(W3281));
  NANDX1 G4210 (.A1(W2800), .A2(I991), .ZN(W3280));
  NANDX1 G4211 (.A1(W922), .A2(W1097), .ZN(O481));
  NANDX1 G4212 (.A1(W2541), .A2(W2965), .ZN(O374));
  NANDX1 G4213 (.A1(W706), .A2(I430), .ZN(W1036));
  NANDX1 G4214 (.A1(W3162), .A2(W2444), .ZN(W3328));
  NANDX1 G4215 (.A1(W1649), .A2(W3035), .ZN(W3329));
  NANDX1 G4216 (.A1(I170), .A2(I469), .ZN(O405));
  NANDX1 G4217 (.A1(W2548), .A2(I242), .ZN(O375));
  NANDX1 G4218 (.A1(W2913), .A2(W441), .ZN(W3277));
  NANDX1 G4219 (.A1(W2854), .A2(W2611), .ZN(O483));
  NANDX1 G4220 (.A1(W592), .A2(W1516), .ZN(W3199));
  NANDX1 G4221 (.A1(W1822), .A2(W3148), .ZN(W3377));
  NANDX1 G4222 (.A1(W3001), .A2(W212), .ZN(O457));
  NANDX1 G4223 (.A1(I843), .A2(W3325), .ZN(W3484));
  NANDX1 G4224 (.A1(W1463), .A2(W1860), .ZN(O377));
  NANDX1 G4225 (.A1(I100), .A2(I650), .ZN(W3447));
  NANDX1 G4226 (.A1(W2595), .A2(W3410), .ZN(O476));
  NANDX1 G4227 (.A1(W670), .A2(I620), .ZN(W3359));
  NANDX1 G4228 (.A1(W2363), .A2(W1655), .ZN(O475));
  NANDX1 G4229 (.A1(W1812), .A2(W1834), .ZN(O474));
  NANDX1 G4230 (.A1(W1857), .A2(W2640), .ZN(W3444));
  NANDX1 G4231 (.A1(W457), .A2(I38), .ZN(O44));
  NANDX1 G4232 (.A1(W1107), .A2(W3027), .ZN(O411));
  NANDX1 G4233 (.A1(I326), .A2(W2415), .ZN(W3358));
  NANDX1 G4234 (.A1(W1990), .A2(W2266), .ZN(W3462));
  NANDX1 G4235 (.A1(W973), .A2(W587), .ZN(W1095));
  NANDX1 G4236 (.A1(W603), .A2(W838), .ZN(W3164));
  NANDX1 G4237 (.A1(I170), .A2(W2086), .ZN(O390));
  NANDX1 G4238 (.A1(W422), .A2(W3023), .ZN(W3242));
  NANDX1 G4239 (.A1(W649), .A2(I575), .ZN(W1022));
  NANDX1 G4240 (.A1(W542), .A2(I236), .ZN(O414));
  NANDX1 G4241 (.A1(W346), .A2(I968), .ZN(O387));
  NANDX1 G4242 (.A1(W1056), .A2(W2664), .ZN(W3355));
  NANDX1 G4243 (.A1(W2864), .A2(W1439), .ZN(O437));
  NANDX1 G4244 (.A1(W2057), .A2(W402), .ZN(W3243));
  NANDX1 G4245 (.A1(I299), .A2(W224), .ZN(W3167));
  NANDX1 G4246 (.A1(W1995), .A2(W1039), .ZN(W3353));
  NANDX1 G4247 (.A1(W63), .A2(W1086), .ZN(W3250));
  NANDX1 G4248 (.A1(W2831), .A2(W9), .ZN(W3248));
  NANDX1 G4249 (.A1(W2507), .A2(W1170), .ZN(W3455));
  NANDX1 G4250 (.A1(W541), .A2(W563), .ZN(W3352));
  NANDX1 G4251 (.A1(W202), .A2(W3181), .ZN(W3349));
  NANDX1 G4252 (.A1(I203), .A2(I378), .ZN(W1025));
  NANDX1 G4253 (.A1(W3014), .A2(W1896), .ZN(W3350));
  NANDX1 G4254 (.A1(I633), .A2(I170), .ZN(O386));
  NANDX1 G4255 (.A1(W936), .A2(W258), .ZN(W1031));
  NANDX1 G4256 (.A1(W260), .A2(W2836), .ZN(W3152));
  NANDX1 G4257 (.A1(I174), .A2(W1648), .ZN(W3155));
  NANDX1 G4258 (.A1(W103), .A2(W2273), .ZN(W3156));
  NANDX1 G4259 (.A1(W1263), .A2(W2911), .ZN(W3182));
  NANDX1 G4260 (.A1(W1386), .A2(W2012), .ZN(O407));
  NANDX1 G4261 (.A1(I863), .A2(W1838), .ZN(W3262));
  NANDX1 G4262 (.A1(W2025), .A2(W2656), .ZN(O465));
  NANDX1 G4263 (.A1(W845), .A2(I890), .ZN(W1066));
  NANDX1 G4264 (.A1(I152), .A2(W644), .ZN(O42));
  NANDX1 G4265 (.A1(W897), .A2(W2877), .ZN(O480));
  NANDX1 G4266 (.A1(I227), .A2(W69), .ZN(W1064));
  NANDX1 G4267 (.A1(I816), .A2(I81), .ZN(W3160));
  NANDX1 G4268 (.A1(W2688), .A2(I696), .ZN(W3331));
  NANDX1 G4269 (.A1(W464), .A2(W3113), .ZN(W3259));
  NANDX1 G4270 (.A1(W1085), .A2(W1164), .ZN(W3179));
  NANDX1 G4271 (.A1(I443), .A2(I230), .ZN(W1062));
  NANDX1 G4272 (.A1(W2290), .A2(W3079), .ZN(O436));
  NANDX1 G4273 (.A1(I642), .A2(I603), .ZN(W3258));
  NANDX1 G4274 (.A1(I263), .A2(I442), .ZN(W1093));
  NANDX1 G4275 (.A1(W743), .A2(W535), .ZN(W1127));
  NANDX1 G4276 (.A1(W418), .A2(I447), .ZN(W1061));
  NANDX1 G4277 (.A1(W108), .A2(W2036), .ZN(W3163));
  NANDX1 G4278 (.A1(I28), .A2(I376), .ZN(O478));
  NANDX1 G4279 (.A1(I634), .A2(I96), .ZN(W1102));
  NANDX1 G4280 (.A1(W232), .A2(W210), .ZN(W3442));
  NANDX1 G4281 (.A1(W2639), .A2(W1517), .ZN(W3468));
  NANDX1 G4282 (.A1(W1554), .A2(W51), .ZN(W3312));
  NANDX1 G4283 (.A1(I297), .A2(W1915), .ZN(W3121));
  NANDX1 G4284 (.A1(I319), .A2(I430), .ZN(W1045));
  NANDX1 G4285 (.A1(W2729), .A2(I168), .ZN(W3287));
  NANDX1 G4286 (.A1(W1062), .A2(W829), .ZN(W1073));
  NANDX1 G4287 (.A1(W672), .A2(I175), .ZN(O40));
  NANDX1 G4288 (.A1(W768), .A2(W871), .ZN(W1141));
  NANDX1 G4289 (.A1(W2996), .A2(W1147), .ZN(W3212));
  NANDX1 G4290 (.A1(I516), .A2(I256), .ZN(W1117));
  NANDX1 G4291 (.A1(W1478), .A2(W1334), .ZN(W3106));
  NANDX1 G4292 (.A1(W2482), .A2(W33), .ZN(W3109));
  NANDX1 G4293 (.A1(W3270), .A2(W157), .ZN(O428));
  NANDX1 G4294 (.A1(W1249), .A2(W1476), .ZN(W3302));
  NANDX1 G4295 (.A1(W2441), .A2(I887), .ZN(W3123));
  NANDX1 G4296 (.A1(W2379), .A2(W2400), .ZN(O450));
  NANDX1 G4297 (.A1(I672), .A2(W2652), .ZN(W3414));
  NANDX1 G4298 (.A1(I900), .A2(W2633), .ZN(W3390));
  NANDX1 G4299 (.A1(W366), .A2(W802), .ZN(W1114));
  NANDX1 G4300 (.A1(I787), .A2(I652), .ZN(W1113));
  NANDX1 G4301 (.A1(I505), .A2(W257), .ZN(W3495));
  NANDX1 G4302 (.A1(W2572), .A2(W2758), .ZN(W3408));
  NANDX1 G4303 (.A1(I583), .A2(W1891), .ZN(W3293));
  NANDX1 G4304 (.A1(W1192), .A2(W934), .ZN(W3112));
  NANDX1 G4305 (.A1(W185), .A2(W2812), .ZN(W3411));
  NANDX1 G4306 (.A1(W2793), .A2(W1442), .ZN(O400));
  NANDX1 G4307 (.A1(W845), .A2(I800), .ZN(W1146));
  NANDX1 G4308 (.A1(W754), .A2(W278), .ZN(W3410));
  NANDX1 G4309 (.A1(W1178), .A2(W2740), .ZN(W3320));
  NANDX1 G4310 (.A1(W2334), .A2(W931), .ZN(W3115));
  NANDX1 G4311 (.A1(W1661), .A2(W1073), .ZN(W3292));
  NANDX1 G4312 (.A1(I88), .A2(I536), .ZN(W1115));
  NANDX1 G4313 (.A1(W1174), .A2(W2270), .ZN(W3396));
  NANDX1 G4314 (.A1(W1979), .A2(W888), .ZN(W3307));
  NANDX1 G4315 (.A1(I542), .A2(W2154), .ZN(W3116));
  NANDX1 G4316 (.A1(I944), .A2(W977), .ZN(W1082));
  NANDX1 G4317 (.A1(W54), .A2(W1059), .ZN(W1074));
  NANDX1 G4318 (.A1(W256), .A2(I420), .ZN(O451));
  NANDX1 G4319 (.A1(W2019), .A2(I450), .ZN(W3120));
  NANDX1 G4320 (.A1(W1790), .A2(I595), .ZN(W3288));
  NANDX1 G4321 (.A1(I647), .A2(W723), .ZN(W3110));
  NANDX1 G4322 (.A1(I245), .A2(W708), .ZN(W3298));
  NANDX1 G4323 (.A1(W265), .A2(W774), .ZN(W1077));
  NANDX1 G4324 (.A1(W2389), .A2(I592), .ZN(O488));
  NANDX1 G4325 (.A1(W2286), .A2(I746), .ZN(W3400));
  NANDX1 G4326 (.A1(W3284), .A2(W1337), .ZN(W3319));
  NANDX1 G4327 (.A1(W238), .A2(I842), .ZN(W1043));
  NANDX1 G4328 (.A1(W2794), .A2(I737), .ZN(W3318));
  NANDX1 G4329 (.A1(W44), .A2(I660), .ZN(W3218));
  NANDX1 G4330 (.A1(W2932), .A2(W2225), .ZN(O449));
  NANDX1 G4331 (.A1(I421), .A2(I774), .ZN(W1071));
  NANDX1 G4332 (.A1(W2944), .A2(I17), .ZN(W3315));
  NANDX1 G4333 (.A1(W2856), .A2(W2308), .ZN(W3314));
  NANDX1 G4334 (.A1(I549), .A2(W486), .ZN(W1139));
  INVX1 G4335 (.I(W1353), .ZN(W1462));
  INVX1 G4336 (.I(I576), .ZN(W288));
  INVX1 G4337 (.I(I448), .ZN(W224));
  INVX1 G4338 (.I(W1445), .ZN(W3731));
  INVX1 G4339 (.I(I426), .ZN(W213));
  INVX1 G4340 (.I(I188), .ZN(O1736));
  INVX1 G4341 (.I(W3648), .ZN(O1735));
  INVX1 G4342 (.I(W359), .ZN(O1734));
  INVX1 G4343 (.I(W2024), .ZN(O1856));
  INVX1 G4344 (.I(W3524), .ZN(W3689));
  INVX1 G4345 (.I(W4221), .ZN(O1733));
  INVX1 G4346 (.I(W1981), .ZN(O158));
  INVX1 G4347 (.I(W5273), .ZN(W5682));
  INVX1 G4348 (.I(W2081), .ZN(W2139));
  INVX1 G4349 (.I(W642), .ZN(W1056));
  INVX1 G4350 (.I(W305), .ZN(W3733));
  INVX1 G4351 (.I(W1333), .ZN(W2041));
  INVX1 G4352 (.I(W619), .ZN(W2157));
  INVX1 G4353 (.I(W1987), .ZN(O1729));
  INVX1 G4354 (.I(W1936), .ZN(O1728));
  INVX1 G4355 (.I(W4330), .ZN(W5874));
  INVX1 G4356 (.I(W1858), .ZN(W2024));
  INVX1 G4357 (.I(W4723), .ZN(O1706));
  INVX1 G4358 (.I(W58), .ZN(O41));
  INVX1 G4359 (.I(W4647), .ZN(W5866));
  INVX1 G4360 (.I(W174), .ZN(O1746));
  INVX1 G4361 (.I(W451), .ZN(O555));
  INVX1 G4362 (.I(I584), .ZN(W292));
  INVX1 G4363 (.I(W3248), .ZN(W3366));
  INVX1 G4364 (.I(W784), .ZN(W3748));
  INVX1 G4365 (.I(I528), .ZN(W264));
  INVX1 G4366 (.I(I318), .ZN(W1464));
  INVX1 G4367 (.I(I424), .ZN(W212));
  INVX1 G4368 (.I(W4342), .ZN(O1743));
  INVX1 G4369 (.I(W1528), .ZN(O1883));
  INVX1 G4370 (.I(W1332), .ZN(O1882));
  INVX1 G4371 (.I(W1487), .ZN(W2045));
  INVX1 G4372 (.I(W2504), .ZN(W3730));
  INVX1 G4373 (.I(W4985), .ZN(O1741));
  INVX1 G4374 (.I(W2379), .ZN(W3395));
  INVX1 G4375 (.I(W1144), .ZN(W2135));
  INVX1 G4376 (.I(W3701), .ZN(O1693));
  INVX1 G4377 (.I(W5852), .ZN(O1875));
  INVX1 G4378 (.I(I612), .ZN(O1739));
  INVX1 G4379 (.I(W199), .ZN(O164));
  INVX1 G4380 (.I(W412), .ZN(W1459));
  INVX1 G4381 (.I(I760), .ZN(W1044));
  INVX1 G4382 (.I(W2814), .ZN(O1865));
  INVX1 G4383 (.I(W906), .ZN(W2151));
  INVX1 G4384 (.I(W1357), .ZN(O552));
  INVX1 G4385 (.I(W2432), .ZN(O1717));
  INVX1 G4386 (.I(I873), .ZN(W2036));
  INVX1 G4387 (.I(W1882), .ZN(W2035));
  INVX1 G4388 (.I(I560), .ZN(W280));
  INVX1 G4389 (.I(W156), .ZN(O1715));
  INVX1 G4390 (.I(W451), .ZN(W2028));
  INVX1 G4391 (.I(W834), .ZN(W958));
  INVX1 G4392 (.I(W2523), .ZN(W3738));
  INVX1 G4393 (.I(I280), .ZN(W1452));
  INVX1 G4394 (.I(I570), .ZN(W285));
  INVX1 G4395 (.I(W4522), .ZN(O1870));
  INVX1 G4396 (.I(I276), .ZN(O1874));
  INVX1 G4397 (.I(W2487), .ZN(O438));
  INVX1 G4398 (.I(W2568), .ZN(O1711));
  INVX1 G4399 (.I(W678), .ZN(W2032));
  INVX1 G4400 (.I(W1446), .ZN(O1702));
  INVX1 G4401 (.I(W1407), .ZN(W2031));
  INVX1 G4402 (.I(I568), .ZN(W284));
  INVX1 G4403 (.I(W988), .ZN(O553));
  INVX1 G4404 (.I(I755), .ZN(W2027));
  INVX1 G4405 (.I(W2068), .ZN(W3361));
  INVX1 G4406 (.I(I544), .ZN(W272));
  INVX1 G4407 (.I(W1288), .ZN(O163));
  INVX1 G4408 (.I(I224), .ZN(W1501));
  INVX1 G4409 (.I(W4258), .ZN(O1860));
  INVX1 G4410 (.I(W1112), .ZN(W2144));
  INVX1 G4411 (.I(W224), .ZN(O1709));
  INVX1 G4412 (.I(W1320), .ZN(W1450));
  INVX1 G4413 (.I(I165), .ZN(W2039));
  INVX1 G4414 (.I(W2816), .ZN(W5700));
  INVX1 G4415 (.I(W2006), .ZN(W3364));
  INVX1 G4416 (.I(I758), .ZN(O1862));
  INVX1 G4417 (.I(W3395), .ZN(O571));
  INVX1 G4418 (.I(I60), .ZN(W2148));
  INVX1 G4419 (.I(I572), .ZN(W286));
  INVX1 G4420 (.I(W4661), .ZN(O1721));
  INVX1 G4421 (.I(W1592), .ZN(W2037));
  INVX1 G4422 (.I(I552), .ZN(W276));
  INVX1 G4423 (.I(W2978), .ZN(O1705));
  INVX1 G4424 (.I(W604), .ZN(W941));
  INVX1 G4425 (.I(W4753), .ZN(O1698));
  INVX1 G4426 (.I(I702), .ZN(O1699));
  INVX1 G4427 (.I(W1800), .ZN(W3360));
  INVX1 G4428 (.I(W4329), .ZN(O1799));
  INVX1 G4429 (.I(W4686), .ZN(O1806));
  INVX1 G4430 (.I(I486), .ZN(W243));
  INVX1 G4431 (.I(W5658), .ZN(O1835));
  INVX1 G4432 (.I(W2191), .ZN(W5843));
  INVX1 G4433 (.I(I595), .ZN(W5806));
  INVX1 G4434 (.I(W584), .ZN(W1489));
  INVX1 G4435 (.I(W2635), .ZN(O1837));
  INVX1 G4436 (.I(W5658), .ZN(O1805));
  INVX1 G4437 (.I(I161), .ZN(O148));
  INVX1 G4438 (.I(W5213), .ZN(O1802));
  INVX1 G4439 (.I(W5254), .ZN(O1801));
  INVX1 G4440 (.I(W1589), .ZN(W2060));
  INVX1 G4441 (.I(W5474), .ZN(O1840));
  INVX1 G4442 (.I(W3243), .ZN(W3388));
  INVX1 G4443 (.I(W1940), .ZN(W3712));
  INVX1 G4444 (.I(W1006), .ZN(W2095));
  INVX1 G4445 (.I(W3691), .ZN(W3713));
  INVX1 G4446 (.I(W1728), .ZN(O1841));
  INVX1 G4447 (.I(I712), .ZN(W1053));
  INVX1 G4448 (.I(W330), .ZN(W3715));
  INVX1 G4449 (.I(W2957), .ZN(O558));
  INVX1 G4450 (.I(W5582), .ZN(O1793));
  INVX1 G4451 (.I(I460), .ZN(W230));
  INVX1 G4452 (.I(I576), .ZN(W1492));
  INVX1 G4453 (.I(W2049), .ZN(O152));
  INVX1 G4454 (.I(W2569), .ZN(O1659));
  INVX1 G4455 (.I(I496), .ZN(W248));
  INVX1 G4456 (.I(I482), .ZN(W3703));
  INVX1 G4457 (.I(I798), .ZN(O1826));
  INVX1 G4458 (.I(W922), .ZN(O1825));
  INVX1 G4459 (.I(W4367), .ZN(O1824));
  INVX1 G4460 (.I(I690), .ZN(O144));
  INVX1 G4461 (.I(W152), .ZN(W1486));
  INVX1 G4462 (.I(W783), .ZN(W3386));
  INVX1 G4463 (.I(W394), .ZN(O37));
  INVX1 G4464 (.I(W1482), .ZN(W1487));
  INVX1 G4465 (.I(W962), .ZN(O1822));
  INVX1 G4466 (.I(W421), .ZN(W2073));
  INVX1 G4467 (.I(W1883), .ZN(W2074));
  INVX1 G4468 (.I(I472), .ZN(W236));
  INVX1 G4469 (.I(W76), .ZN(O70));
  INVX1 G4470 (.I(I817), .ZN(W2102));
  INVX1 G4471 (.I(W1390), .ZN(W2077));
  INVX1 G4472 (.I(I464), .ZN(W232));
  INVX1 G4473 (.I(W1859), .ZN(W2067));
  INVX1 G4474 (.I(W478), .ZN(O1832));
  INVX1 G4475 (.I(W541), .ZN(O447));
  INVX1 G4476 (.I(I995), .ZN(W1479));
  INVX1 G4477 (.I(W328), .ZN(W2086));
  INVX1 G4478 (.I(W979), .ZN(W2087));
  INVX1 G4479 (.I(W2974), .ZN(O1811));
  INVX1 G4480 (.I(W743), .ZN(W1050));
  INVX1 G4481 (.I(W164), .ZN(W1477));
  INVX1 G4482 (.I(W1865), .ZN(O1834));
  INVX1 G4483 (.I(W2772), .ZN(O1807));
  INVX1 G4484 (.I(I531), .ZN(W2049));
  INVX1 G4485 (.I(W778), .ZN(O565));
  INVX1 G4486 (.I(I512), .ZN(W256));
  INVX1 G4487 (.I(W1376), .ZN(O1767));
  INVX1 G4488 (.I(I520), .ZN(W5860));
  INVX1 G4489 (.I(I514), .ZN(W257));
  INVX1 G4490 (.I(I939), .ZN(O1765));
  INVX1 G4491 (.I(W4128), .ZN(O1764));
  INVX1 G4492 (.I(W740), .ZN(O72));
  INVX1 G4493 (.I(W312), .ZN(W2120));
  INVX1 G4494 (.I(W4617), .ZN(O1762));
  INVX1 G4495 (.I(W449), .ZN(W2121));
  INVX1 G4496 (.I(W1363), .ZN(W1468));
  INVX1 G4497 (.I(I968), .ZN(W2123));
  INVX1 G4498 (.I(W1316), .ZN(W2118));
  INVX1 G4499 (.I(W609), .ZN(W2125));
  INVX1 G4500 (.I(W1970), .ZN(O1756));
  INVX1 G4501 (.I(W2912), .ZN(O1755));
  INVX1 G4502 (.I(W1450), .ZN(W2126));
  INVX1 G4503 (.I(W1365), .ZN(O1850));
  INVX1 G4504 (.I(I426), .ZN(W2127));
  INVX1 G4505 (.I(W2273), .ZN(O1753));
  INVX1 G4506 (.I(W3837), .ZN(O1752));
  INVX1 G4507 (.I(I654), .ZN(W3726));
  INVX1 G4508 (.I(I452), .ZN(W226));
  INVX1 G4509 (.I(I522), .ZN(W261));
  INVX1 G4510 (.I(I612), .ZN(O1749));
  INVX1 G4511 (.I(W2082), .ZN(W3727));
  INVX1 G4512 (.I(W3221), .ZN(W5776));
  INVX1 G4513 (.I(I175), .ZN(O153));
  INVX1 G4514 (.I(I607), .ZN(W2104));
  INVX1 G4515 (.I(W1570), .ZN(W2056));
  INVX1 G4516 (.I(W1247), .ZN(O1786));
  INVX1 G4517 (.I(W1281), .ZN(O1784));
  INVX1 G4518 (.I(W4394), .ZN(O1783));
  INVX1 G4519 (.I(W3196), .ZN(O1782));
  INVX1 G4520 (.I(W3283), .ZN(W3393));
  INVX1 G4521 (.I(I126), .ZN(W3719));
  INVX1 G4522 (.I(W5492), .ZN(O1780));
  INVX1 G4523 (.I(I688), .ZN(W2108));
  INVX1 G4524 (.I(W1977), .ZN(O1778));
  INVX1 G4525 (.I(I758), .ZN(W1494));
  INVX1 G4526 (.I(W1273), .ZN(O567));
  INVX1 G4527 (.I(W751), .ZN(W2109));
  INVX1 G4528 (.I(W731), .ZN(W2110));
  INVX1 G4529 (.I(W3202), .ZN(W3720));
  INVX1 G4530 (.I(W403), .ZN(W2112));
  INVX1 G4531 (.I(W1257), .ZN(O1773));
  INVX1 G4532 (.I(I520), .ZN(O443));
  INVX1 G4533 (.I(W3011), .ZN(W5858));
  INVX1 G4534 (.I(W1035), .ZN(W3368));
  INVX1 G4535 (.I(W1599), .ZN(O556));
  INVX1 G4536 (.I(W1380), .ZN(O564));
  INVX1 G4537 (.I(W101), .ZN(W1469));
  INVX1 G4538 (.I(I512), .ZN(W2117));
  INVX1 G4539 (.I(W1503), .ZN(W5482));
  INVX1 G4540 (.I(I511), .ZN(W5474));
  INVX1 G4541 (.I(W461), .ZN(W1400));
  INVX1 G4542 (.I(W276), .ZN(W2307));
  INVX1 G4543 (.I(I213), .ZN(W1070));
  INVX1 G4544 (.I(W1025), .ZN(O598));
  INVX1 G4545 (.I(W2011), .ZN(W2304));
  INVX1 G4546 (.I(W2098), .ZN(W2303));
  INVX1 G4547 (.I(W3709), .ZN(O1546));
  INVX1 G4548 (.I(W3292), .ZN(O601));
  INVX1 G4549 (.I(W830), .ZN(W3801));
  INVX1 G4550 (.I(W2875), .ZN(O596));
  INVX1 G4551 (.I(W76), .ZN(W1069));
  INVX1 G4552 (.I(I429), .ZN(W3798));
  INVX1 G4553 (.I(I92), .ZN(O1549));
  INVX1 G4554 (.I(W2903), .ZN(O1550));
  INVX1 G4555 (.I(W824), .ZN(W1403));
  INVX1 G4556 (.I(W1325), .ZN(O192));
  INVX1 G4557 (.I(I750), .ZN(W375));
  INVX1 G4558 (.I(I592), .ZN(W2326));
  INVX1 G4559 (.I(I748), .ZN(W374));
  INVX1 G4560 (.I(W2396), .ZN(W5453));
  INVX1 G4561 (.I(W737), .ZN(W3317));
  INVX1 G4562 (.I(W4335), .ZN(W5457));
  INVX1 G4563 (.I(W131), .ZN(W2319));
  INVX1 G4564 (.I(I738), .ZN(W369));
  INVX1 G4565 (.I(W3104), .ZN(O432));
  INVX1 G4566 (.I(W568), .ZN(O191));
  INVX1 G4567 (.I(W1254), .ZN(W1398));
  INVX1 G4568 (.I(I253), .ZN(O1534));
  INVX1 G4569 (.I(W3750), .ZN(O1535));
  INVX1 G4570 (.I(I732), .ZN(W366));
  INVX1 G4571 (.I(W5325), .ZN(O1537));
  INVX1 G4572 (.I(W3569), .ZN(W3808));
  INVX1 G4573 (.I(W1926), .ZN(W5519));
  INVX1 G4574 (.I(I702), .ZN(W351));
  INVX1 G4575 (.I(W1093), .ZN(W2282));
  INVX1 G4576 (.I(W4939), .ZN(O1567));
  INVX1 G4577 (.I(W708), .ZN(W927));
  INVX1 G4578 (.I(W2369), .ZN(W5515));
  INVX1 G4579 (.I(I698), .ZN(W349));
  INVX1 G4580 (.I(W923), .ZN(W2277));
  INVX1 G4581 (.I(W1448), .ZN(W3789));
  INVX1 G4582 (.I(I49), .ZN(W5510));
  INVX1 G4583 (.I(I489), .ZN(O592));
  INVX1 G4584 (.I(W1746), .ZN(W2274));
  INVX1 G4585 (.I(I688), .ZN(W344));
  INVX1 G4586 (.I(W594), .ZN(O1576));
  INVX1 G4587 (.I(W157), .ZN(W3786));
  INVX1 G4588 (.I(W519), .ZN(W1068));
  INVX1 G4589 (.I(W905), .ZN(W2269));
  INVX1 G4590 (.I(I82), .ZN(W2287));
  INVX1 G4591 (.I(I590), .ZN(W3327));
  INVX1 G4592 (.I(W504), .ZN(W1405));
  INVX1 G4593 (.I(I716), .ZN(W358));
  INVX1 G4594 (.I(W1190), .ZN(W1406));
  INVX1 G4595 (.I(I477), .ZN(W5496));
  INVX1 G4596 (.I(W4902), .ZN(O1554));
  INVX1 G4597 (.I(W2360), .ZN(O1556));
  INVX1 G4598 (.I(W571), .ZN(W926));
  INVX1 G4599 (.I(W2219), .ZN(O193));
  INVX1 G4600 (.I(W1857), .ZN(O1560));
  INVX1 G4601 (.I(W67), .ZN(W3330));
  INVX1 G4602 (.I(I330), .ZN(O1562));
  INVX1 G4603 (.I(I102), .ZN(W2285));
  INVX1 G4604 (.I(I708), .ZN(O5));
  INVX1 G4605 (.I(W1647), .ZN(W3791));
  INVX1 G4606 (.I(W2251), .ZN(O186));
  INVX1 G4607 (.I(I999), .ZN(W3305));
  INVX1 G4608 (.I(W797), .ZN(W2355));
  INVX1 G4609 (.I(I946), .ZN(W1388));
  INVX1 G4610 (.I(W1625), .ZN(O1483));
  INVX1 G4611 (.I(W1318), .ZN(W2353));
  INVX1 G4612 (.I(W2912), .ZN(O1484));
  INVX1 G4613 (.I(W1788), .ZN(W3828));
  INVX1 G4614 (.I(W4355), .ZN(W5399));
  INVX1 G4615 (.I(I782), .ZN(W391));
  INVX1 G4616 (.I(W1744), .ZN(W3304));
  INVX1 G4617 (.I(W3966), .ZN(O1487));
  INVX1 G4618 (.I(W2815), .ZN(O1488));
  INVX1 G4619 (.I(W780), .ZN(W5404));
  INVX1 G4620 (.I(W501), .ZN(O1489));
  INVX1 G4621 (.I(I600), .ZN(W916));
  INVX1 G4622 (.I(W806), .ZN(O1491));
  INVX1 G4623 (.I(W332), .ZN(O199));
  INVX1 G4624 (.I(W3847), .ZN(O1472));
  INVX1 G4625 (.I(I162), .ZN(W3839));
  INVX1 G4626 (.I(I794), .ZN(W397));
  INVX1 G4627 (.I(W1213), .ZN(O1466));
  INVX1 G4628 (.I(W3471), .ZN(O1468));
  INVX1 G4629 (.I(W1653), .ZN(W2363));
  INVX1 G4630 (.I(W618), .ZN(W2362));
  INVX1 G4631 (.I(I737), .ZN(W913));
  INVX1 G4632 (.I(I400), .ZN(W2360));
  INVX1 G4633 (.I(W719), .ZN(W1391));
  INVX1 G4634 (.I(W2162), .ZN(O1473));
  INVX1 G4635 (.I(W1070), .ZN(W2359));
  INVX1 G4636 (.I(W1261), .ZN(W5386));
  INVX1 G4637 (.I(W4109), .ZN(O1475));
  INVX1 G4638 (.I(I788), .ZN(W394));
  INVX1 G4639 (.I(W512), .ZN(W1386));
  INVX1 G4640 (.I(W1718), .ZN(O1478));
  INVX1 G4641 (.I(I760), .ZN(W380));
  INVX1 G4642 (.I(W3768), .ZN(O1508));
  INVX1 G4643 (.I(W3059), .ZN(O1509));
  INVX1 G4644 (.I(I822), .ZN(W3309));
  INVX1 G4645 (.I(I580), .ZN(O1512));
  INVX1 G4646 (.I(W2218), .ZN(W2334));
  INVX1 G4647 (.I(W5290), .ZN(W5435));
  INVX1 G4648 (.I(W2223), .ZN(W2333));
  INVX1 G4649 (.I(I762), .ZN(O7));
  INVX1 G4650 (.I(W1158), .ZN(W1394));
  INVX1 G4651 (.I(I756), .ZN(W378));
  INVX1 G4652 (.I(I200), .ZN(W2330));
  INVX1 G4653 (.I(W1184), .ZN(W2329));
  INVX1 G4654 (.I(W983), .ZN(O1518));
  INVX1 G4655 (.I(W3255), .ZN(O1519));
  INVX1 G4656 (.I(W4868), .ZN(O1520));
  INVX1 G4657 (.I(W766), .ZN(W2328));
  INVX1 G4658 (.I(W3247), .ZN(O1499));
  INVX1 G4659 (.I(I774), .ZN(W387));
  INVX1 G4660 (.I(W90), .ZN(W2346));
  INVX1 G4661 (.I(W2090), .ZN(W3306));
  INVX1 G4662 (.I(W3641), .ZN(O1495));
  INVX1 G4663 (.I(W2601), .ZN(W5414));
  INVX1 G4664 (.I(W1260), .ZN(O1496));
  INVX1 G4665 (.I(W2401), .ZN(O1497));
  INVX1 G4666 (.I(W4274), .ZN(O1498));
  INVX1 G4667 (.I(I844), .ZN(O1578));
  INVX1 G4668 (.I(W3657), .ZN(O606));
  INVX1 G4669 (.I(W3784), .ZN(O605));
  INVX1 G4670 (.I(W637), .ZN(O1502));
  INVX1 G4671 (.I(I768), .ZN(O8));
  INVX1 G4672 (.I(I914), .ZN(W2340));
  INVX1 G4673 (.I(W394), .ZN(W917));
  INVX1 G4674 (.I(W3420), .ZN(O1506));
  INVX1 G4675 (.I(I701), .ZN(W2198));
  INVX1 G4676 (.I(W4123), .ZN(W5622));
  INVX1 G4677 (.I(W1914), .ZN(W5623));
  INVX1 G4678 (.I(W1050), .ZN(W3345));
  INVX1 G4679 (.I(W1702), .ZN(O171));
  INVX1 G4680 (.I(W2100), .ZN(O1653));
  INVX1 G4681 (.I(W135), .ZN(W5627));
  INVX1 G4682 (.I(W1963), .ZN(W2201));
  INVX1 G4683 (.I(I138), .ZN(W2200));
  INVX1 G4684 (.I(W2459), .ZN(W3343));
  INVX1 G4685 (.I(W3594), .ZN(O1656));
  INVX1 G4686 (.I(I616), .ZN(W308));
  INVX1 G4687 (.I(W4968), .ZN(O1658));
  INVX1 G4688 (.I(I517), .ZN(W2365));
  INVX1 G4689 (.I(I108), .ZN(W3346));
  INVX1 G4690 (.I(W1378), .ZN(W2196));
  INVX1 G4691 (.I(I610), .ZN(W305));
  INVX1 G4692 (.I(W3135), .ZN(O435));
  INVX1 G4693 (.I(W1363), .ZN(O1635));
  INVX1 G4694 (.I(I235), .ZN(W2215));
  INVX1 G4695 (.I(I868), .ZN(W2213));
  INVX1 G4696 (.I(W2968), .ZN(O1638));
  INVX1 G4697 (.I(I46), .ZN(W3765));
  INVX1 G4698 (.I(I75), .ZN(O1640));
  INVX1 G4699 (.I(W3321), .ZN(O1642));
  INVX1 G4700 (.I(I71), .ZN(O1643));
  INVX1 G4701 (.I(I923), .ZN(W1437));
  INVX1 G4702 (.I(W398), .ZN(O1645));
  INVX1 G4703 (.I(W2004), .ZN(W2209));
  INVX1 G4704 (.I(W4074), .ZN(W5615));
  INVX1 G4705 (.I(I626), .ZN(W313));
  INVX1 G4706 (.I(W2025), .ZN(W2206));
  INVX1 G4707 (.I(W3975), .ZN(O1648));
  INVX1 G4708 (.I(W3671), .ZN(W5619));
  INVX1 G4709 (.I(I590), .ZN(W295));
  INVX1 G4710 (.I(I598), .ZN(W299));
  INVX1 G4711 (.I(W4271), .ZN(W5657));
  INVX1 G4712 (.I(I945), .ZN(W1444));
  INVX1 G4713 (.I(W2160), .ZN(W3347));
  INVX1 G4714 (.I(W1289), .ZN(W3348));
  INVX1 G4715 (.I(W913), .ZN(O166));
  INVX1 G4716 (.I(W696), .ZN(W938));
  INVX1 G4717 (.I(I592), .ZN(W296));
  INVX1 G4718 (.I(W1724), .ZN(O578));
  INVX1 G4719 (.I(W884), .ZN(O574));
  INVX1 G4720 (.I(W1956), .ZN(W2173));
  INVX1 G4721 (.I(W1648), .ZN(O1683));
  INVX1 G4722 (.I(W5141), .ZN(O1684));
  INVX1 G4723 (.I(W4004), .ZN(O1685));
  INVX1 G4724 (.I(I624), .ZN(O1686));
  INVX1 G4725 (.I(I588), .ZN(W294));
  INVX1 G4726 (.I(W5409), .ZN(O1670));
  INVX1 G4727 (.I(W2010), .ZN(W2194));
  INVX1 G4728 (.I(I68), .ZN(W1439));
  INVX1 G4729 (.I(W1892), .ZN(O1664));
  INVX1 G4730 (.I(W2647), .ZN(O1665));
  INVX1 G4731 (.I(W1637), .ZN(W2191));
  INVX1 G4732 (.I(W1094), .ZN(W3757));
  INVX1 G4733 (.I(W2089), .ZN(W2189));
  INVX1 G4734 (.I(I132), .ZN(W936));
  INVX1 G4735 (.I(I335), .ZN(W2217));
  INVX1 G4736 (.I(I267), .ZN(O67));
  INVX1 G4737 (.I(I858), .ZN(O168));
  INVX1 G4738 (.I(W872), .ZN(W2183));
  INVX1 G4739 (.I(I179), .ZN(O167));
  INVX1 G4740 (.I(W3527), .ZN(O1675));
  INVX1 G4741 (.I(I349), .ZN(W5653));
  INVX1 G4742 (.I(W5275), .ZN(O1676));
  INVX1 G4743 (.I(W848), .ZN(W3776));
  INVX1 G4744 (.I(I335), .ZN(W2256));
  INVX1 G4745 (.I(W3050), .ZN(O1593));
  INVX1 G4746 (.I(W603), .ZN(W2255));
  INVX1 G4747 (.I(W1328), .ZN(O587));
  INVX1 G4748 (.I(I974), .ZN(W2252));
  INVX1 G4749 (.I(W804), .ZN(W2251));
  INVX1 G4750 (.I(W1107), .ZN(O586));
  INVX1 G4751 (.I(W3330), .ZN(O1600));
  INVX1 G4752 (.I(W208), .ZN(W2257));
  INVX1 G4753 (.I(W3027), .ZN(O1602));
  INVX1 G4754 (.I(I557), .ZN(W2248));
  INVX1 G4755 (.I(I266), .ZN(O1603));
  INVX1 G4756 (.I(W1484), .ZN(W3775));
  INVX1 G4757 (.I(I758), .ZN(W5561));
  INVX1 G4758 (.I(W1095), .ZN(W3774));
  INVX1 G4759 (.I(W193), .ZN(O181));
  INVX1 G4760 (.I(W766), .ZN(O1585));
  INVX1 G4761 (.I(W152), .ZN(W3784));
  INVX1 G4762 (.I(W3780), .ZN(W3783));
  INVX1 G4763 (.I(W2462), .ZN(W5531));
  INVX1 G4764 (.I(W1114), .ZN(W2264));
  INVX1 G4765 (.I(I936), .ZN(W929));
  INVX1 G4766 (.I(I498), .ZN(W2262));
  INVX1 G4767 (.I(W3398), .ZN(O1583));
  INVX1 G4768 (.I(W93), .ZN(W2261));
  INVX1 G4769 (.I(I666), .ZN(W333));
  INVX1 G4770 (.I(W3131), .ZN(O588));
  INVX1 G4771 (.I(W2739), .ZN(O1587));
  INVX1 G4772 (.I(W4334), .ZN(O1588));
  INVX1 G4773 (.I(W521), .ZN(O1589));
  INVX1 G4774 (.I(W1678), .ZN(W5543));
  INVX1 G4775 (.I(W4786), .ZN(O1591));
  INVX1 G4776 (.I(W908), .ZN(O1592));
  INVX1 G4777 (.I(W382), .ZN(W2228));
  INVX1 G4778 (.I(I576), .ZN(W5582));
  INVX1 G4779 (.I(I652), .ZN(W326));
  INVX1 G4780 (.I(W1982), .ZN(O1621));
  INVX1 G4781 (.I(I650), .ZN(W325));
  INVX1 G4782 (.I(W117), .ZN(O178));
  INVX1 G4783 (.I(W1528), .ZN(W3770));
  INVX1 G4784 (.I(W474), .ZN(W2229));
  INVX1 G4785 (.I(I644), .ZN(W322));
  INVX1 G4786 (.I(W1052), .ZN(W5581));
  INVX1 G4787 (.I(I828), .ZN(W2227));
  INVX1 G4788 (.I(W4878), .ZN(O1626));
  INVX1 G4789 (.I(I393), .ZN(W931));
  INVX1 G4790 (.I(I285), .ZN(W1429));
  INVX1 G4791 (.I(I247), .ZN(W2221));
  INVX1 G4792 (.I(W1519), .ZN(W2220));
  INVX1 G4793 (.I(W182), .ZN(W2218));
  INVX1 G4794 (.I(W3086), .ZN(O1689));
  INVX1 G4795 (.I(W939), .ZN(W2232));
  INVX1 G4796 (.I(W997), .ZN(W1428));
  INVX1 G4797 (.I(W1685), .ZN(W2235));
  INVX1 G4798 (.I(W2181), .ZN(W2236));
  INVX1 G4799 (.I(W1489), .ZN(W2237));
  INVX1 G4800 (.I(W2481), .ZN(O1616));
  INVX1 G4801 (.I(W4295), .ZN(O1615));
  INVX1 G4802 (.I(W1951), .ZN(O1614));
  INVX1 G4803 (.I(W1038), .ZN(W2238));
  INVX1 G4804 (.I(W1221), .ZN(W3771));
  INVX1 G4805 (.I(W372), .ZN(O585));
  INVX1 G4806 (.I(W166), .ZN(W1424));
  INVX1 G4807 (.I(I662), .ZN(W331));
  INVX1 G4808 (.I(I525), .ZN(W1422));
  INVX1 G4809 (.I(W1261), .ZN(O1607));
  INVX1 G4810 (.I(W364), .ZN(W1590));
  INVX1 G4811 (.I(W1672), .ZN(W3479));
  INVX1 G4812 (.I(W168), .ZN(W1587));
  INVX1 G4813 (.I(W835), .ZN(W1760));
  INVX1 G4814 (.I(I148), .ZN(W74));
  INVX1 G4815 (.I(W2279), .ZN(O504));
  INVX1 G4816 (.I(I18), .ZN(W1757));
  INVX1 G4817 (.I(W1860), .ZN(W3481));
  INVX1 G4818 (.I(W1526), .ZN(O103));
  INVX1 G4819 (.I(W5613), .ZN(O2249));
  INVX1 G4820 (.I(I142), .ZN(W71));
  INVX1 G4821 (.I(I140), .ZN(W70));
  INVX1 G4822 (.I(W1745), .ZN(O2262));
  INVX1 G4823 (.I(I138), .ZN(W69));
  INVX1 G4824 (.I(W2312), .ZN(W3482));
  INVX1 G4825 (.I(W130), .ZN(O502));
  INVX1 G4826 (.I(I132), .ZN(W66));
  INVX1 G4827 (.I(W4922), .ZN(O2267));
  INVX1 G4828 (.I(I158), .ZN(W79));
  INVX1 G4829 (.I(W5931), .ZN(O2232));
  INVX1 G4830 (.I(W1602), .ZN(W3566));
  INVX1 G4831 (.I(W649), .ZN(O2233));
  INVX1 G4832 (.I(W1512), .ZN(O2234));
  INVX1 G4833 (.I(W4589), .ZN(O2235));
  INVX1 G4834 (.I(W3058), .ZN(W3565));
  INVX1 G4835 (.I(W3541), .ZN(W3564));
  INVX1 G4836 (.I(I596), .ZN(W3562));
  INVX1 G4837 (.I(W2306), .ZN(O2268));
  INVX1 G4838 (.I(I95), .ZN(W1770));
  INVX1 G4839 (.I(W805), .ZN(O2242));
  INVX1 G4840 (.I(W1096), .ZN(W1769));
  INVX1 G4841 (.I(I154), .ZN(W77));
  INVX1 G4842 (.I(I583), .ZN(O2245));
  INVX1 G4843 (.I(W816), .ZN(W993));
  INVX1 G4844 (.I(I121), .ZN(O105));
  INVX1 G4845 (.I(W806), .ZN(W1766));
  INVX1 G4846 (.I(W3106), .ZN(W3550));
  INVX1 G4847 (.I(W1502), .ZN(W1598));
  INVX1 G4848 (.I(W3327), .ZN(O2285));
  INVX1 G4849 (.I(W3135), .ZN(W3483));
  INVX1 G4850 (.I(W5587), .ZN(O2287));
  INVX1 G4851 (.I(I323), .ZN(O2288));
  INVX1 G4852 (.I(I118), .ZN(W59));
  INVX1 G4853 (.I(W2534), .ZN(W3551));
  INVX1 G4854 (.I(W3190), .ZN(O2291));
  INVX1 G4855 (.I(I584), .ZN(W1597));
  INVX1 G4856 (.I(W6329), .ZN(O2293));
  INVX1 G4857 (.I(W349), .ZN(O2294));
  INVX1 G4858 (.I(I648), .ZN(W1734));
  INVX1 G4859 (.I(W1756), .ZN(O2297));
  INVX1 G4860 (.I(W2451), .ZN(O2298));
  INVX1 G4861 (.I(I762), .ZN(W3548));
  INVX1 G4862 (.I(W280), .ZN(O2300));
  INVX1 G4863 (.I(W5199), .ZN(O2301));
  INVX1 G4864 (.I(W769), .ZN(O2277));
  INVX1 G4865 (.I(I130), .ZN(W65));
  INVX1 G4866 (.I(W288), .ZN(O2270));
  INVX1 G4867 (.I(I799), .ZN(O82));
  INVX1 G4868 (.I(I151), .ZN(W996));
  INVX1 G4869 (.I(W3744), .ZN(O2273));
  INVX1 G4870 (.I(W2154), .ZN(O501));
  INVX1 G4871 (.I(W71), .ZN(W1594));
  INVX1 G4872 (.I(W904), .ZN(W1595));
  INVX1 G4873 (.I(I166), .ZN(W83));
  INVX1 G4874 (.I(I128), .ZN(W64));
  INVX1 G4875 (.I(I964), .ZN(O2278));
  INVX1 G4876 (.I(I126), .ZN(W63));
  INVX1 G4877 (.I(I124), .ZN(W62));
  INVX1 G4878 (.I(W799), .ZN(O2281));
  INVX1 G4879 (.I(W662), .ZN(W1742));
  INVX1 G4880 (.I(W5807), .ZN(O2282));
  INVX1 G4881 (.I(W1082), .ZN(W3574));
  INVX1 G4882 (.I(W1227), .ZN(O2182));
  INVX1 G4883 (.I(W5250), .ZN(O2183));
  INVX1 G4884 (.I(I901), .ZN(W1020));
  INVX1 G4885 (.I(I952), .ZN(W1806));
  INVX1 G4886 (.I(W880), .ZN(W1019));
  INVX1 G4887 (.I(I210), .ZN(W105));
  INVX1 G4888 (.I(I542), .ZN(W1803));
  INVX1 G4889 (.I(W2602), .ZN(W3474));
  INVX1 G4890 (.I(W1372), .ZN(W3471));
  INVX1 G4891 (.I(W3285), .ZN(O2190));
  INVX1 G4892 (.I(W5824), .ZN(W6237));
  INVX1 G4893 (.I(W2284), .ZN(O508));
  INVX1 G4894 (.I(W564), .ZN(O38));
  INVX1 G4895 (.I(W284), .ZN(O2193));
  INVX1 G4896 (.I(I830), .ZN(W6241));
  INVX1 G4897 (.I(W634), .ZN(O109));
  INVX1 G4898 (.I(I204), .ZN(W102));
  INVX1 G4899 (.I(I184), .ZN(W987));
  INVX1 G4900 (.I(W5561), .ZN(O2162));
  INVX1 G4901 (.I(W1664), .ZN(O2163));
  INVX1 G4902 (.I(W4), .ZN(O2164));
  INVX1 G4903 (.I(W931), .ZN(W3463));
  INVX1 G4904 (.I(W1380), .ZN(W1571));
  INVX1 G4905 (.I(W1319), .ZN(W1820));
  INVX1 G4906 (.I(W972), .ZN(W3586));
  INVX1 G4907 (.I(W103), .ZN(W986));
  INVX1 G4908 (.I(W1460), .ZN(W1578));
  INVX1 G4909 (.I(W541), .ZN(W1814));
  INVX1 G4910 (.I(W3070), .ZN(O2176));
  INVX1 G4911 (.I(W2300), .ZN(O2177));
  INVX1 G4912 (.I(W5824), .ZN(O2178));
  INVX1 G4913 (.I(I106), .ZN(W3581));
  INVX1 G4914 (.I(W2498), .ZN(W6223));
  INVX1 G4915 (.I(W296), .ZN(O477));
  INVX1 G4916 (.I(W571), .ZN(W1782));
  INVX1 G4917 (.I(W2863), .ZN(O2214));
  INVX1 G4918 (.I(W2229), .ZN(O2215));
  INVX1 G4919 (.I(I206), .ZN(W1786));
  INVX1 G4920 (.I(W2277), .ZN(O2217));
  INVX1 G4921 (.I(W448), .ZN(W1581));
  INVX1 G4922 (.I(W1111), .ZN(O2218));
  INVX1 G4923 (.I(I905), .ZN(W1784));
  INVX1 G4924 (.I(I518), .ZN(W1783));
  INVX1 G4925 (.I(I182), .ZN(W91));
  INVX1 G4926 (.I(W3277), .ZN(O2222));
  INVX1 G4927 (.I(W1149), .ZN(O2223));
  INVX1 G4928 (.I(I176), .ZN(W88));
  INVX1 G4929 (.I(W1502), .ZN(W1781));
  INVX1 G4930 (.I(W632), .ZN(W1780));
  INVX1 G4931 (.I(I172), .ZN(W86));
  INVX1 G4932 (.I(W223), .ZN(W1778));
  INVX1 G4933 (.I(W780), .ZN(W3567));
  INVX1 G4934 (.I(I879), .ZN(O108));
  INVX1 G4935 (.I(W1501), .ZN(W1796));
  INVX1 G4936 (.I(I200), .ZN(W100));
  INVX1 G4937 (.I(I198), .ZN(O2));
  INVX1 G4938 (.I(I223), .ZN(W1795));
  INVX1 G4939 (.I(W178), .ZN(O2201));
  INVX1 G4940 (.I(W1079), .ZN(O479));
  INVX1 G4941 (.I(I207), .ZN(W1793));
  INVX1 G4942 (.I(W1488), .ZN(W1792));
  INVX1 G4943 (.I(W3775), .ZN(O2302));
  INVX1 G4944 (.I(W1612), .ZN(W3569));
  INVX1 G4945 (.I(W41), .ZN(O2208));
  INVX1 G4946 (.I(I726), .ZN(W1788));
  INVX1 G4947 (.I(I188), .ZN(W94));
  INVX1 G4948 (.I(I186), .ZN(W93));
  INVX1 G4949 (.I(I710), .ZN(W1580));
  INVX1 G4950 (.I(W5076), .ZN(O2213));
  INVX1 G4951 (.I(W2708), .ZN(O2404));
  INVX1 G4952 (.I(W2449), .ZN(O2396));
  INVX1 G4953 (.I(I40), .ZN(W20));
  INVX1 G4954 (.I(W1626), .ZN(O2398));
  INVX1 G4955 (.I(W1284), .ZN(W1670));
  INVX1 G4956 (.I(I36), .ZN(W18));
  INVX1 G4957 (.I(W476), .ZN(O2401));
  INVX1 G4958 (.I(W212), .ZN(W1669));
  INVX1 G4959 (.I(W140), .ZN(W1667));
  INVX1 G4960 (.I(W1180), .ZN(O2395));
  INVX1 G4961 (.I(I34), .ZN(W17));
  INVX1 G4962 (.I(W3135), .ZN(O2406));
  INVX1 G4963 (.I(I32), .ZN(W16));
  INVX1 G4964 (.I(W809), .ZN(W1012));
  INVX1 G4965 (.I(I558), .ZN(O2409));
  INVX1 G4966 (.I(W4984), .ZN(O2410));
  INVX1 G4967 (.I(W2253), .ZN(O2411));
  INVX1 G4968 (.I(W3452), .ZN(W3520));
  INVX1 G4969 (.I(W5165), .ZN(O2386));
  INVX1 G4970 (.I(I462), .ZN(O496));
  INVX1 G4971 (.I(W5666), .ZN(O2379));
  INVX1 G4972 (.I(I350), .ZN(W3497));
  INVX1 G4973 (.I(I46), .ZN(W23));
  INVX1 G4974 (.I(I937), .ZN(W1004));
  INVX1 G4975 (.I(W2888), .ZN(W3498));
  INVX1 G4976 (.I(I526), .ZN(W3526));
  INVX1 G4977 (.I(W352), .ZN(W3499));
  INVX1 G4978 (.I(I498), .ZN(W1007));
  INVX1 G4979 (.I(W2012), .ZN(W3524));
  INVX1 G4980 (.I(W958), .ZN(W1674));
  INVX1 G4981 (.I(W6267), .ZN(O2389));
  INVX1 G4982 (.I(W66), .ZN(O2390));
  INVX1 G4983 (.I(W878), .ZN(W3500));
  INVX1 G4984 (.I(W3075), .ZN(W3522));
  INVX1 G4985 (.I(W4376), .ZN(O2393));
  INVX1 G4986 (.I(W1408), .ZN(O2394));
  INVX1 G4987 (.I(W1051), .ZN(W1647));
  INVX1 G4988 (.I(I14), .ZN(W7));
  INVX1 G4989 (.I(W1686), .ZN(O2433));
  INVX1 G4990 (.I(W2565), .ZN(W3504));
  INVX1 G4991 (.I(I64), .ZN(W1632));
  INVX1 G4992 (.I(W5331), .ZN(O2436));
  INVX1 G4993 (.I(W32), .ZN(O91));
  INVX1 G4994 (.I(W3784), .ZN(O2438));
  INVX1 G4995 (.I(W995), .ZN(O492));
  INVX1 G4996 (.I(W1668), .ZN(O2431));
  INVX1 G4997 (.I(W1203), .ZN(O90));
  INVX1 G4998 (.I(W1664), .ZN(O2442));
  INVX1 G4999 (.I(I727), .ZN(W1010));
  INVX1 G5000 (.I(W1043), .ZN(W1635));
  INVX1 G5001 (.I(W921), .ZN(W1636));
  INVX1 G5002 (.I(W2495), .ZN(O2446));
  INVX1 G5003 (.I(W1782), .ZN(O490));
  INVX1 G5004 (.I(W2000), .ZN(O491));
  INVX1 G5005 (.I(W377), .ZN(O494));
  INVX1 G5006 (.I(W2769), .ZN(O2414));
  INVX1 G5007 (.I(W1173), .ZN(W1662));
  INVX1 G5008 (.I(W1174), .ZN(W3502));
  INVX1 G5009 (.I(W1121), .ZN(O2417));
  INVX1 G5010 (.I(I24), .ZN(W12));
  INVX1 G5011 (.I(W5210), .ZN(O2419));
  INVX1 G5012 (.I(W1642), .ZN(W1658));
  INVX1 G5013 (.I(W2571), .ZN(O2422));
  INVX1 G5014 (.I(I114), .ZN(W1682));
  INVX1 G5015 (.I(W5055), .ZN(O2424));
  INVX1 G5016 (.I(W1521), .ZN(W1655));
  INVX1 G5017 (.I(W705), .ZN(W3515));
  INVX1 G5018 (.I(W842), .ZN(O2427));
  INVX1 G5019 (.I(W39), .ZN(W1653));
  INVX1 G5020 (.I(W2892), .ZN(O2429));
  INVX1 G5021 (.I(W4315), .ZN(O2430));
  INVX1 G5022 (.I(W1691), .ZN(W1717));
  INVX1 G5023 (.I(W2753), .ZN(W3546));
  INVX1 G5024 (.I(W1035), .ZN(W1604));
  INVX1 G5025 (.I(W917), .ZN(O2323));
  INVX1 G5026 (.I(W1388), .ZN(W3486));
  INVX1 G5027 (.I(I88), .ZN(W44));
  INVX1 G5028 (.I(W1623), .ZN(O2326));
  INVX1 G5029 (.I(I86), .ZN(W43));
  INVX1 G5030 (.I(W331), .ZN(O39));
  INVX1 G5031 (.I(W1200), .ZN(W1724));
  INVX1 G5032 (.I(W3636), .ZN(O2330));
  INVX1 G5033 (.I(W638), .ZN(W1715));
  INVX1 G5034 (.I(W6226), .ZN(O2332));
  INVX1 G5035 (.I(I82), .ZN(W41));
  INVX1 G5036 (.I(W4542), .ZN(O2334));
  INVX1 G5037 (.I(W1254), .ZN(W1714));
  INVX1 G5038 (.I(W1524), .ZN(W1712));
  INVX1 G5039 (.I(I76), .ZN(W38));
  INVX1 G5040 (.I(I104), .ZN(W52));
  INVX1 G5041 (.I(W1525), .ZN(W1601));
  INVX1 G5042 (.I(W2099), .ZN(O2305));
  INVX1 G5043 (.I(W402), .ZN(W1729));
  INVX1 G5044 (.I(I542), .ZN(W1728));
  INVX1 G5045 (.I(W2674), .ZN(O2308));
  INVX1 G5046 (.I(W7), .ZN(W1602));
  INVX1 G5047 (.I(W5866), .ZN(O2310));
  INVX1 G5048 (.I(I106), .ZN(W53));
  INVX1 G5049 (.I(I773), .ZN(W1708));
  INVX1 G5050 (.I(I832), .ZN(W1603));
  INVX1 G5051 (.I(I100), .ZN(W50));
  INVX1 G5052 (.I(I98), .ZN(W49));
  INVX1 G5053 (.I(W3223), .ZN(O2316));
  INVX1 G5054 (.I(I96), .ZN(W48));
  INVX1 G5055 (.I(I65), .ZN(W1725));
  INVX1 G5056 (.I(I92), .ZN(W46));
  INVX1 G5057 (.I(W579), .ZN(W1003));
  INVX1 G5058 (.I(W2680), .ZN(O2359));
  INVX1 G5059 (.I(I58), .ZN(W29));
  INVX1 G5060 (.I(W970), .ZN(O87));
  INVX1 G5061 (.I(W4032), .ZN(O2362));
  INVX1 G5062 (.I(W1301), .ZN(W3536));
  INVX1 G5063 (.I(W553), .ZN(W1623));
  INVX1 G5064 (.I(W4767), .ZN(O2366));
  INVX1 G5065 (.I(I468), .ZN(W3534));
  INVX1 G5066 (.I(W756), .ZN(O498));
  INVX1 G5067 (.I(W5531), .ZN(O2369));
  INVX1 G5068 (.I(I62), .ZN(W1685));
  INVX1 G5069 (.I(W3250), .ZN(W3532));
  INVX1 G5070 (.I(W1673), .ZN(O2372));
  INVX1 G5071 (.I(W5400), .ZN(O2373));
  INVX1 G5072 (.I(I34), .ZN(W1013));
  INVX1 G5073 (.I(I52), .ZN(W26));
  INVX1 G5074 (.I(W5314), .ZN(O2376));
  INVX1 G5075 (.I(W254), .ZN(W1614));
  INVX1 G5076 (.I(W1235), .ZN(W1612));
  INVX1 G5077 (.I(W3348), .ZN(O2342));
  INVX1 G5078 (.I(I72), .ZN(W36));
  INVX1 G5079 (.I(W104), .ZN(W1706));
  INVX1 G5080 (.I(I711), .ZN(W1613));
  INVX1 G5081 (.I(I68), .ZN(W34));
  INVX1 G5082 (.I(W250), .ZN(O486));
  INVX1 G5083 (.I(I432), .ZN(O96));
  INVX1 G5084 (.I(W1028), .ZN(O2161));
  INVX1 G5085 (.I(I66), .ZN(W33));
  INVX1 G5086 (.I(W185), .ZN(W3494));
  INVX1 G5087 (.I(I62), .ZN(W31));
  INVX1 G5088 (.I(W515), .ZN(W1618));
  INVX1 G5089 (.I(W80), .ZN(W1002));
  INVX1 G5090 (.I(W4808), .ZN(O2356));
  INVX1 G5091 (.I(W98), .ZN(W1619));
  INVX1 G5092 (.I(W361), .ZN(O1978));
  INVX1 G5093 (.I(W743), .ZN(W3654));
  INVX1 G5094 (.I(W1826), .ZN(O1971));
  INVX1 G5095 (.I(W3296), .ZN(W3421));
  INVX1 G5096 (.I(W4608), .ZN(O1973));
  INVX1 G5097 (.I(I368), .ZN(W184));
  INVX1 G5098 (.I(I366), .ZN(W183));
  INVX1 G5099 (.I(W854), .ZN(W3422));
  INVX1 G5100 (.I(W27), .ZN(W1959));
  INVX1 G5101 (.I(I222), .ZN(W1964));
  INVX1 G5102 (.I(W2941), .ZN(O541));
  INVX1 G5103 (.I(I203), .ZN(O1980));
  INVX1 G5104 (.I(W3182), .ZN(O456));
  INVX1 G5105 (.I(I362), .ZN(W181));
  INVX1 G5106 (.I(I706), .ZN(W1954));
  INVX1 G5107 (.I(I528), .ZN(W1953));
  INVX1 G5108 (.I(W3281), .ZN(O539));
  INVX1 G5109 (.I(W1073), .ZN(W1951));
  INVX1 G5110 (.I(I376), .ZN(W188));
  INVX1 G5111 (.I(W2921), .ZN(O544));
  INVX1 G5112 (.I(I734), .ZN(O454));
  INVX1 G5113 (.I(W5863), .ZN(O1955));
  INVX1 G5114 (.I(I380), .ZN(W190));
  INVX1 G5115 (.I(W189), .ZN(W1519));
  INVX1 G5116 (.I(W1733), .ZN(W3658));
  INVX1 G5117 (.I(I378), .ZN(W189));
  INVX1 G5118 (.I(I380), .ZN(O1960));
  INVX1 G5119 (.I(W2632), .ZN(W3646));
  INVX1 G5120 (.I(I613), .ZN(W1521));
  INVX1 G5121 (.I(I269), .ZN(W1038));
  INVX1 G5122 (.I(W392), .ZN(W1037));
  INVX1 G5123 (.I(W2923), .ZN(W3419));
  INVX1 G5124 (.I(W4028), .ZN(O1964));
  INVX1 G5125 (.I(W4554), .ZN(O1965));
  INVX1 G5126 (.I(I372), .ZN(W186));
  INVX1 G5127 (.I(W4492), .ZN(O1967));
  INVX1 G5128 (.I(W56), .ZN(W1534));
  INVX1 G5129 (.I(W4063), .ZN(W6034));
  INVX1 G5130 (.I(I240), .ZN(W1933));
  INVX1 G5131 (.I(I340), .ZN(W170));
  INVX1 G5132 (.I(W5000), .ZN(O2006));
  INVX1 G5133 (.I(W5577), .ZN(O2007));
  INVX1 G5134 (.I(I695), .ZN(W6039));
  INVX1 G5135 (.I(I819), .ZN(O459));
  INVX1 G5136 (.I(W1302), .ZN(O2009));
  INVX1 G5137 (.I(I342), .ZN(W171));
  INVX1 G5138 (.I(W432), .ZN(W1034));
  INVX1 G5139 (.I(I332), .ZN(W166));
  INVX1 G5140 (.I(W2712), .ZN(O534));
  INVX1 G5141 (.I(I586), .ZN(W1927));
  INVX1 G5142 (.I(I217), .ZN(W971));
  INVX1 G5143 (.I(W1456), .ZN(W1925));
  INVX1 G5144 (.I(W1078), .ZN(O2018));
  INVX1 G5145 (.I(W4174), .ZN(O2019));
  INVX1 G5146 (.I(W1769), .ZN(W3640));
  INVX1 G5147 (.I(W1154), .ZN(W3425));
  INVX1 G5148 (.I(I358), .ZN(W179));
  INVX1 G5149 (.I(I390), .ZN(O537));
  INVX1 G5150 (.I(W1833), .ZN(O1990));
  INVX1 G5151 (.I(W1231), .ZN(O1991));
  INVX1 G5152 (.I(W43), .ZN(W3428));
  INVX1 G5153 (.I(I877), .ZN(O128));
  INVX1 G5154 (.I(W1007), .ZN(W1941));
  INVX1 G5155 (.I(W2248), .ZN(O1952));
  INVX1 G5156 (.I(I842), .ZN(W1939));
  INVX1 G5157 (.I(W429), .ZN(W3430));
  INVX1 G5158 (.I(I120), .ZN(W3431));
  INVX1 G5159 (.I(W2997), .ZN(O1999));
  INVX1 G5160 (.I(W810), .ZN(O536));
  INVX1 G5161 (.I(I344), .ZN(W172));
  INVX1 G5162 (.I(W2410), .ZN(O458));
  INVX1 G5163 (.I(W158), .ZN(W5928));
  INVX1 G5164 (.I(W1878), .ZN(O1902));
  INVX1 G5165 (.I(I103), .ZN(W2010));
  INVX1 G5166 (.I(W1501), .ZN(W2009));
  INVX1 G5167 (.I(I723), .ZN(W3674));
  INVX1 G5168 (.I(I547), .ZN(W2007));
  INVX1 G5169 (.I(W231), .ZN(W3406));
  INVX1 G5170 (.I(W1464), .ZN(O1908));
  INVX1 G5171 (.I(W167), .ZN(W3407));
  INVX1 G5172 (.I(W451), .ZN(O548));
  INVX1 G5173 (.I(W485), .ZN(O1910));
  INVX1 G5174 (.I(W49), .ZN(W2004));
  INVX1 G5175 (.I(W4642), .ZN(W5931));
  INVX1 G5176 (.I(I410), .ZN(W205));
  INVX1 G5177 (.I(I313), .ZN(W2003));
  INVX1 G5178 (.I(W994), .ZN(W1507));
  INVX1 G5179 (.I(W867), .ZN(W3671));
  INVX1 G5180 (.I(W441), .ZN(W1509));
  INVX1 G5181 (.I(I418), .ZN(W209));
  INVX1 G5182 (.I(I98), .ZN(W2020));
  INVX1 G5183 (.I(W5679), .ZN(O1887));
  INVX1 G5184 (.I(W1705), .ZN(O1888));
  INVX1 G5185 (.I(W3287), .ZN(W3680));
  INVX1 G5186 (.I(W1450), .ZN(W3403));
  INVX1 G5187 (.I(W119), .ZN(O453));
  INVX1 G5188 (.I(W2396), .ZN(O1892));
  INVX1 G5189 (.I(W1947), .ZN(W3677));
  INVX1 G5190 (.I(W3494), .ZN(W3670));
  INVX1 G5191 (.I(W5776), .ZN(O1894));
  INVX1 G5192 (.I(W1707), .ZN(W2015));
  INVX1 G5193 (.I(W4146), .ZN(O1896));
  INVX1 G5194 (.I(W17), .ZN(W3676));
  INVX1 G5195 (.I(W1846), .ZN(W2012));
  INVX1 G5196 (.I(W517), .ZN(O1899));
  INVX1 G5197 (.I(W4379), .ZN(O1900));
  INVX1 G5198 (.I(I382), .ZN(W191));
  INVX1 G5199 (.I(I394), .ZN(W197));
  INVX1 G5200 (.I(W829), .ZN(W3413));
  INVX1 G5201 (.I(W5386), .ZN(O1938));
  INVX1 G5202 (.I(W515), .ZN(W1984));
  INVX1 G5203 (.I(W5010), .ZN(O1940));
  INVX1 G5204 (.I(W264), .ZN(W1983));
  INVX1 G5205 (.I(W1340), .ZN(W3663));
  INVX1 G5206 (.I(W295), .ZN(W1515));
  INVX1 G5207 (.I(W5567), .ZN(O1935));
  INVX1 G5208 (.I(W369), .ZN(W1979));
  INVX1 G5209 (.I(I744), .ZN(O1945));
  INVX1 G5210 (.I(W4615), .ZN(O1946));
  INVX1 G5211 (.I(W2589), .ZN(W3662));
  INVX1 G5212 (.I(W236), .ZN(W3415));
  INVX1 G5213 (.I(I431), .ZN(W1975));
  INVX1 G5214 (.I(W952), .ZN(O1950));
  INVX1 G5215 (.I(I117), .ZN(W1517));
  INVX1 G5216 (.I(W797), .ZN(W1512));
  INVX1 G5217 (.I(I402), .ZN(W201));
  INVX1 G5218 (.I(W1351), .ZN(W1510));
  INVX1 G5219 (.I(W5748), .ZN(O1919));
  INVX1 G5220 (.I(I356), .ZN(O1921));
  INVX1 G5221 (.I(I398), .ZN(W199));
  INVX1 G5222 (.I(W2169), .ZN(O1924));
  INVX1 G5223 (.I(I464), .ZN(W1992));
  INVX1 G5224 (.I(W985), .ZN(O1926));
  INVX1 G5225 (.I(W3457), .ZN(W3630));
  INVX1 G5226 (.I(I396), .ZN(W198));
  INVX1 G5227 (.I(W2965), .ZN(O1929));
  INVX1 G5228 (.I(W1380), .ZN(W1989));
  INVX1 G5229 (.I(I594), .ZN(W1987));
  INVX1 G5230 (.I(I624), .ZN(O1932));
  INVX1 G5231 (.I(W4298), .ZN(O1933));
  INVX1 G5232 (.I(W3205), .ZN(W3666));
  INVX1 G5233 (.I(I229), .ZN(W3605));
  INVX1 G5234 (.I(I992), .ZN(W1867));
  INVX1 G5235 (.I(W1342), .ZN(W1554));
  INVX1 G5236 (.I(I822), .ZN(O116));
  INVX1 G5237 (.I(W615), .ZN(O2111));
  INVX1 G5238 (.I(W2124), .ZN(W3607));
  INVX1 G5239 (.I(W79), .ZN(W1862));
  INVX1 G5240 (.I(I715), .ZN(W980));
  INVX1 G5241 (.I(W1746), .ZN(W1859));
  INVX1 G5242 (.I(I953), .ZN(W1026));
  INVX1 G5243 (.I(W5985), .ZN(O2116));
  INVX1 G5244 (.I(W1247), .ZN(O471));
  INVX1 G5245 (.I(W1470), .ZN(W1856));
  INVX1 G5246 (.I(W3960), .ZN(O2119));
  INVX1 G5247 (.I(I839), .ZN(O2120));
  INVX1 G5248 (.I(I771), .ZN(O2121));
  INVX1 G5249 (.I(W183), .ZN(O2123));
  INVX1 G5250 (.I(I945), .ZN(W3602));
  INVX1 G5251 (.I(W1015), .ZN(O118));
  INVX1 G5252 (.I(I658), .ZN(W1878));
  INVX1 G5253 (.I(I7), .ZN(O2091));
  INVX1 G5254 (.I(W5057), .ZN(O2092));
  INVX1 G5255 (.I(W1933), .ZN(O2093));
  INVX1 G5256 (.I(W610), .ZN(W3446));
  INVX1 G5257 (.I(W826), .ZN(O2094));
  INVX1 G5258 (.I(W3771), .ZN(O2096));
  INVX1 G5259 (.I(I235), .ZN(O2097));
  INVX1 G5260 (.I(W5425), .ZN(O2125));
  INVX1 G5261 (.I(W1742), .ZN(O2099));
  INVX1 G5262 (.I(W3687), .ZN(O2100));
  INVX1 G5263 (.I(I291), .ZN(W1029));
  INVX1 G5264 (.I(I264), .ZN(W132));
  INVX1 G5265 (.I(W3070), .ZN(W3610));
  INVX1 G5266 (.I(W1365), .ZN(W1871));
  INVX1 G5267 (.I(W3300), .ZN(O470));
  INVX1 G5268 (.I(I415), .ZN(W1869));
  INVX1 G5269 (.I(W48), .ZN(W1567));
  INVX1 G5270 (.I(W3224), .ZN(O2144));
  INVX1 G5271 (.I(W4712), .ZN(W6186));
  INVX1 G5272 (.I(W592), .ZN(W3597));
  INVX1 G5273 (.I(W2270), .ZN(O517));
  INVX1 G5274 (.I(I630), .ZN(W1838));
  INVX1 G5275 (.I(I918), .ZN(O516));
  INVX1 G5276 (.I(W2514), .ZN(W3457));
  INVX1 G5277 (.I(I688), .ZN(W3458));
  INVX1 G5278 (.I(W1484), .ZN(O518));
  INVX1 G5279 (.I(W5139), .ZN(O2153));
  INVX1 G5280 (.I(W1843), .ZN(O2154));
  INVX1 G5281 (.I(I145), .ZN(O513));
  INVX1 G5282 (.I(I365), .ZN(O114));
  INVX1 G5283 (.I(W816), .ZN(W1827));
  INVX1 G5284 (.I(W4881), .ZN(O2158));
  INVX1 G5285 (.I(I520), .ZN(W1826));
  INVX1 G5286 (.I(I100), .ZN(O2160));
  INVX1 G5287 (.I(W326), .ZN(W3456));
  INVX1 G5288 (.I(W326), .ZN(W1852));
  INVX1 G5289 (.I(W3729), .ZN(O2127));
  INVX1 G5290 (.I(W281), .ZN(W1850));
  INVX1 G5291 (.I(W3957), .ZN(O2130));
  INVX1 G5292 (.I(I272), .ZN(W1849));
  INVX1 G5293 (.I(I250), .ZN(W125));
  INVX1 G5294 (.I(W2524), .ZN(O2133));
  INVX1 G5295 (.I(I238), .ZN(W1848));
  INVX1 G5296 (.I(W488), .ZN(W1030));
  INVX1 G5297 (.I(W1785), .ZN(O2136));
  INVX1 G5298 (.I(W121), .ZN(W981));
  INVX1 G5299 (.I(W802), .ZN(W1843));
  INVX1 G5300 (.I(I357), .ZN(W1563));
  INVX1 G5301 (.I(W449), .ZN(O2140));
  INVX1 G5302 (.I(W3297), .ZN(O2141));
  INVX1 G5303 (.I(W4641), .ZN(O2142));
  INVX1 G5304 (.I(I525), .ZN(W974));
  INVX1 G5305 (.I(I266), .ZN(W1910));
  INVX1 G5306 (.I(W5987), .ZN(O2040));
  INVX1 G5307 (.I(I310), .ZN(W155));
  INVX1 G5308 (.I(W1518), .ZN(O2041));
  INVX1 G5309 (.I(W983), .ZN(O2042));
  INVX1 G5310 (.I(W3992), .ZN(O2043));
  INVX1 G5311 (.I(W2478), .ZN(O2044));
  INVX1 G5312 (.I(I712), .ZN(W1539));
  INVX1 G5313 (.I(W4291), .ZN(O2038));
  INVX1 G5314 (.I(I306), .ZN(W153));
  INVX1 G5315 (.I(W1686), .ZN(O464));
  INVX1 G5316 (.I(I555), .ZN(W1906));
  INVX1 G5317 (.I(W898), .ZN(W3622));
  INVX1 G5318 (.I(W2608), .ZN(W6087));
  INVX1 G5319 (.I(W500), .ZN(W3441));
  INVX1 G5320 (.I(W2287), .ZN(O2052));
  INVX1 G5321 (.I(I445), .ZN(W1902));
  INVX1 G5322 (.I(W1263), .ZN(O2028));
  INVX1 G5323 (.I(W4726), .ZN(O2021));
  INVX1 G5324 (.I(W2752), .ZN(O2022));
  INVX1 G5325 (.I(W616), .ZN(O126));
  INVX1 G5326 (.I(W3118), .ZN(O2023));
  INVX1 G5327 (.I(I326), .ZN(W163));
  INVX1 G5328 (.I(W283), .ZN(O125));
  INVX1 G5329 (.I(I324), .ZN(W162));
  INVX1 G5330 (.I(I843), .ZN(O2027));
  INVX1 G5331 (.I(I332), .ZN(W1542));
  INVX1 G5332 (.I(I320), .ZN(W160));
  INVX1 G5333 (.I(W3045), .ZN(O531));
  INVX1 G5334 (.I(W213), .ZN(O2031));
  INVX1 G5335 (.I(W1001), .ZN(W1538));
  INVX1 G5336 (.I(I301), .ZN(W1915));
  INVX1 G5337 (.I(W1049), .ZN(O529));
  INVX1 G5338 (.I(W616), .ZN(W1912));
  INVX1 G5339 (.I(W783), .ZN(W1883));
  INVX1 G5340 (.I(W1137), .ZN(O526));
  INVX1 G5341 (.I(I254), .ZN(W1545));
  INVX1 G5342 (.I(W665), .ZN(W1889));
  INVX1 G5343 (.I(W766), .ZN(W1546));
  INVX1 G5344 (.I(W3913), .ZN(O2075));
  INVX1 G5345 (.I(I286), .ZN(W143));
  INVX1 G5346 (.I(W2987), .ZN(O525));
  INVX1 G5347 (.I(I80), .ZN(O2079));
  INVX1 G5348 (.I(I292), .ZN(W146));
  INVX1 G5349 (.I(I280), .ZN(W140));
  INVX1 G5350 (.I(I278), .ZN(W139));
  INVX1 G5351 (.I(I623), .ZN(W1882));
  INVX1 G5352 (.I(W1517), .ZN(O466));
  INVX1 G5353 (.I(I274), .ZN(W137));
  INVX1 G5354 (.I(W2160), .ZN(O2087));
  INVX1 G5355 (.I(W4659), .ZN(O2088));
  INVX1 G5356 (.I(I272), .ZN(W136));
  INVX1 G5357 (.I(W494), .ZN(W1894));
  INVX1 G5358 (.I(W3257), .ZN(O2055));
  INVX1 G5359 (.I(W795), .ZN(W1900));
  INVX1 G5360 (.I(I808), .ZN(W1899));
  INVX1 G5361 (.I(W3980), .ZN(O2058));
  INVX1 G5362 (.I(W1073), .ZN(W1898));
  INVX1 G5363 (.I(W1989), .ZN(O2060));
  INVX1 G5364 (.I(W881), .ZN(W1896));
  INVX1 G5365 (.I(W731), .ZN(W1544));
  INVX1 G5366 (.I(W2187), .ZN(W3402));
  INVX1 G5367 (.I(W5267), .ZN(W6101));
  INVX1 G5368 (.I(W1171), .ZN(O2064));
  INVX1 G5369 (.I(W1210), .ZN(O121));
  INVX1 G5370 (.I(W1157), .ZN(W1892));
  INVX1 G5371 (.I(W3770), .ZN(O2067));
  INVX1 G5372 (.I(I294), .ZN(W147));
  INVX1 G5373 (.I(W5296), .ZN(O2069));
  INVX1 G5374 (.I(W879), .ZN(W1236));
  INVX1 G5375 (.I(W247), .ZN(W4567));
  INVX1 G5376 (.I(W4204), .ZN(O954));
  INVX1 G5377 (.I(W2163), .ZN(O955));
  INVX1 G5378 (.I(W4416), .ZN(O956));
  INVX1 G5379 (.I(W2886), .ZN(O711));
  INVX1 G5380 (.I(I92), .ZN(W1235));
  INVX1 G5381 (.I(W1985), .ZN(O308));
  INVX1 G5382 (.I(W1465), .ZN(O958));
  INVX1 G5383 (.I(W1296), .ZN(O953));
  INVX1 G5384 (.I(W2821), .ZN(O391));
  INVX1 G5385 (.I(W1557), .ZN(W2854));
  INVX1 G5386 (.I(W2139), .ZN(W4579));
  INVX1 G5387 (.I(I746), .ZN(O29));
  INVX1 G5388 (.I(W2708), .ZN(O304));
  INVX1 G5389 (.I(W3063), .ZN(W4582));
  INVX1 G5390 (.I(W981), .ZN(W3177));
  INVX1 G5391 (.I(W738), .ZN(W4584));
  INVX1 G5392 (.I(W646), .ZN(W680));
  INVX1 G5393 (.I(W3730), .ZN(W4549));
  INVX1 G5394 (.I(I72), .ZN(W833));
  INVX1 G5395 (.I(W2323), .ZN(O945));
  INVX1 G5396 (.I(I458), .ZN(W834));
  INVX1 G5397 (.I(I672), .ZN(W2868));
  INVX1 G5398 (.I(W97), .ZN(O389));
  INVX1 G5399 (.I(W3421), .ZN(W4555));
  INVX1 G5400 (.I(I209), .ZN(W681));
  INVX1 G5401 (.I(W1085), .ZN(W2849));
  INVX1 G5402 (.I(W2460), .ZN(W3174));
  INVX1 G5403 (.I(W2545), .ZN(O714));
  INVX1 G5404 (.I(W286), .ZN(W4560));
  INVX1 G5405 (.I(I797), .ZN(O949));
  INVX1 G5406 (.I(W782), .ZN(O713));
  INVX1 G5407 (.I(W68), .ZN(W1233));
  INVX1 G5408 (.I(W1036), .ZN(W2862));
  INVX1 G5409 (.I(W873), .ZN(O952));
  INVX1 G5410 (.I(W658), .ZN(W662));
  INVX1 G5411 (.I(W4113), .ZN(W4605));
  INVX1 G5412 (.I(W1062), .ZN(W1240));
  INVX1 G5413 (.I(W34), .ZN(W2836));
  INVX1 G5414 (.I(W475), .ZN(W2835));
  INVX1 G5415 (.I(W173), .ZN(W4609));
  INVX1 G5416 (.I(W2124), .ZN(W3180));
  INVX1 G5417 (.I(I565), .ZN(O707));
  INVX1 G5418 (.I(W2746), .ZN(O974));
  INVX1 G5419 (.I(W923), .ZN(W2838));
  INVX1 G5420 (.I(W1314), .ZN(O975));
  INVX1 G5421 (.I(W569), .ZN(W661));
  INVX1 G5422 (.I(W2781), .ZN(O976));
  INVX1 G5423 (.I(W1940), .ZN(W4617));
  INVX1 G5424 (.I(W1861), .ZN(W2832));
  INVX1 G5425 (.I(W3502), .ZN(O978));
  INVX1 G5426 (.I(W235), .ZN(W660));
  INVX1 G5427 (.I(I702), .ZN(W1126));
  INVX1 G5428 (.I(W4148), .ZN(O967));
  INVX1 G5429 (.I(W3634), .ZN(W4586));
  INVX1 G5430 (.I(I983), .ZN(O963));
  INVX1 G5431 (.I(W276), .ZN(O302));
  INVX1 G5432 (.I(W429), .ZN(W669));
  INVX1 G5433 (.I(I925), .ZN(W2846));
  INVX1 G5434 (.I(W1484), .ZN(O965));
  INVX1 G5435 (.I(I711), .ZN(W4593));
  INVX1 G5436 (.I(W670), .ZN(W2843));
  INVX1 G5437 (.I(W4410), .ZN(W4548));
  INVX1 G5438 (.I(I742), .ZN(W4596));
  INVX1 G5439 (.I(W2964), .ZN(W4597));
  INVX1 G5440 (.I(W1545), .ZN(W4598));
  INVX1 G5441 (.I(W970), .ZN(O968));
  INVX1 G5442 (.I(W765), .ZN(W4051));
  INVX1 G5443 (.I(W2010), .ZN(W2840));
  INVX1 G5444 (.I(W129), .ZN(W2839));
  INVX1 G5445 (.I(W701), .ZN(W1219));
  INVX1 G5446 (.I(W1237), .ZN(O916));
  INVX1 G5447 (.I(W968), .ZN(O917));
  INVX1 G5448 (.I(W2423), .ZN(W4079));
  INVX1 G5449 (.I(W3117), .ZN(O918));
  INVX1 G5450 (.I(W365), .ZN(W4497));
  INVX1 G5451 (.I(W3796), .ZN(W4499));
  INVX1 G5452 (.I(W1707), .ZN(O919));
  INVX1 G5453 (.I(W590), .ZN(W4501));
  INVX1 G5454 (.I(W3775), .ZN(W4492));
  INVX1 G5455 (.I(W3634), .ZN(O920));
  INVX1 G5456 (.I(W2598), .ZN(W4077));
  INVX1 G5457 (.I(W1488), .ZN(W4505));
  INVX1 G5458 (.I(I11), .ZN(W701));
  INVX1 G5459 (.I(W1905), .ZN(O921));
  INVX1 G5460 (.I(W4380), .ZN(W4509));
  INVX1 G5461 (.I(W913), .ZN(O922));
  INVX1 G5462 (.I(W510), .ZN(W700));
  INVX1 G5463 (.I(W3025), .ZN(W4484));
  INVX1 G5464 (.I(W2842), .ZN(W2908));
  INVX1 G5465 (.I(I213), .ZN(W2907));
  INVX1 G5466 (.I(W495), .ZN(W4478));
  INVX1 G5467 (.I(I222), .ZN(O909));
  INVX1 G5468 (.I(I999), .ZN(W704));
  INVX1 G5469 (.I(W2277), .ZN(O910));
  INVX1 G5470 (.I(W2760), .ZN(W4482));
  INVX1 G5471 (.I(W2013), .ZN(O322));
  INVX1 G5472 (.I(W1472), .ZN(W3166));
  INVX1 G5473 (.I(I8), .ZN(W1217));
  INVX1 G5474 (.I(W3335), .ZN(W4486));
  INVX1 G5475 (.I(W21), .ZN(O912));
  INVX1 G5476 (.I(W338), .ZN(O913));
  INVX1 G5477 (.I(W546), .ZN(W1218));
  INVX1 G5478 (.I(I938), .ZN(O915));
  INVX1 G5479 (.I(W1748), .ZN(W2903));
  INVX1 G5480 (.I(I967), .ZN(O388));
  INVX1 G5481 (.I(I347), .ZN(W690));
  INVX1 G5482 (.I(W2664), .ZN(O721));
  INVX1 G5483 (.I(W3430), .ZN(O720));
  INVX1 G5484 (.I(W685), .ZN(W830));
  INVX1 G5485 (.I(I911), .ZN(W2883));
  INVX1 G5486 (.I(W2170), .ZN(O316));
  INVX1 G5487 (.I(I401), .ZN(W4537));
  INVX1 G5488 (.I(W1292), .ZN(O315));
  INVX1 G5489 (.I(I91), .ZN(W691));
  INVX1 G5490 (.I(W528), .ZN(W4067));
  INVX1 G5491 (.I(W2725), .ZN(O939));
  INVX1 G5492 (.I(I262), .ZN(W684));
  INVX1 G5493 (.I(W1615), .ZN(W3169));
  INVX1 G5494 (.I(W15), .ZN(W3170));
  INVX1 G5495 (.I(W913), .ZN(W2873));
  INVX1 G5496 (.I(W2269), .ZN(O943));
  INVX1 G5497 (.I(W2372), .ZN(W3172));
  INVX1 G5498 (.I(W2026), .ZN(W4074));
  INVX1 G5499 (.I(W1041), .ZN(O925));
  INVX1 G5500 (.I(I727), .ZN(W699));
  INVX1 G5501 (.I(I308), .ZN(W1222));
  INVX1 G5502 (.I(I782), .ZN(O926));
  INVX1 G5503 (.I(W2062), .ZN(W2895));
  INVX1 G5504 (.I(W4182), .ZN(W4518));
  INVX1 G5505 (.I(W4368), .ZN(W4519));
  INVX1 G5506 (.I(I250), .ZN(W696));
  INVX1 G5507 (.I(W3257), .ZN(O980));
  INVX1 G5508 (.I(W3921), .ZN(W4073));
  INVX1 G5509 (.I(I437), .ZN(W1223));
  INVX1 G5510 (.I(I456), .ZN(W1224));
  INVX1 G5511 (.I(W3498), .ZN(W4526));
  INVX1 G5512 (.I(W1150), .ZN(W2889));
  INVX1 G5513 (.I(W661), .ZN(W2888));
  INVX1 G5514 (.I(W1772), .ZN(O930));
  INVX1 G5515 (.I(W1655), .ZN(W2763));
  INVX1 G5516 (.I(W3582), .ZN(O1032));
  INVX1 G5517 (.I(W2639), .ZN(O1033));
  INVX1 G5518 (.I(W67), .ZN(W2766));
  INVX1 G5519 (.I(W3956), .ZN(O1035));
  INVX1 G5520 (.I(W589), .ZN(W626));
  INVX1 G5521 (.I(W1582), .ZN(W2765));
  INVX1 G5522 (.I(W499), .ZN(W4726));
  INVX1 G5523 (.I(I773), .ZN(W624));
  INVX1 G5524 (.I(I165), .ZN(O1031));
  INVX1 G5525 (.I(W2979), .ZN(W4015));
  INVX1 G5526 (.I(W4245), .ZN(O1039));
  INVX1 G5527 (.I(W1492), .ZN(O281));
  INVX1 G5528 (.I(W1340), .ZN(W4732));
  INVX1 G5529 (.I(W1942), .ZN(O1041));
  INVX1 G5530 (.I(I322), .ZN(W2760));
  INVX1 G5531 (.I(I502), .ZN(W4014));
  INVX1 G5532 (.I(I848), .ZN(W620));
  INVX1 G5533 (.I(I485), .ZN(W4019));
  INVX1 G5534 (.I(W3641), .ZN(O1019));
  INVX1 G5535 (.I(W197), .ZN(W2775));
  INVX1 G5536 (.I(W110), .ZN(W631));
  INVX1 G5537 (.I(W1085), .ZN(W2773));
  INVX1 G5538 (.I(W285), .ZN(O1022));
  INVX1 G5539 (.I(W65), .ZN(W630));
  INVX1 G5540 (.I(I796), .ZN(W2772));
  INVX1 G5541 (.I(W2386), .ZN(W2771));
  INVX1 G5542 (.I(W258), .ZN(W847));
  INVX1 G5543 (.I(W4635), .ZN(O1026));
  INVX1 G5544 (.I(I446), .ZN(W1118));
  INVX1 G5545 (.I(W4458), .ZN(W4712));
  INVX1 G5546 (.I(I719), .ZN(W4713));
  INVX1 G5547 (.I(W1155), .ZN(O1028));
  INVX1 G5548 (.I(W1705), .ZN(W3201));
  INVX1 G5549 (.I(W190), .ZN(O1029));
  INVX1 G5550 (.I(W40), .ZN(O283));
  INVX1 G5551 (.I(I605), .ZN(W609));
  INVX1 G5552 (.I(I153), .ZN(W2744));
  INVX1 G5553 (.I(W464), .ZN(W1116));
  INVX1 G5554 (.I(W3924), .ZN(W4758));
  INVX1 G5555 (.I(W2104), .ZN(O1055));
  INVX1 G5556 (.I(W507), .ZN(W612));
  INVX1 G5557 (.I(W941), .ZN(W2742));
  INVX1 G5558 (.I(I229), .ZN(W610));
  INVX1 G5559 (.I(W116), .ZN(O275));
  INVX1 G5560 (.I(W406), .ZN(W2746));
  INVX1 G5561 (.I(W3722), .ZN(W4765));
  INVX1 G5562 (.I(W403), .ZN(W607));
  INVX1 G5563 (.I(I683), .ZN(W1271));
  INVX1 G5564 (.I(W242), .ZN(O274));
  INVX1 G5565 (.I(I919), .ZN(W605));
  INVX1 G5566 (.I(W521), .ZN(W604));
  INVX1 G5567 (.I(W3947), .ZN(W4006));
  INVX1 G5568 (.I(W582), .ZN(W1273));
  INVX1 G5569 (.I(W284), .ZN(O1049));
  INVX1 G5570 (.I(W1661), .ZN(O1045));
  INVX1 G5571 (.I(I977), .ZN(O279));
  INVX1 G5572 (.I(W1254), .ZN(W2755));
  INVX1 G5573 (.I(W2750), .ZN(W2754));
  INVX1 G5574 (.I(W1585), .ZN(W3203));
  INVX1 G5575 (.I(W2670), .ZN(O690));
  INVX1 G5576 (.I(I444), .ZN(W4744));
  INVX1 G5577 (.I(W168), .ZN(W4745));
  INVX1 G5578 (.I(W924), .ZN(W2776));
  INVX1 G5579 (.I(W63), .ZN(W2750));
  INVX1 G5580 (.I(W415), .ZN(O399));
  INVX1 G5581 (.I(W217), .ZN(W1269));
  INVX1 G5582 (.I(I991), .ZN(O1050));
  INVX1 G5583 (.I(W4094), .ZN(O1051));
  INVX1 G5584 (.I(I730), .ZN(W615));
  INVX1 G5585 (.I(W4629), .ZN(W4753));
  INVX1 G5586 (.I(W3912), .ZN(O991));
  INVX1 G5587 (.I(I528), .ZN(W842));
  INVX1 G5588 (.I(W3062), .ZN(W4037));
  INVX1 G5589 (.I(W1343), .ZN(O292));
  INVX1 G5590 (.I(I91), .ZN(W1251));
  INVX1 G5591 (.I(W137), .ZN(W4646));
  INVX1 G5592 (.I(W586), .ZN(W843));
  INVX1 G5593 (.I(I797), .ZN(W4648));
  INVX1 G5594 (.I(W1381), .ZN(O990));
  INVX1 G5595 (.I(W3444), .ZN(W4641));
  INVX1 G5596 (.I(W4008), .ZN(O992));
  INVX1 G5597 (.I(W36), .ZN(O701));
  INVX1 G5598 (.I(W72), .ZN(W645));
  INVX1 G5599 (.I(W3902), .ZN(W4655));
  INVX1 G5600 (.I(W2281), .ZN(W4656));
  INVX1 G5601 (.I(W11), .ZN(O700));
  INVX1 G5602 (.I(W3636), .ZN(W4032));
  INVX1 G5603 (.I(W277), .ZN(W1120));
  INVX1 G5604 (.I(I414), .ZN(W839));
  INVX1 G5605 (.I(W1963), .ZN(W4624));
  INVX1 G5606 (.I(I113), .ZN(W1242));
  INVX1 G5607 (.I(W286), .ZN(W3183));
  INVX1 G5608 (.I(W2149), .ZN(O298));
  INVX1 G5609 (.I(W3399), .ZN(W4628));
  INVX1 G5610 (.I(I834), .ZN(O57));
  INVX1 G5611 (.I(W1116), .ZN(W4044));
  INVX1 G5612 (.I(W437), .ZN(W2824));
  INVX1 G5613 (.I(W929), .ZN(W1255));
  INVX1 G5614 (.I(W2122), .ZN(W4042));
  INVX1 G5615 (.I(I166), .ZN(W2821));
  INVX1 G5616 (.I(I481), .ZN(W1125));
  INVX1 G5617 (.I(W74), .ZN(W1124));
  INVX1 G5618 (.I(W333), .ZN(W2818));
  INVX1 G5619 (.I(W1429), .ZN(W4638));
  INVX1 G5620 (.I(I60), .ZN(W1246));
  INVX1 G5621 (.I(W1289), .ZN(O287));
  INVX1 G5622 (.I(W866), .ZN(W4682));
  INVX1 G5623 (.I(W1489), .ZN(O1009));
  INVX1 G5624 (.I(I441), .ZN(W638));
  INVX1 G5625 (.I(W397), .ZN(W637));
  INVX1 G5626 (.I(I216), .ZN(O20));
  INVX1 G5627 (.I(W2688), .ZN(W2785));
  INVX1 G5628 (.I(W4267), .ZN(O1012));
  INVX1 G5629 (.I(W2336), .ZN(W4689));
  INVX1 G5630 (.I(I407), .ZN(O1007));
  INVX1 G5631 (.I(I452), .ZN(W634));
  INVX1 G5632 (.I(W1702), .ZN(W2783));
  INVX1 G5633 (.I(W2404), .ZN(W2782));
  INVX1 G5634 (.I(W185), .ZN(O286));
  INVX1 G5635 (.I(W1745), .ZN(W2779));
  INVX1 G5636 (.I(W6), .ZN(W3198));
  INVX1 G5637 (.I(W218), .ZN(W4697));
  INVX1 G5638 (.I(W274), .ZN(O1018));
  INVX1 G5639 (.I(W2161), .ZN(O1001));
  INVX1 G5640 (.I(W13), .ZN(O290));
  INVX1 G5641 (.I(W1587), .ZN(W2798));
  INVX1 G5642 (.I(I578), .ZN(W3192));
  INVX1 G5643 (.I(W2465), .ZN(O997));
  INVX1 G5644 (.I(W1226), .ZN(W1256));
  INVX1 G5645 (.I(W2161), .ZN(W3194));
  INVX1 G5646 (.I(I94), .ZN(W1257));
  INVX1 G5647 (.I(W1407), .ZN(O696));
  INVX1 G5648 (.I(I18), .ZN(W2909));
  INVX1 G5649 (.I(W3575), .ZN(O1002));
  INVX1 G5650 (.I(W1755), .ZN(O289));
  INVX1 G5651 (.I(W2501), .ZN(W4024));
  INVX1 G5652 (.I(W1805), .ZN(W2788));
  INVX1 G5653 (.I(W3457), .ZN(W4677));
  INVX1 G5654 (.I(I641), .ZN(O1005));
  INVX1 G5655 (.I(I968), .ZN(W4023));
  INVX1 G5656 (.I(W239), .ZN(W3038));
  INVX1 G5657 (.I(W3337), .ZN(O749));
  INVX1 G5658 (.I(I743), .ZN(W1170));
  INVX1 G5659 (.I(I808), .ZN(W767));
  INVX1 G5660 (.I(W146), .ZN(W4271));
  INVX1 G5661 (.I(I658), .ZN(W4272));
  INVX1 G5662 (.I(W2957), .ZN(W3127));
  INVX1 G5663 (.I(I339), .ZN(W4135));
  INVX1 G5664 (.I(W599), .ZN(W4275));
  INVX1 G5665 (.I(I660), .ZN(O351));
  INVX1 G5666 (.I(W3042), .ZN(W4277));
  INVX1 G5667 (.I(W4175), .ZN(O813));
  INVX1 G5668 (.I(W207), .ZN(W4279));
  INVX1 G5669 (.I(I745), .ZN(W766));
  INVX1 G5670 (.I(W878), .ZN(W3037));
  INVX1 G5671 (.I(W934), .ZN(W1171));
  INVX1 G5672 (.I(W1402), .ZN(W3035));
  INVX1 G5673 (.I(W356), .ZN(W1172));
  INVX1 G5674 (.I(W406), .ZN(W4257));
  INVX1 G5675 (.I(W304), .ZN(W3054));
  INVX1 G5676 (.I(I310), .ZN(W4249));
  INVX1 G5677 (.I(W569), .ZN(O354));
  INVX1 G5678 (.I(W863), .ZN(W4251));
  INVX1 G5679 (.I(W231), .ZN(W773));
  INVX1 G5680 (.I(W2597), .ZN(W3051));
  INVX1 G5681 (.I(W3413), .ZN(W4255));
  INVX1 G5682 (.I(W2516), .ZN(W4256));
  INVX1 G5683 (.I(I892), .ZN(W3128));
  INVX1 G5684 (.I(W1676), .ZN(W4258));
  INVX1 G5685 (.I(W658), .ZN(W4259));
  INVX1 G5686 (.I(W292), .ZN(O47));
  INVX1 G5687 (.I(W1620), .ZN(W4140));
  INVX1 G5688 (.I(W2900), .ZN(W3125));
  INVX1 G5689 (.I(W682), .ZN(W3046));
  INVX1 G5690 (.I(I134), .ZN(W3044));
  INVX1 G5691 (.I(W749), .ZN(W4266));
  INVX1 G5692 (.I(W3707), .ZN(W4312));
  INVX1 G5693 (.I(W3084), .ZN(W4303));
  INVX1 G5694 (.I(I953), .ZN(W1180));
  INVX1 G5695 (.I(W730), .ZN(W1181));
  INVX1 G5696 (.I(W1118), .ZN(O50));
  INVX1 G5697 (.I(W524), .ZN(O821));
  INVX1 G5698 (.I(I820), .ZN(O746));
  INVX1 G5699 (.I(I843), .ZN(W1184));
  INVX1 G5700 (.I(W2456), .ZN(O824));
  INVX1 G5701 (.I(W58), .ZN(W807));
  INVX1 G5702 (.I(W712), .ZN(W809));
  INVX1 G5703 (.I(W1070), .ZN(O825));
  INVX1 G5704 (.I(I536), .ZN(W4315));
  INVX1 G5705 (.I(W2579), .ZN(W3014));
  INVX1 G5706 (.I(W1970), .ZN(W4124));
  INVX1 G5707 (.I(W1566), .ZN(W4319));
  INVX1 G5708 (.I(W2989), .ZN(O344));
  INVX1 G5709 (.I(W1991), .ZN(W4123));
  INVX1 G5710 (.I(W248), .ZN(W4294));
  INVX1 G5711 (.I(W1045), .ZN(W3129));
  INVX1 G5712 (.I(I584), .ZN(W805));
  INVX1 G5713 (.I(I454), .ZN(O49));
  INVX1 G5714 (.I(I160), .ZN(W762));
  INVX1 G5715 (.I(W2898), .ZN(W3130));
  INVX1 G5716 (.I(W101), .ZN(W4291));
  INVX1 G5717 (.I(W3287), .ZN(W4292));
  INVX1 G5718 (.I(I267), .ZN(W760));
  INVX1 G5719 (.I(I485), .ZN(O752));
  INVX1 G5720 (.I(W963), .ZN(W1177));
  INVX1 G5721 (.I(W657), .ZN(W759));
  INVX1 G5722 (.I(W3281), .ZN(W4297));
  INVX1 G5723 (.I(W443), .ZN(W3131));
  INVX1 G5724 (.I(I873), .ZN(W4299));
  INVX1 G5725 (.I(I404), .ZN(W3024));
  INVX1 G5726 (.I(W751), .ZN(W758));
  INVX1 G5727 (.I(W1982), .ZN(O369));
  INVX1 G5728 (.I(I0), .ZN(W789));
  INVX1 G5729 (.I(I974), .ZN(O363));
  INVX1 G5730 (.I(W744), .ZN(W4187));
  INVX1 G5731 (.I(W1012), .ZN(W4188));
  INVX1 G5732 (.I(W3003), .ZN(O770));
  INVX1 G5733 (.I(I963), .ZN(W4190));
  INVX1 G5734 (.I(I849), .ZN(W796));
  INVX1 G5735 (.I(W242), .ZN(O772));
  INVX1 G5736 (.I(W3884), .ZN(W4162));
  INVX1 G5737 (.I(W779), .ZN(W4195));
  INVX1 G5738 (.I(W2953), .ZN(W3086));
  INVX1 G5739 (.I(W857), .ZN(O774));
  INVX1 G5740 (.I(W868), .ZN(W4198));
  INVX1 G5741 (.I(W3116), .ZN(O775));
  INVX1 G5742 (.I(W2558), .ZN(O361));
  INVX1 G5743 (.I(I464), .ZN(O27));
  INVX1 G5744 (.I(W425), .ZN(W4204));
  INVX1 G5745 (.I(W2009), .ZN(W3097));
  INVX1 G5746 (.I(W3742), .ZN(O764));
  INVX1 G5747 (.I(W2823), .ZN(W3102));
  INVX1 G5748 (.I(W919), .ZN(W1148));
  INVX1 G5749 (.I(I285), .ZN(W4171));
  INVX1 G5750 (.I(I753), .ZN(W1151));
  INVX1 G5751 (.I(I168), .ZN(W3099));
  INVX1 G5752 (.I(W170), .ZN(W3098));
  INVX1 G5753 (.I(W2471), .ZN(W4175));
  INVX1 G5754 (.I(W1732), .ZN(O359));
  INVX1 G5755 (.I(W2586), .ZN(O366));
  INVX1 G5756 (.I(W3952), .ZN(W4164));
  INVX1 G5757 (.I(W2967), .ZN(W4179));
  INVX1 G5758 (.I(W230), .ZN(W4180));
  INVX1 G5759 (.I(I274), .ZN(O767));
  INVX1 G5760 (.I(W2723), .ZN(O762));
  INVX1 G5761 (.I(W521), .ZN(W1153));
  INVX1 G5762 (.I(W866), .ZN(W1142));
  INVX1 G5763 (.I(W921), .ZN(O794));
  INVX1 G5764 (.I(I546), .ZN(W4227));
  INVX1 G5765 (.I(W1700), .ZN(O795));
  INVX1 G5766 (.I(W272), .ZN(W1144));
  INVX1 G5767 (.I(W536), .ZN(O798));
  INVX1 G5768 (.I(W2519), .ZN(W3068));
  INVX1 G5769 (.I(W2247), .ZN(W4233));
  INVX1 G5770 (.I(W165), .ZN(W4234));
  INVX1 G5771 (.I(W976), .ZN(O755));
  INVX1 G5772 (.I(W23), .ZN(O48));
  INVX1 G5773 (.I(W957), .ZN(O801));
  INVX1 G5774 (.I(I544), .ZN(W800));
  INVX1 G5775 (.I(W3542), .ZN(W4241));
  INVX1 G5776 (.I(W2765), .ZN(W3061));
  INVX1 G5777 (.I(W1832), .ZN(W3059));
  INVX1 G5778 (.I(W1559), .ZN(W3058));
  INVX1 G5779 (.I(W2073), .ZN(W3057));
  INVX1 G5780 (.I(W1720), .ZN(O785));
  INVX1 G5781 (.I(W1330), .ZN(W4206));
  INVX1 G5782 (.I(W1099), .ZN(O780));
  INVX1 G5783 (.I(I608), .ZN(O781));
  INVX1 G5784 (.I(W1768), .ZN(W4209));
  INVX1 G5785 (.I(W2158), .ZN(O782));
  INVX1 G5786 (.I(I592), .ZN(W785));
  INVX1 G5787 (.I(W126), .ZN(W4212));
  INVX1 G5788 (.I(I915), .ZN(O759));
  INVX1 G5789 (.I(W878), .ZN(W3008));
  INVX1 G5790 (.I(W175), .ZN(W782));
  INVX1 G5791 (.I(I337), .ZN(W3079));
  INVX1 G5792 (.I(W1326), .ZN(O788));
  INVX1 G5793 (.I(W2899), .ZN(W3077));
  INVX1 G5794 (.I(I957), .ZN(W4221));
  INVX1 G5795 (.I(W2148), .ZN(O370));
  INVX1 G5796 (.I(I322), .ZN(W3075));
  INVX1 G5797 (.I(W2580), .ZN(O875));
  INVX1 G5798 (.I(W143), .ZN(O868));
  INVX1 G5799 (.I(I755), .ZN(O334));
  INVX1 G5800 (.I(W271), .ZN(O54));
  INVX1 G5801 (.I(W91), .ZN(W721));
  INVX1 G5802 (.I(I929), .ZN(W4092));
  INVX1 G5803 (.I(W269), .ZN(W3157));
  INVX1 G5804 (.I(W4327), .ZN(O874));
  INVX1 G5805 (.I(W564), .ZN(W4427));
  INVX1 G5806 (.I(I122), .ZN(W2950));
  INVX1 G5807 (.I(W2051), .ZN(O385));
  INVX1 G5808 (.I(W1273), .ZN(W2939));
  INVX1 G5809 (.I(W4161), .ZN(W4431));
  INVX1 G5810 (.I(W1072), .ZN(O876));
  INVX1 G5811 (.I(W892), .ZN(O877));
  INVX1 G5812 (.I(W2228), .ZN(O331));
  INVX1 G5813 (.I(W437), .ZN(W1210));
  INVX1 G5814 (.I(I162), .ZN(W2936));
  INVX1 G5815 (.I(W589), .ZN(O383));
  INVX1 G5816 (.I(W1946), .ZN(W3150));
  INVX1 G5817 (.I(I947), .ZN(W2960));
  INVX1 G5818 (.I(W3774), .ZN(W4098));
  INVX1 G5819 (.I(W3796), .ZN(W4402));
  INVX1 G5820 (.I(W2676), .ZN(O858));
  INVX1 G5821 (.I(W176), .ZN(O859));
  INVX1 G5822 (.I(W10), .ZN(W727));
  INVX1 G5823 (.I(W907), .ZN(W4406));
  INVX1 G5824 (.I(W2386), .ZN(O330));
  INVX1 G5825 (.I(I178), .ZN(W2957));
  INVX1 G5826 (.I(W2055), .ZN(W2956));
  INVX1 G5827 (.I(W59), .ZN(W4410));
  INVX1 G5828 (.I(I340), .ZN(W817));
  INVX1 G5829 (.I(W1839), .ZN(W2954));
  INVX1 G5830 (.I(W1911), .ZN(W2953));
  INVX1 G5831 (.I(W735), .ZN(W1202));
  INVX1 G5832 (.I(I671), .ZN(W725));
  INVX1 G5833 (.I(W531), .ZN(W825));
  INVX1 G5834 (.I(W1999), .ZN(W2919));
  INVX1 G5835 (.I(W2907), .ZN(O324));
  INVX1 G5836 (.I(W765), .ZN(W2917));
  INVX1 G5837 (.I(W2024), .ZN(O894));
  INVX1 G5838 (.I(W290), .ZN(W710));
  INVX1 G5839 (.I(W2319), .ZN(W2916));
  INVX1 G5840 (.I(W1080), .ZN(W4082));
  INVX1 G5841 (.I(W484), .ZN(W2914));
  INVX1 G5842 (.I(W508), .ZN(W1215));
  INVX1 G5843 (.I(I827), .ZN(W709));
  INVX1 G5844 (.I(I384), .ZN(W708));
  INVX1 G5845 (.I(W2135), .ZN(W2912));
  INVX1 G5846 (.I(I269), .ZN(O901));
  INVX1 G5847 (.I(I426), .ZN(W706));
  INVX1 G5848 (.I(W1598), .ZN(O903));
  INVX1 G5849 (.I(W533), .ZN(W2910));
  INVX1 G5850 (.I(W679), .ZN(W705));
  INVX1 G5851 (.I(I615), .ZN(W2925));
  INVX1 G5852 (.I(W645), .ZN(W1211));
  INVX1 G5853 (.I(I620), .ZN(W1212));
  INVX1 G5854 (.I(W3036), .ZN(O728));
  INVX1 G5855 (.I(W3229), .ZN(W4441));
  INVX1 G5856 (.I(W1587), .ZN(O882));
  INVX1 G5857 (.I(W1668), .ZN(W3159));
  INVX1 G5858 (.I(W826), .ZN(O327));
  INVX1 G5859 (.I(W2397), .ZN(W4447));
  INVX1 G5860 (.I(W682), .ZN(W728));
  INVX1 G5861 (.I(W2268), .ZN(O887));
  INVX1 G5862 (.I(W2140), .ZN(W2924));
  INVX1 G5863 (.I(W2421), .ZN(O888));
  INVX1 G5864 (.I(I16), .ZN(W716));
  INVX1 G5865 (.I(W957), .ZN(W4085));
  INVX1 G5866 (.I(W704), .ZN(W823));
  INVX1 G5867 (.I(W1559), .ZN(W3162));
  INVX1 G5868 (.I(I628), .ZN(W4352));
  INVX1 G5869 (.I(I543), .ZN(W747));
  INVX1 G5870 (.I(I444), .ZN(W1134));
  INVX1 G5871 (.I(W967), .ZN(W2992));
  INVX1 G5872 (.I(I707), .ZN(O839));
  INVX1 G5873 (.I(W1870), .ZN(W4113));
  INVX1 G5874 (.I(W1819), .ZN(O339));
  INVX1 G5875 (.I(W2375), .ZN(O841));
  INVX1 G5876 (.I(W643), .ZN(O842));
  INVX1 G5877 (.I(W3), .ZN(W2995));
  INVX1 G5878 (.I(W1139), .ZN(W4353));
  INVX1 G5879 (.I(W210), .ZN(W2988));
  INVX1 G5880 (.I(W606), .ZN(W4355));
  INVX1 G5881 (.I(W1489), .ZN(W2987));
  INVX1 G5882 (.I(I12), .ZN(O24));
  INVX1 G5883 (.I(I609), .ZN(O844));
  INVX1 G5884 (.I(I350), .ZN(W1193));
  INVX1 G5885 (.I(W4065), .ZN(O845));
  INVX1 G5886 (.I(W687), .ZN(W751));
  INVX1 G5887 (.I(W142), .ZN(W1136));
  INVX1 G5888 (.I(W1481), .ZN(O829));
  INVX1 G5889 (.I(W1569), .ZN(W3138));
  INVX1 G5890 (.I(W4253), .ZN(W4327));
  INVX1 G5891 (.I(W174), .ZN(O831));
  INVX1 G5892 (.I(W41), .ZN(W3004));
  INVX1 G5893 (.I(W391), .ZN(W4330));
  INVX1 G5894 (.I(W989), .ZN(W4331));
  INVX1 G5895 (.I(W2471), .ZN(O338));
  INVX1 G5896 (.I(W3127), .ZN(W4333));
  INVX1 G5897 (.I(W3316), .ZN(W4334));
  INVX1 G5898 (.I(I970), .ZN(O742));
  INVX1 G5899 (.I(I587), .ZN(W1190));
  INVX1 G5900 (.I(W2794), .ZN(O341));
  INVX1 G5901 (.I(W2446), .ZN(O740));
  INVX1 G5902 (.I(I892), .ZN(W1191));
  INVX1 G5903 (.I(I696), .ZN(W814));
  INVX1 G5904 (.I(W74), .ZN(W4379));
  INVX1 G5905 (.I(W1621), .ZN(O736));
  INVX1 G5906 (.I(W2694), .ZN(W2972));
  INVX1 G5907 (.I(W401), .ZN(O379));
  INVX1 G5908 (.I(W1459), .ZN(W4104));
  INVX1 G5909 (.I(W1255), .ZN(O852));
  INVX1 G5910 (.I(W76), .ZN(W2967));
  INVX1 G5911 (.I(W320), .ZN(O336));
  INVX1 G5912 (.I(W290), .ZN(O737));
  INVX1 G5913 (.I(W2699), .ZN(O382));
  INVX1 G5914 (.I(W2014), .ZN(O855));
  INVX1 G5915 (.I(W804), .ZN(W815));
  INVX1 G5916 (.I(W710), .ZN(W4393));
  INVX1 G5917 (.I(W2643), .ZN(O335));
  INVX1 G5918 (.I(W2721), .ZN(W4395));
  INVX1 G5919 (.I(W2494), .ZN(W4396));
  INVX1 G5920 (.I(I339), .ZN(W4397));
  INVX1 G5921 (.I(W323), .ZN(O738));
  INVX1 G5922 (.I(I261), .ZN(W1132));
  INVX1 G5923 (.I(W2190), .ZN(W4111));
  INVX1 G5924 (.I(W369), .ZN(W740));
  INVX1 G5925 (.I(W981), .ZN(W1194));
  INVX1 G5926 (.I(W3205), .ZN(W4366));
  INVX1 G5927 (.I(I871), .ZN(W4367));
  INVX1 G5928 (.I(W605), .ZN(W2981));
  INVX1 G5929 (.I(I305), .ZN(W4369));
  INVX1 G5930 (.I(W1954), .ZN(O1065));
  INVX1 G5931 (.I(W2661), .ZN(W2979));
  INVX1 G5932 (.I(W1444), .ZN(W2978));
  INVX1 G5933 (.I(W1368), .ZN(W3144));
  INVX1 G5934 (.I(W214), .ZN(W2975));
  INVX1 G5935 (.I(W4157), .ZN(O850));
  INVX1 G5936 (.I(W4284), .ZN(W4376));
  INVX1 G5937 (.I(W1291), .ZN(W4377));
  INVX1 G5938 (.I(W3353), .ZN(W5175));
  INVX1 G5939 (.I(I793), .ZN(W3894));
  INVX1 G5940 (.I(W3107), .ZN(W5168));
  INVX1 G5941 (.I(I57), .ZN(O1317));
  INVX1 G5942 (.I(W3389), .ZN(O637));
  INVX1 G5943 (.I(I222), .ZN(O1319));
  INVX1 G5944 (.I(I616), .ZN(O1320));
  INVX1 G5945 (.I(W1273), .ZN(W2492));
  INVX1 G5946 (.I(W183), .ZN(W893));
  INVX1 G5947 (.I(W5113), .ZN(O1315));
  INVX1 G5948 (.I(I934), .ZN(W467));
  INVX1 G5949 (.I(W4085), .ZN(O1324));
  INVX1 G5950 (.I(W767), .ZN(O1325));
  INVX1 G5951 (.I(W1697), .ZN(W5180));
  INVX1 G5952 (.I(I930), .ZN(W465));
  INVX1 G5953 (.I(W3398), .ZN(W5182));
  INVX1 G5954 (.I(W1104), .ZN(W3890));
  INVX1 G5955 (.I(W2701), .ZN(O635));
  INVX1 G5956 (.I(W1245), .ZN(W2501));
  INVX1 G5957 (.I(W3489), .ZN(W5149));
  INVX1 G5958 (.I(W1256), .ZN(O1302));
  INVX1 G5959 (.I(W32), .ZN(O1303));
  INVX1 G5960 (.I(I954), .ZN(W477));
  INVX1 G5961 (.I(I491), .ZN(O1305));
  INVX1 G5962 (.I(I332), .ZN(O222));
  INVX1 G5963 (.I(W1021), .ZN(O1307));
  INVX1 G5964 (.I(W2925), .ZN(W5156));
  INVX1 G5965 (.I(I320), .ZN(W3888));
  INVX1 G5966 (.I(I950), .ZN(W475));
  INVX1 G5967 (.I(I948), .ZN(W474));
  INVX1 G5968 (.I(W190), .ZN(W1342));
  INVX1 G5969 (.I(W2795), .ZN(W3897));
  INVX1 G5970 (.I(W3099), .ZN(W3264));
  INVX1 G5971 (.I(W970), .ZN(O1314));
  INVX1 G5972 (.I(W1129), .ZN(O417));
  INVX1 G5973 (.I(I811), .ZN(W2495));
  INVX1 G5974 (.I(W1927), .ZN(O1345));
  INVX1 G5975 (.I(W4906), .ZN(O1341));
  INVX1 G5976 (.I(W642), .ZN(W5204));
  INVX1 G5977 (.I(W2709), .ZN(O1342));
  INVX1 G5978 (.I(W2127), .ZN(O632));
  INVX1 G5979 (.I(W3603), .ZN(W3881));
  INVX1 G5980 (.I(I156), .ZN(W895));
  INVX1 G5981 (.I(W1216), .ZN(O1344));
  INVX1 G5982 (.I(I339), .ZN(W2469));
  INVX1 G5983 (.I(W3863), .ZN(W3883));
  INVX1 G5984 (.I(I816), .ZN(O631));
  INVX1 G5985 (.I(I696), .ZN(W2466));
  INVX1 G5986 (.I(W2213), .ZN(W5215));
  INVX1 G5987 (.I(W1492), .ZN(O1347));
  INVX1 G5988 (.I(W3264), .ZN(O1348));
  INVX1 G5989 (.I(I872), .ZN(W2465));
  INVX1 G5990 (.I(W1549), .ZN(W2464));
  INVX1 G5991 (.I(W4937), .ZN(O1350));
  INVX1 G5992 (.I(W2541), .ZN(W3269));
  INVX1 G5993 (.I(W2478), .ZN(W3887));
  INVX1 G5994 (.I(I912), .ZN(O1327));
  INVX1 G5995 (.I(W2004), .ZN(W2485));
  INVX1 G5996 (.I(W2371), .ZN(W2484));
  INVX1 G5997 (.I(W873), .ZN(W1350));
  INVX1 G5998 (.I(I721), .ZN(W3267));
  INVX1 G5999 (.I(W349), .ZN(W2481));
  INVX1 G6000 (.I(W1387), .ZN(O217));
  INVX1 G6001 (.I(W1584), .ZN(W5148));
  INVX1 G6002 (.I(W1885), .ZN(W2478));
  INVX1 G6003 (.I(W2609), .ZN(O1335));
  INVX1 G6004 (.I(I368), .ZN(W3270));
  INVX1 G6005 (.I(W4302), .ZN(O1337));
  INVX1 G6006 (.I(W2408), .ZN(W2476));
  INVX1 G6007 (.I(W684), .ZN(W2475));
  INVX1 G6008 (.I(W513), .ZN(W1352));
  INVX1 G6009 (.I(W2118), .ZN(O1269));
  INVX1 G6010 (.I(W1471), .ZN(O1262));
  INVX1 G6011 (.I(I996), .ZN(W498));
  INVX1 G6012 (.I(W428), .ZN(W2541));
  INVX1 G6013 (.I(W4749), .ZN(O1264));
  INVX1 G6014 (.I(I458), .ZN(W885));
  INVX1 G6015 (.I(W2410), .ZN(O643));
  INVX1 G6016 (.I(W1793), .ZN(W2538));
  INVX1 G6017 (.I(I338), .ZN(O642));
  INVX1 G6018 (.I(I728), .ZN(W884));
  INVX1 G6019 (.I(W1783), .ZN(W5100));
  INVX1 G6020 (.I(W1997), .ZN(W2535));
  INVX1 G6021 (.I(W3665), .ZN(O1271));
  INVX1 G6022 (.I(W160), .ZN(W2533));
  INVX1 G6023 (.I(W3275), .ZN(W3913));
  INVX1 G6024 (.I(W2835), .ZN(O1274));
  INVX1 G6025 (.I(W2215), .ZN(W3912));
  INVX1 G6026 (.I(W321), .ZN(W2530));
  INVX1 G6027 (.I(W373), .ZN(W1330));
  INVX1 G6028 (.I(W2059), .ZN(O647));
  INVX1 G6029 (.I(W1030), .ZN(W2551));
  INVX1 G6030 (.I(W72), .ZN(O646));
  INVX1 G6031 (.I(W1841), .ZN(W2548));
  INVX1 G6032 (.I(W791), .ZN(O231));
  INVX1 G6033 (.I(I517), .ZN(O1255));
  INVX1 G6034 (.I(I724), .ZN(W501));
  INVX1 G6035 (.I(W1889), .ZN(W5080));
  INVX1 G6036 (.I(W1517), .ZN(W2529));
  INVX1 G6037 (.I(I85), .ZN(O1258));
  INVX1 G6038 (.I(W4965), .ZN(O1259));
  INVX1 G6039 (.I(W423), .ZN(W5084));
  INVX1 G6040 (.I(W895), .ZN(W3921));
  INVX1 G6041 (.I(W1335), .ZN(O1260));
  INVX1 G6042 (.I(I874), .ZN(W883));
  INVX1 G6043 (.I(W3352), .ZN(O1261));
  INVX1 G6044 (.I(W4413), .ZN(O1297));
  INVX1 G6045 (.I(W2802), .ZN(O1290));
  INVX1 G6046 (.I(W4148), .ZN(O1292));
  INVX1 G6047 (.I(W4279), .ZN(O1293));
  INVX1 G6048 (.I(W1757), .ZN(O223));
  INVX1 G6049 (.I(W1662), .ZN(O1295));
  INVX1 G6050 (.I(W2334), .ZN(W5135));
  INVX1 G6051 (.I(W473), .ZN(W889));
  INVX1 G6052 (.I(I977), .ZN(W3903));
  INVX1 G6053 (.I(W810), .ZN(W1338));
  INVX1 G6054 (.I(W2552), .ZN(W5139));
  INVX1 G6055 (.I(I777), .ZN(W890));
  INVX1 G6056 (.I(W2914), .ZN(W3260));
  INVX1 G6057 (.I(W2535), .ZN(O416));
  INVX1 G6058 (.I(I960), .ZN(W480));
  INVX1 G6059 (.I(I958), .ZN(W479));
  INVX1 G6060 (.I(W4748), .ZN(O1300));
  INVX1 G6061 (.I(I525), .ZN(W3898));
  INVX1 G6062 (.I(W1722), .ZN(O224));
  INVX1 G6063 (.I(I984), .ZN(W492));
  INVX1 G6064 (.I(W3523), .ZN(W3911));
  INVX1 G6065 (.I(W3049), .ZN(W3257));
  INVX1 G6066 (.I(W964), .ZN(W2524));
  INVX1 G6067 (.I(W2380), .ZN(W3907));
  INVX1 G6068 (.I(I978), .ZN(W489));
  INVX1 G6069 (.I(I19), .ZN(W1334));
  INVX1 G6070 (.I(W941), .ZN(W1337));
  INVX1 G6071 (.I(W2002), .ZN(W3273));
  INVX1 G6072 (.I(W2671), .ZN(O640));
  INVX1 G6073 (.I(W1406), .ZN(W5122));
  INVX1 G6074 (.I(W4369), .ZN(O1286));
  INVX1 G6075 (.I(I488), .ZN(W2515));
  INVX1 G6076 (.I(W844), .ZN(W2514));
  INVX1 G6077 (.I(I970), .ZN(W485));
  INVX1 G6078 (.I(W3347), .ZN(W5127));
  INVX1 G6079 (.I(W2807), .ZN(W5327));
  INVX1 G6080 (.I(W156), .ZN(O424));
  INVX1 G6081 (.I(W3905), .ZN(O1421));
  INVX1 G6082 (.I(W3444), .ZN(O1422));
  INVX1 G6083 (.I(I195), .ZN(O1423));
  INVX1 G6084 (.I(W529), .ZN(W908));
  INVX1 G6085 (.I(W3748), .ZN(O1426));
  INVX1 G6086 (.I(I910), .ZN(O611));
  INVX1 G6087 (.I(I773), .ZN(O204));
  INVX1 G6088 (.I(I423), .ZN(W3848));
  INVX1 G6089 (.I(W2189), .ZN(O1428));
  INVX1 G6090 (.I(W178), .ZN(O35));
  INVX1 G6091 (.I(I731), .ZN(W1081));
  INVX1 G6092 (.I(I323), .ZN(O1431));
  INVX1 G6093 (.I(I354), .ZN(W1382));
  INVX1 G6094 (.I(W2714), .ZN(O765));
  INVX1 G6095 (.I(I822), .ZN(W411));
  INVX1 G6096 (.I(W663), .ZN(W910));
  INVX1 G6097 (.I(I836), .ZN(W418));
  INVX1 G6098 (.I(W1853), .ZN(W2410));
  INVX1 G6099 (.I(W1002), .ZN(O206));
  INVX1 G6100 (.I(I846), .ZN(W423));
  INVX1 G6101 (.I(I662), .ZN(W2407));
  INVX1 G6102 (.I(I844), .ZN(W422));
  INVX1 G6103 (.I(W571), .ZN(W905));
  INVX1 G6104 (.I(I840), .ZN(W420));
  INVX1 G6105 (.I(W1283), .ZN(W1372));
  INVX1 G6106 (.I(W2027), .ZN(O1436));
  INVX1 G6107 (.I(I834), .ZN(W417));
  INVX1 G6108 (.I(W135), .ZN(W2404));
  INVX1 G6109 (.I(I191), .ZN(W3852));
  INVX1 G6110 (.I(W1175), .ZN(O1412));
  INVX1 G6111 (.I(W76), .ZN(W1375));
  INVX1 G6112 (.I(I946), .ZN(O1415));
  INVX1 G6113 (.I(W4812), .ZN(W5314));
  INVX1 G6114 (.I(W832), .ZN(W1083));
  INVX1 G6115 (.I(W208), .ZN(O1455));
  INVX1 G6116 (.I(W1939), .ZN(O1449));
  INVX1 G6117 (.I(W555), .ZN(W2372));
  INVX1 G6118 (.I(W453), .ZN(W5357));
  INVX1 G6119 (.I(I137), .ZN(W1385));
  INVX1 G6120 (.I(W293), .ZN(W3834));
  INVX1 G6121 (.I(I806), .ZN(W403));
  INVX1 G6122 (.I(W2979), .ZN(O1454));
  INVX1 G6123 (.I(I804), .ZN(W402));
  INVX1 G6124 (.I(W2883), .ZN(W3297));
  INVX1 G6125 (.I(W2311), .ZN(O1456));
  INVX1 G6126 (.I(W2223), .ZN(O1457));
  INVX1 G6127 (.I(I802), .ZN(W401));
  INVX1 G6128 (.I(W2803), .ZN(O1459));
  INVX1 G6129 (.I(I693), .ZN(O201));
  INVX1 G6130 (.I(I800), .ZN(W400));
  INVX1 G6131 (.I(W60), .ZN(W2367));
  INVX1 G6132 (.I(W1704), .ZN(O200));
  INVX1 G6133 (.I(W2141), .ZN(W2379));
  INVX1 G6134 (.I(W1052), .ZN(W1080));
  INVX1 G6135 (.I(W1616), .ZN(W2381));
  INVX1 G6136 (.I(W1731), .ZN(W2380));
  INVX1 G6137 (.I(W1539), .ZN(O1439));
  INVX1 G6138 (.I(W1871), .ZN(O1440));
  INVX1 G6139 (.I(I570), .ZN(O1441));
  INVX1 G6140 (.I(W4362), .ZN(O1442));
  INVX1 G6141 (.I(I385), .ZN(W5345));
  INVX1 G6142 (.I(I117), .ZN(W2411));
  INVX1 G6143 (.I(I647), .ZN(W1383));
  INVX1 G6144 (.I(I185), .ZN(W2377));
  INVX1 G6145 (.I(W244), .ZN(W1079));
  INVX1 G6146 (.I(W3652), .ZN(O1446));
  INVX1 G6147 (.I(W235), .ZN(W2375));
  INVX1 G6148 (.I(W2936), .ZN(O1447));
  INVX1 G6149 (.I(W320), .ZN(W1384));
  INVX1 G6150 (.I(I665), .ZN(W1365));
  INVX1 G6151 (.I(W4527), .ZN(O1363));
  INVX1 G6152 (.I(W88), .ZN(O1364));
  INVX1 G6153 (.I(W1636), .ZN(O1365));
  INVX1 G6154 (.I(I878), .ZN(W1359));
  INVX1 G6155 (.I(W849), .ZN(O1367));
  INVX1 G6156 (.I(W1146), .ZN(W1361));
  INVX1 G6157 (.I(W918), .ZN(W2444));
  INVX1 G6158 (.I(W856), .ZN(W901));
  INVX1 G6159 (.I(I890), .ZN(W445));
  INVX1 G6160 (.I(W5101), .ZN(O1373));
  INVX1 G6161 (.I(W21), .ZN(W1366));
  INVX1 G6162 (.I(W591), .ZN(W2438));
  INVX1 G6163 (.I(I882), .ZN(W441));
  INVX1 G6164 (.I(I637), .ZN(W2436));
  INVX1 G6165 (.I(I496), .ZN(O212));
  INVX1 G6166 (.I(W884), .ZN(W2434));
  INVX1 G6167 (.I(W3454), .ZN(O623));
  INVX1 G6168 (.I(W3384), .ZN(O627));
  INVX1 G6169 (.I(W309), .ZN(O421));
  INVX1 G6170 (.I(W1779), .ZN(W5224));
  INVX1 G6171 (.I(W3583), .ZN(W3874));
  INVX1 G6172 (.I(W609), .ZN(W897));
  INVX1 G6173 (.I(W3599), .ZN(O628));
  INVX1 G6174 (.I(W868), .ZN(W2456));
  INVX1 G6175 (.I(W4052), .ZN(O1354));
  INVX1 G6176 (.I(I898), .ZN(W449));
  INVX1 G6177 (.I(W949), .ZN(W2432));
  INVX1 G6178 (.I(W45), .ZN(W3275));
  INVX1 G6179 (.I(W309), .ZN(W1088));
  INVX1 G6180 (.I(I896), .ZN(W448));
  INVX1 G6181 (.I(W3174), .ZN(O625));
  INVX1 G6182 (.I(W1869), .ZN(O1360));
  INVX1 G6183 (.I(W1527), .ZN(O216));
  INVX1 G6184 (.I(W151), .ZN(W1087));
  INVX1 G6185 (.I(W4073), .ZN(O1398));
  INVX1 G6186 (.I(W2293), .ZN(O1394));
  INVX1 G6187 (.I(W128), .ZN(W5280));
  INVX1 G6188 (.I(W711), .ZN(W2419));
  INVX1 G6189 (.I(W492), .ZN(O208));
  INVX1 G6190 (.I(W449), .ZN(W2417));
  INVX1 G6191 (.I(W1033), .ZN(O1396));
  INVX1 G6192 (.I(W697), .ZN(O207));
  INVX1 G6193 (.I(W2610), .ZN(O618));
  INVX1 G6194 (.I(I773), .ZN(W2420));
  INVX1 G6195 (.I(I100), .ZN(W2414));
  INVX1 G6196 (.I(I854), .ZN(W427));
  INVX1 G6197 (.I(I337), .ZN(W5290));
  INVX1 G6198 (.I(W2877), .ZN(O1400));
  INVX1 G6199 (.I(W205), .ZN(W2413));
  INVX1 G6200 (.I(W3750), .ZN(O1402));
  INVX1 G6201 (.I(I366), .ZN(O617));
  INVX1 G6202 (.I(I850), .ZN(W425));
  INVX1 G6203 (.I(W1988), .ZN(O620));
  INVX1 G6204 (.I(W1763), .ZN(W3860));
  INVX1 G6205 (.I(W544), .ZN(W1367));
  INVX1 G6206 (.I(W1740), .ZN(O209));
  INVX1 G6207 (.I(W5143), .ZN(O1384));
  INVX1 G6208 (.I(W605), .ZN(W2428));
  INVX1 G6209 (.I(W1717), .ZN(W2427));
  INVX1 G6210 (.I(W2302), .ZN(W3283));
  INVX1 G6211 (.I(I890), .ZN(W904));
  INVX1 G6212 (.I(I153), .ZN(O233));
  INVX1 G6213 (.I(I868), .ZN(W434));
  INVX1 G6214 (.I(W163), .ZN(O1390));
  INVX1 G6215 (.I(W2130), .ZN(W3286));
  INVX1 G6216 (.I(I866), .ZN(W433));
  INVX1 G6217 (.I(W2282), .ZN(W5275));
  INVX1 G6218 (.I(I864), .ZN(W432));
  INVX1 G6219 (.I(W4883), .ZN(O1392));
  INVX1 G6220 (.I(W1602), .ZN(O1128));
  INVX1 G6221 (.I(I890), .ZN(W3986));
  INVX1 G6222 (.I(I730), .ZN(O1124));
  INVX1 G6223 (.I(W2793), .ZN(W4868));
  INVX1 G6224 (.I(W1862), .ZN(W3985));
  INVX1 G6225 (.I(W403), .ZN(O16));
  INVX1 G6226 (.I(W1712), .ZN(O264));
  INVX1 G6227 (.I(W430), .ZN(W2684));
  INVX1 G6228 (.I(W4600), .ZN(O1127));
  INVX1 G6229 (.I(W4180), .ZN(W4865));
  INVX1 G6230 (.I(I121), .ZN(W1111));
  INVX1 G6231 (.I(W4662), .ZN(W4877));
  INVX1 G6232 (.I(I616), .ZN(W1290));
  INVX1 G6233 (.I(W1708), .ZN(W4880));
  INVX1 G6234 (.I(W1098), .ZN(O402));
  INVX1 G6235 (.I(I797), .ZN(W858));
  INVX1 G6236 (.I(W23), .ZN(W4883));
  INVX1 G6237 (.I(W3446), .ZN(O1131));
  INVX1 G6238 (.I(I390), .ZN(W4856));
  INVX1 G6239 (.I(I324), .ZN(W580));
  INVX1 G6240 (.I(W1067), .ZN(W3213));
  INVX1 G6241 (.I(W2744), .ZN(O1115));
  INVX1 G6242 (.I(W64), .ZN(W1286));
  INVX1 G6243 (.I(W3216), .ZN(W4852));
  INVX1 G6244 (.I(W461), .ZN(O1116));
  INVX1 G6245 (.I(W2492), .ZN(O1117));
  INVX1 G6246 (.I(I20), .ZN(W2693));
  INVX1 G6247 (.I(W2631), .ZN(O403));
  INVX1 G6248 (.I(I464), .ZN(W578));
  INVX1 G6249 (.I(W818), .ZN(W2692));
  INVX1 G6250 (.I(W68), .ZN(W4859));
  INVX1 G6251 (.I(W2451), .ZN(O266));
  INVX1 G6252 (.I(I746), .ZN(W4861));
  INVX1 G6253 (.I(W187), .ZN(W575));
  INVX1 G6254 (.I(I682), .ZN(O401));
  INVX1 G6255 (.I(W2041), .ZN(O265));
  INVX1 G6256 (.I(I147), .ZN(W1296));
  INVX1 G6257 (.I(I446), .ZN(O404));
  INVX1 G6258 (.I(W4299), .ZN(W4904));
  INVX1 G6259 (.I(I413), .ZN(W863));
  INVX1 G6260 (.I(W419), .ZN(W864));
  INVX1 G6261 (.I(I7), .ZN(W563));
  INVX1 G6262 (.I(W3359), .ZN(W4908));
  INVX1 G6263 (.I(I547), .ZN(W4909));
  INVX1 G6264 (.I(W59), .ZN(W2661));
  INVX1 G6265 (.I(W2229), .ZN(W4902));
  INVX1 G6266 (.I(W1474), .ZN(W2658));
  INVX1 G6267 (.I(W2010), .ZN(O1151));
  INVX1 G6268 (.I(W2552), .ZN(W4915));
  INVX1 G6269 (.I(I31), .ZN(W558));
  INVX1 G6270 (.I(W2815), .ZN(O1152));
  INVX1 G6271 (.I(W1552), .ZN(W3969));
  INVX1 G6272 (.I(W329), .ZN(W2656));
  INVX1 G6273 (.I(W2060), .ZN(W2655));
  INVX1 G6274 (.I(I84), .ZN(W3975));
  INVX1 G6275 (.I(I797), .ZN(W1292));
  INVX1 G6276 (.I(W727), .ZN(W3221));
  INVX1 G6277 (.I(W2958), .ZN(O1135));
  INVX1 G6278 (.I(I147), .ZN(W566));
  INVX1 G6279 (.I(W679), .ZN(W2672));
  INVX1 G6280 (.I(W1655), .ZN(W3225));
  INVX1 G6281 (.I(W479), .ZN(W2670));
  INVX1 G6282 (.I(W1280), .ZN(W3976));
  INVX1 G6283 (.I(W385), .ZN(W581));
  INVX1 G6284 (.I(W1885), .ZN(W4895));
  INVX1 G6285 (.I(W2048), .ZN(O258));
  INVX1 G6286 (.I(W4019), .ZN(W4897));
  INVX1 G6287 (.I(I858), .ZN(O31));
  INVX1 G6288 (.I(W2961), .ZN(O1141));
  INVX1 G6289 (.I(W3933), .ZN(O1142));
  INVX1 G6290 (.I(W2487), .ZN(W2665));
  INVX1 G6291 (.I(W932), .ZN(W2723));
  INVX1 G6292 (.I(I23), .ZN(W852));
  INVX1 G6293 (.I(W1376), .ZN(O271));
  INVX1 G6294 (.I(W351), .ZN(W2727));
  INVX1 G6295 (.I(I70), .ZN(O1080));
  INVX1 G6296 (.I(I175), .ZN(W4001));
  INVX1 G6297 (.I(W2522), .ZN(W2725));
  INVX1 G6298 (.I(W230), .ZN(W2724));
  INVX1 G6299 (.I(W3832), .ZN(O1082));
  INVX1 G6300 (.I(W168), .ZN(W4791));
  INVX1 G6301 (.I(W1), .ZN(W593));
  INVX1 G6302 (.I(W2845), .ZN(O1083));
  INVX1 G6303 (.I(W1790), .ZN(W4803));
  INVX1 G6304 (.I(W4343), .ZN(O1084));
  INVX1 G6305 (.I(W351), .ZN(O1085));
  INVX1 G6306 (.I(W3519), .ZN(W4000));
  INVX1 G6307 (.I(W3820), .ZN(W3999));
  INVX1 G6308 (.I(W1183), .ZN(W1279));
  INVX1 G6309 (.I(W35), .ZN(W597));
  INVX1 G6310 (.I(W525), .ZN(O18));
  INVX1 G6311 (.I(W2575), .ZN(O1067));
  INVX1 G6312 (.I(I294), .ZN(W601));
  INVX1 G6313 (.I(I595), .ZN(W600));
  INVX1 G6314 (.I(W3350), .ZN(O1070));
  INVX1 G6315 (.I(I247), .ZN(W599));
  INVX1 G6316 (.I(I596), .ZN(W851));
  INVX1 G6317 (.I(W2262), .ZN(O1072));
  INVX1 G6318 (.I(W2153), .ZN(O687));
  INVX1 G6319 (.I(I388), .ZN(W1274));
  INVX1 G6320 (.I(W3403), .ZN(W4004));
  INVX1 G6321 (.I(W4399), .ZN(W4786));
  INVX1 G6322 (.I(W2872), .ZN(W4787));
  INVX1 G6323 (.I(W2723), .ZN(O272));
  INVX1 G6324 (.I(W926), .ZN(W1275));
  INVX1 G6325 (.I(W213), .ZN(W3208));
  INVX1 G6326 (.I(W4272), .ZN(O1107));
  INVX1 G6327 (.I(W2760), .ZN(O1100));
  INVX1 G6328 (.I(W222), .ZN(W585));
  INVX1 G6329 (.I(I705), .ZN(O58));
  INVX1 G6330 (.I(W1156), .ZN(O1102));
  INVX1 G6331 (.I(I5), .ZN(W3211));
  INVX1 G6332 (.I(W141), .ZN(W583));
  INVX1 G6333 (.I(W3104), .ZN(O1105));
  INVX1 G6334 (.I(I368), .ZN(O1106));
  INVX1 G6335 (.I(W966), .ZN(W1284));
  INVX1 G6336 (.I(W3784), .ZN(O680));
  INVX1 G6337 (.I(W3726), .ZN(W4840));
  INVX1 G6338 (.I(I412), .ZN(O1108));
  INVX1 G6339 (.I(W3707), .ZN(O1109));
  INVX1 G6340 (.I(W1894), .ZN(O267));
  INVX1 G6341 (.I(W102), .ZN(W2697));
  INVX1 G6342 (.I(W1500), .ZN(W2696));
  INVX1 G6343 (.I(W4239), .ZN(O1113));
  INVX1 G6344 (.I(W2902), .ZN(O683));
  INVX1 G6345 (.I(W600), .ZN(W2718));
  INVX1 G6346 (.I(W1668), .ZN(W4812));
  INVX1 G6347 (.I(W2467), .ZN(W2715));
  INVX1 G6348 (.I(I540), .ZN(W2713));
  INVX1 G6349 (.I(I464), .ZN(W2712));
  INVX1 G6350 (.I(I875), .ZN(O685));
  INVX1 G6351 (.I(W4203), .ZN(O1092));
  INVX1 G6352 (.I(W2744), .ZN(O684));
  INVX1 G6353 (.I(W706), .ZN(W865));
  INVX1 G6354 (.I(W3111), .ZN(O1095));
  INVX1 G6355 (.I(W2750), .ZN(O682));
  INVX1 G6356 (.I(W1423), .ZN(O1098));
  INVX1 G6357 (.I(W764), .ZN(W2705));
  INVX1 G6358 (.I(W2356), .ZN(O1099));
  INVX1 G6359 (.I(W439), .ZN(W2704));
  INVX1 G6360 (.I(I780), .ZN(W586));
  INVX1 G6361 (.I(W1043), .ZN(W1320));
  INVX1 G6362 (.I(W2766), .ZN(O1210));
  INVX1 G6363 (.I(W515), .ZN(W2590));
  INVX1 G6364 (.I(W2306), .ZN(W2589));
  INVX1 G6365 (.I(W2979), .ZN(W3942));
  INVX1 G6366 (.I(I940), .ZN(O239));
  INVX1 G6367 (.I(W1210), .ZN(W1318));
  INVX1 G6368 (.I(W349), .ZN(W2583));
  INVX1 G6369 (.I(W3567), .ZN(O657));
  INVX1 G6370 (.I(I614), .ZN(W1316));
  INVX1 G6371 (.I(I890), .ZN(O1221));
  INVX1 G6372 (.I(W2305), .ZN(W2578));
  INVX1 G6373 (.I(I409), .ZN(W2577));
  INVX1 G6374 (.I(W2194), .ZN(W5029));
  INVX1 G6375 (.I(I74), .ZN(W518));
  INVX1 G6376 (.I(W565), .ZN(W875));
  INVX1 G6377 (.I(I673), .ZN(W3937));
  INVX1 G6378 (.I(I145), .ZN(W516));
  INVX1 G6379 (.I(W2228), .ZN(W2598));
  INVX1 G6380 (.I(I977), .ZN(O1203));
  INVX1 G6381 (.I(I136), .ZN(O409));
  INVX1 G6382 (.I(W161), .ZN(W1313));
  INVX1 G6383 (.I(W1399), .ZN(O1204));
  INVX1 G6384 (.I(W735), .ZN(W871));
  INVX1 G6385 (.I(W353), .ZN(W1314));
  INVX1 G6386 (.I(W649), .ZN(W5001));
  INVX1 G6387 (.I(W331), .ZN(W5002));
  INVX1 G6388 (.I(W3381), .ZN(O1225));
  INVX1 G6389 (.I(W801), .ZN(W1104));
  INVX1 G6390 (.I(W477), .ZN(W1103));
  INVX1 G6391 (.I(W398), .ZN(W528));
  INVX1 G6392 (.I(I992), .ZN(O241));
  INVX1 G6393 (.I(W1394), .ZN(W5009));
  INVX1 G6394 (.I(W336), .ZN(W5010));
  INVX1 G6395 (.I(W838), .ZN(W2593));
  INVX1 G6396 (.I(I710), .ZN(W2592));
  INVX1 G6397 (.I(W243), .ZN(W2558));
  INVX1 G6398 (.I(W1105), .ZN(O1240));
  INVX1 G6399 (.I(W1906), .ZN(O1241));
  INVX1 G6400 (.I(W4880), .ZN(W5055));
  INVX1 G6401 (.I(W443), .ZN(W879));
  INVX1 G6402 (.I(W3711), .ZN(W5057));
  INVX1 G6403 (.I(I592), .ZN(W1097));
  INVX1 G6404 (.I(W747), .ZN(O650));
  INVX1 G6405 (.I(W4780), .ZN(O1244));
  INVX1 G6406 (.I(I57), .ZN(W1099));
  INVX1 G6407 (.I(W570), .ZN(W1328));
  INVX1 G6408 (.I(I0), .ZN(W0));
  INVX1 G6409 (.I(W3080), .ZN(W5066));
  INVX1 G6410 (.I(I406), .ZN(W3924));
  INVX1 G6411 (.I(W4281), .ZN(O1249));
  INVX1 G6412 (.I(W3818), .ZN(O1250));
  INVX1 G6413 (.I(W78), .ZN(W506));
  INVX1 G6414 (.I(W3461), .ZN(O1252));
  INVX1 G6415 (.I(W3064), .ZN(O1233));
  INVX1 G6416 (.I(W449), .ZN(W3936));
  INVX1 G6417 (.I(W1277), .ZN(W1325));
  INVX1 G6418 (.I(W2045), .ZN(O1228));
  INVX1 G6419 (.I(W2413), .ZN(O1229));
  INVX1 G6420 (.I(W841), .ZN(W876));
  INVX1 G6421 (.I(W286), .ZN(O14));
  INVX1 G6422 (.I(W819), .ZN(W2569));
  INVX1 G6423 (.I(W3809), .ZN(W5043));
  INVX1 G6424 (.I(I536), .ZN(O1202));
  INVX1 G6425 (.I(I848), .ZN(W2568));
  INVX1 G6426 (.I(W125), .ZN(O43));
  INVX1 G6427 (.I(I708), .ZN(W2566));
  INVX1 G6428 (.I(W268), .ZN(W878));
  INVX1 G6429 (.I(W4996), .ZN(W5049));
  INVX1 G6430 (.I(I210), .ZN(W2564));
  INVX1 G6431 (.I(I347), .ZN(W510));
  INVX1 G6432 (.I(W101), .ZN(W868));
  INVX1 G6433 (.I(W2303), .ZN(O1165));
  INVX1 G6434 (.I(W2201), .ZN(W2635));
  INVX1 G6435 (.I(W3918), .ZN(O668));
  INVX1 G6436 (.I(W536), .ZN(O1168));
  INVX1 G6437 (.I(W682), .ZN(W4945));
  INVX1 G6438 (.I(W4352), .ZN(O1169));
  INVX1 G6439 (.I(W4780), .ZN(O1170));
  INVX1 G6440 (.I(W886), .ZN(W2633));
  INVX1 G6441 (.I(W891), .ZN(O59));
  INVX1 G6442 (.I(I206), .ZN(O1172));
  INVX1 G6443 (.I(I962), .ZN(O1173));
  INVX1 G6444 (.I(W740), .ZN(O60));
  INVX1 G6445 (.I(W109), .ZN(W4953));
  INVX1 G6446 (.I(I6), .ZN(W549));
  INVX1 G6447 (.I(W3932), .ZN(O1176));
  INVX1 G6448 (.I(W3442), .ZN(O1177));
  INVX1 G6449 (.I(W771), .ZN(W2629));
  INVX1 G6450 (.I(W2221), .ZN(O1161));
  INVX1 G6451 (.I(W1267), .ZN(W2653));
  INVX1 G6452 (.I(I564), .ZN(W1298));
  INVX1 G6453 (.I(W2025), .ZN(W3967));
  INVX1 G6454 (.I(W1358), .ZN(W2647));
  INVX1 G6455 (.I(I338), .ZN(W2645));
  INVX1 G6456 (.I(I808), .ZN(O251));
  INVX1 G6457 (.I(W1377), .ZN(O1159));
  INVX1 G6458 (.I(W1215), .ZN(O1160));
  INVX1 G6459 (.I(W323), .ZN(W1307));
  INVX1 G6460 (.I(W4560), .ZN(O1162));
  INVX1 G6461 (.I(W2015), .ZN(W2642));
  INVX1 G6462 (.I(W970), .ZN(W1303));
  INVX1 G6463 (.I(W142), .ZN(W3964));
  INVX1 G6464 (.I(I261), .ZN(W3231));
  INVX1 G6465 (.I(W222), .ZN(W552));
  INVX1 G6466 (.I(W3480), .ZN(O669));
  INVX1 G6467 (.I(W33), .ZN(W537));
  INVX1 G6468 (.I(W2868), .ZN(O408));
  INVX1 G6469 (.I(W1657), .ZN(O664));
  INVX1 G6470 (.I(W634), .ZN(W3952));
  INVX1 G6471 (.I(W72), .ZN(W540));
  INVX1 G6472 (.I(W2602), .ZN(W2610));
  INVX1 G6473 (.I(W2354), .ZN(W2609));
  INVX1 G6474 (.I(W2343), .ZN(W2608));
  INVX1 G6475 (.I(W3360), .ZN(O663));
  INVX1 G6476 (.I(W2015), .ZN(O1188));
  INVX1 G6477 (.I(W3711), .ZN(W4986));
  INVX1 G6478 (.I(W1634), .ZN(W3950));
  INVX1 G6479 (.I(I217), .ZN(O62));
  INVX1 G6480 (.I(W865), .ZN(O244));
  INVX1 G6481 (.I(I382), .ZN(O15));
  INVX1 G6482 (.I(W1670), .ZN(O1199));
  INVX1 G6483 (.I(I626), .ZN(W870));
  INVX1 G6484 (.I(W1427), .ZN(O1201));
  INVX1 G6485 (.I(W1796), .ZN(O1184));
  INVX1 G6486 (.I(W4597), .ZN(W4959));
  INVX1 G6487 (.I(W1539), .ZN(O1180));
  INVX1 G6488 (.I(W1127), .ZN(W2627));
  INVX1 G6489 (.I(I814), .ZN(W1308));
  INVX1 G6490 (.I(W170), .ZN(W869));
  INVX1 G6491 (.I(W678), .ZN(O666));
  INVX1 G6492 (.I(W467), .ZN(W2621));
  INVX1 G6493 (.I(W30), .ZN(W2620));
  INVX1 G6494 (.I(W3697), .ZN(O1463));
  INVX1 G6495 (.I(W1737), .ZN(W4968));
  INVX1 G6496 (.I(I20), .ZN(W1105));
  INVX1 G6497 (.I(W1699), .ZN(W2618));
  INVX1 G6498 (.I(W1365), .ZN(O247));
  INVX1 G6499 (.I(W869), .ZN(W3956));
  INVX1 G6500 (.I(W2486), .ZN(W4973));
  INVX1 G6501 (.I(W1055), .ZN(O246));
endmodule
